magic
tech sky130A
magscale 1 2
timestamp 1653584426
<< locali >>
rect 16221 42211 16255 42313
rect 29009 42007 29043 42245
rect 18797 41599 18831 41701
rect 26801 40035 26835 40137
rect 4261 39423 4295 39593
rect 22569 38811 22603 38913
rect 22845 38811 22879 39049
rect 27169 38947 27203 39049
rect 17141 38335 17175 38437
rect 28549 38335 28583 38437
rect 12541 37655 12575 37757
rect 14013 37655 14047 37825
rect 24685 37655 24719 37825
rect 8585 37179 8619 37417
rect 25053 37247 25087 37349
rect 9045 36771 9079 36873
rect 10149 36635 10183 36737
rect 11161 36567 11195 36805
rect 12173 36567 12207 36805
rect 18521 36635 18555 36873
rect 20453 36771 20487 36873
rect 7941 36023 7975 36329
rect 17417 35003 17451 35173
rect 18061 35003 18095 35241
rect 29101 35071 29135 35173
rect 3709 34527 3743 34697
rect 22661 34459 22695 34629
rect 28365 34459 28399 34561
rect 12817 33507 12851 33609
rect 3341 32895 3375 33065
rect 5457 32997 5549 33031
rect 5457 32827 5491 32997
rect 23213 32827 23247 33065
rect 12541 32215 12575 32453
rect 21649 32215 21683 32385
rect 22201 32215 22235 32317
rect 10885 31807 10919 31977
rect 21005 31671 21039 31977
rect 8125 31127 8159 31365
rect 17233 31195 17267 31433
rect 18429 31331 18463 31433
rect 12449 30583 12483 30821
rect 14749 30583 14783 30753
rect 17417 30039 17451 30277
rect 18245 30107 18279 30141
rect 19809 30107 19843 30209
rect 18245 30073 18429 30107
rect 17141 29631 17175 29733
rect 22477 28951 22511 29257
rect 21741 28543 21775 28713
rect 10793 28407 10827 28509
rect 22385 28407 22419 28441
rect 22385 28373 22569 28407
rect 21649 28067 21683 28169
rect 8953 27863 8987 28033
rect 23857 27863 23891 28169
rect 27537 27863 27571 28169
rect 28825 28067 28859 28169
rect 30205 27863 30239 28033
rect 8493 27319 8527 27489
rect 18889 27319 18923 27489
rect 11161 26775 11195 27013
rect 12541 26775 12575 26945
rect 14105 26911 14139 27081
rect 23581 26775 23615 27013
rect 13093 26299 13127 26537
rect 18153 26231 18187 26401
rect 22569 26299 22603 26469
rect 6101 25279 6135 25449
rect 6193 25279 6227 25381
rect 7941 25211 7975 25381
rect 13921 25279 13955 25449
rect 16221 24735 16255 24837
rect 18889 24599 18923 24769
rect 2329 24123 2363 24361
rect 8125 24191 8159 24361
rect 13737 24191 13771 24361
rect 13679 24157 13771 24191
rect 18061 23511 18095 23681
rect 11345 22491 11379 22729
rect 5917 21947 5951 22185
rect 7481 22083 7515 22185
rect 11805 21879 11839 22117
rect 15669 22083 15703 22185
rect 15669 21879 15703 22049
rect 16071 21913 16313 21947
rect 10609 21403 10643 21505
rect 11989 21471 12023 21641
rect 12817 21403 12851 21573
rect 18153 21403 18187 21505
rect 22477 21335 22511 21641
rect 22753 21539 22787 21641
rect 7665 20859 7699 21029
rect 17785 20791 17819 21097
rect 22569 20791 22603 20961
rect 11379 20417 11563 20451
rect 11529 20315 11563 20417
rect 16497 20315 16531 20485
rect 17877 20247 17911 20485
rect 19441 20247 19475 20485
rect 13645 19839 13679 20009
rect 17785 19703 17819 20009
rect 24225 19839 24259 20009
rect 25053 19839 25087 20009
rect 17727 19669 17819 19703
rect 949 15895 983 19669
rect 11345 19159 11379 19193
rect 11011 19125 11379 19159
rect 16497 19159 16531 19465
rect 17049 19159 17083 19329
rect 17141 19227 17175 19465
rect 18095 19329 18187 19363
rect 18153 19159 18187 19329
rect 18245 19159 18279 19465
rect 19165 19363 19199 19465
rect 27997 19159 28031 19465
rect 9689 18615 9723 18921
rect 13829 18819 13863 18921
rect 17693 18819 17727 18921
rect 13737 18615 13771 18785
rect 27261 18683 27295 18785
rect 3709 18207 3743 18377
rect 6929 18275 6963 18377
rect 24317 18071 24351 18377
rect 26801 18071 26835 18377
rect 29653 18207 29687 18377
rect 11345 17595 11379 17697
rect 11437 17527 11471 17765
rect 12265 17595 12299 17765
rect 12357 17663 12391 17765
rect 23213 17663 23247 17833
rect 12541 17527 12575 17629
rect 17635 17493 17693 17527
rect 17233 17119 17267 17289
rect 17509 17051 17543 17221
rect 24409 16577 24443 16745
rect 24225 16543 24443 16577
rect 16129 16439 16163 16541
rect 24225 16439 24259 16543
rect 23983 16405 24259 16439
rect 5917 16099 5951 16201
rect 16129 16031 16163 16133
rect 16681 15963 16715 16133
rect 24961 16031 24995 16201
rect 25789 16031 25823 16201
rect 13679 15589 13771 15623
rect 7113 15351 7147 15589
rect 7297 15419 7331 15521
rect 13737 15487 13771 15589
rect 13645 15351 13679 15453
rect 24041 15351 24075 15453
rect 14139 15317 14289 15351
rect 4353 14875 4387 15113
rect 15485 14807 15519 15045
rect 16497 15011 16531 15113
rect 17877 15011 17911 15113
rect 24869 14875 24903 14977
rect 9873 14263 9907 14365
rect 15301 14263 15335 14569
rect 17693 14399 17727 14501
rect 8953 13923 8987 14025
rect 14289 13719 14323 13889
rect 15301 13719 15335 13957
rect 23949 13719 23983 13957
rect 29929 13787 29963 13957
rect 15393 13311 15427 13413
rect 18429 13175 18463 13481
rect 28549 13311 28583 13481
rect 4629 12835 4663 12937
rect 10149 12631 10183 12733
rect 4445 11611 4479 11713
rect 8769 10999 8803 11237
rect 29101 11067 29135 11237
rect 7757 10591 7791 10693
rect 8493 10591 8527 10693
rect 20545 10659 20579 10761
rect 7757 10557 7849 10591
rect 10977 10455 11011 10625
rect 16313 9979 16347 10081
rect 5549 9435 5583 9673
rect 8769 9367 8803 9605
rect 8861 9503 8895 9605
rect 24685 9469 24869 9503
rect 24685 9435 24719 9469
rect 2973 8891 3007 8993
rect 4445 8823 4479 9129
rect 5549 9027 5583 9129
rect 8769 8823 8803 8925
rect 20085 8823 20119 8925
rect 22845 8823 22879 8857
rect 22845 8789 23029 8823
rect 3433 8347 3467 8517
rect 24869 8347 24903 8449
rect 25697 8347 25731 8449
rect 9965 7871 9999 7973
rect 11069 7871 11103 7973
rect 27077 7871 27111 8041
rect 9965 7735 9999 7837
rect 6193 7259 6227 7497
rect 32137 6919 32171 8109
rect 12817 6103 12851 6205
rect 27721 6171 27755 6409
rect 4721 5627 4755 5797
rect 29929 5695 29963 5865
rect 15301 5559 15335 5661
rect 26709 5559 26743 5661
rect 6193 5015 6227 5117
rect 16681 5083 16715 5185
rect 18153 4675 18187 4777
rect 949 2431 983 4505
rect 13645 4471 13679 4641
rect 19533 4607 19567 4777
rect 18889 4471 18923 4573
rect 15117 4131 15151 4233
rect 3525 3519 3559 3621
rect 6009 2839 6043 3077
rect 7389 2907 7423 3009
rect 11161 2839 11195 3077
rect 18889 3043 18923 3145
rect 18061 2907 18095 3009
rect 21189 2839 21223 3009
rect 6377 2295 6411 2601
rect 24409 2499 24443 2601
rect 28917 2431 28951 2601
rect 30297 2431 30331 2533
rect 13001 1207 13035 1309
rect 14381 1207 14415 1513
rect 15301 1207 15335 1309
rect 17233 1207 17267 1309
rect 21373 1207 21407 1309
rect 25237 1207 25271 1309
rect 27537 1275 27571 1445
rect 17233 663 17267 969
<< viali >>
rect 4353 42313 4387 42347
rect 7481 42313 7515 42347
rect 16221 42313 16255 42347
rect 21189 42313 21223 42347
rect 22293 42313 22327 42347
rect 4261 42245 4295 42279
rect 23673 42245 23707 42279
rect 29009 42245 29043 42279
rect 1869 42177 1903 42211
rect 2881 42177 2915 42211
rect 7665 42177 7699 42211
rect 8217 42177 8251 42211
rect 9137 42177 9171 42211
rect 10057 42177 10091 42211
rect 12725 42177 12759 42211
rect 15393 42177 15427 42211
rect 15945 42177 15979 42211
rect 16221 42177 16255 42211
rect 16865 42177 16899 42211
rect 18153 42177 18187 42211
rect 20065 42177 20099 42211
rect 22477 42177 22511 42211
rect 23121 42177 23155 42211
rect 24593 42177 24627 42211
rect 25789 42177 25823 42211
rect 26433 42177 26467 42211
rect 27169 42177 27203 42211
rect 28641 42177 28675 42211
rect 3157 42109 3191 42143
rect 9413 42109 9447 42143
rect 13001 42109 13035 42143
rect 17141 42109 17175 42143
rect 18429 42109 18463 42143
rect 19809 42109 19843 42143
rect 27445 42109 27479 42143
rect 28917 42109 28951 42143
rect 3065 42041 3099 42075
rect 9873 42041 9907 42075
rect 16129 42041 16163 42075
rect 17049 42041 17083 42075
rect 17969 42041 18003 42075
rect 24409 42041 24443 42075
rect 29745 42177 29779 42211
rect 30389 42177 30423 42211
rect 31309 42177 31343 42211
rect 30205 42041 30239 42075
rect 31125 42041 31159 42075
rect 1961 41973 1995 42007
rect 2697 41973 2731 42007
rect 8309 41973 8343 42007
rect 8953 41973 8987 42007
rect 9321 41973 9355 42007
rect 12541 41973 12575 42007
rect 12909 41973 12943 42007
rect 15209 41973 15243 42007
rect 16681 41973 16715 42007
rect 18337 41973 18371 42007
rect 22937 41973 22971 42007
rect 23765 41973 23799 42007
rect 25605 41973 25639 42007
rect 26249 41973 26283 42007
rect 26985 41973 27019 42007
rect 27353 41973 27387 42007
rect 28457 41973 28491 42007
rect 28825 41973 28859 42007
rect 29009 41973 29043 42007
rect 29561 41973 29595 42007
rect 6193 41769 6227 41803
rect 8401 41769 8435 41803
rect 19625 41769 19659 41803
rect 26617 41769 26651 41803
rect 3249 41701 3283 41735
rect 9321 41701 9355 41735
rect 18797 41701 18831 41735
rect 25789 41701 25823 41735
rect 29009 41701 29043 41735
rect 6285 41633 6319 41667
rect 9413 41633 9447 41667
rect 18061 41633 18095 41667
rect 19717 41633 19751 41667
rect 26709 41633 26743 41667
rect 29929 41633 29963 41667
rect 1869 41565 1903 41599
rect 2136 41565 2170 41599
rect 3985 41565 4019 41599
rect 4169 41565 4203 41599
rect 4261 41565 4295 41599
rect 4905 41565 4939 41599
rect 5181 41565 5215 41599
rect 5365 41565 5399 41599
rect 6009 41565 6043 41599
rect 7021 41565 7055 41599
rect 9137 41565 9171 41599
rect 10057 41565 10091 41599
rect 12081 41565 12115 41599
rect 12348 41565 12382 41599
rect 14105 41565 14139 41599
rect 15945 41565 15979 41599
rect 16212 41565 16246 41599
rect 18245 41565 18279 41599
rect 18521 41565 18555 41599
rect 18705 41565 18739 41599
rect 18797 41565 18831 41599
rect 19441 41565 19475 41599
rect 20637 41565 20671 41599
rect 22477 41565 22511 41599
rect 24409 41565 24443 41599
rect 26433 41565 26467 41599
rect 27629 41565 27663 41599
rect 27896 41565 27930 41599
rect 29745 41565 29779 41599
rect 30021 41565 30055 41599
rect 30665 41565 30699 41599
rect 31309 41565 31343 41599
rect 4721 41497 4755 41531
rect 7288 41497 7322 41531
rect 8953 41497 8987 41531
rect 10324 41497 10358 41531
rect 14372 41497 14406 41531
rect 20904 41497 20938 41531
rect 22744 41497 22778 41531
rect 24676 41497 24710 41531
rect 3801 41429 3835 41463
rect 5825 41429 5859 41463
rect 11437 41429 11471 41463
rect 13461 41429 13495 41463
rect 15485 41429 15519 41463
rect 17325 41429 17359 41463
rect 19257 41429 19291 41463
rect 22017 41429 22051 41463
rect 23857 41429 23891 41463
rect 26249 41429 26283 41463
rect 29561 41429 29595 41463
rect 30481 41429 30515 41463
rect 31125 41429 31159 41463
rect 10333 41225 10367 41259
rect 13461 41225 13495 41259
rect 15669 41225 15703 41259
rect 8668 41157 8702 41191
rect 14565 41157 14599 41191
rect 18766 41157 18800 41191
rect 25320 41157 25354 41191
rect 27252 41157 27286 41191
rect 1409 41089 1443 41123
rect 1676 41089 1710 41123
rect 3801 41089 3835 41123
rect 4057 41089 4091 41123
rect 6377 41089 6411 41123
rect 6644 41089 6678 41123
rect 8401 41089 8435 41123
rect 10517 41089 10551 41123
rect 11621 41089 11655 41123
rect 11888 41089 11922 41123
rect 13645 41089 13679 41123
rect 13921 41089 13955 41123
rect 14105 41089 14139 41123
rect 14749 41089 14783 41123
rect 15025 41089 15059 41123
rect 15209 41089 15243 41123
rect 15853 41089 15887 41123
rect 16681 41089 16715 41123
rect 16937 41089 16971 41123
rect 18521 41089 18555 41123
rect 20637 41089 20671 41123
rect 21281 41089 21315 41123
rect 22100 41089 22134 41123
rect 23673 41089 23707 41123
rect 23857 41089 23891 41123
rect 26985 41089 27019 41123
rect 28825 41089 28859 41123
rect 29081 41089 29115 41123
rect 30849 41089 30883 41123
rect 10793 41021 10827 41055
rect 16129 41021 16163 41055
rect 21833 41021 21867 41055
rect 24133 41021 24167 41055
rect 25053 41021 25087 41055
rect 20453 40953 20487 40987
rect 30205 40953 30239 40987
rect 2789 40885 2823 40919
rect 5181 40885 5215 40919
rect 7757 40885 7791 40919
rect 9781 40885 9815 40919
rect 10701 40885 10735 40919
rect 13001 40885 13035 40919
rect 16037 40885 16071 40919
rect 18061 40885 18095 40919
rect 19901 40885 19935 40919
rect 21097 40885 21131 40919
rect 23213 40885 23247 40919
rect 24041 40885 24075 40919
rect 26433 40885 26467 40919
rect 28365 40885 28399 40919
rect 30665 40885 30699 40919
rect 1685 40681 1719 40715
rect 3801 40681 3835 40715
rect 7021 40681 7055 40715
rect 16405 40681 16439 40715
rect 22201 40681 22235 40715
rect 23305 40681 23339 40715
rect 27353 40681 27387 40715
rect 28457 40681 28491 40715
rect 7941 40613 7975 40647
rect 2145 40545 2179 40579
rect 8401 40545 8435 40579
rect 9413 40545 9447 40579
rect 19257 40545 19291 40579
rect 29561 40545 29595 40579
rect 1869 40477 1903 40511
rect 2053 40477 2087 40511
rect 2789 40477 2823 40511
rect 3065 40477 3099 40511
rect 3249 40477 3283 40511
rect 3985 40477 4019 40511
rect 4261 40477 4295 40511
rect 4445 40477 4479 40511
rect 8125 40477 8159 40511
rect 8309 40477 8343 40511
rect 11437 40477 11471 40511
rect 11713 40477 11747 40511
rect 11897 40477 11931 40511
rect 13001 40477 13035 40511
rect 13277 40477 13311 40511
rect 13461 40477 13495 40511
rect 14565 40477 14599 40511
rect 16589 40477 16623 40511
rect 16865 40477 16899 40511
rect 17049 40477 17083 40511
rect 17693 40477 17727 40511
rect 17969 40477 18003 40511
rect 18153 40477 18187 40511
rect 19513 40477 19547 40511
rect 21741 40477 21775 40511
rect 22385 40477 22419 40511
rect 22661 40477 22695 40511
rect 22845 40477 22879 40511
rect 23489 40477 23523 40511
rect 23673 40477 23707 40511
rect 23765 40477 23799 40511
rect 24409 40477 24443 40511
rect 26433 40477 26467 40511
rect 26709 40477 26743 40511
rect 26893 40477 26927 40511
rect 27537 40477 27571 40511
rect 27813 40477 27847 40511
rect 27997 40477 28031 40511
rect 28641 40477 28675 40511
rect 28825 40477 28859 40511
rect 28917 40477 28951 40511
rect 29817 40477 29851 40511
rect 2605 40409 2639 40443
rect 5733 40409 5767 40443
rect 9680 40409 9714 40443
rect 14832 40409 14866 40443
rect 24654 40409 24688 40443
rect 10793 40341 10827 40375
rect 11253 40341 11287 40375
rect 12817 40341 12851 40375
rect 15945 40341 15979 40375
rect 17509 40341 17543 40375
rect 20637 40341 20671 40375
rect 21557 40341 21591 40375
rect 25789 40341 25823 40375
rect 26249 40341 26283 40375
rect 30941 40341 30975 40375
rect 3341 40137 3375 40171
rect 5825 40137 5859 40171
rect 7573 40137 7607 40171
rect 8861 40137 8895 40171
rect 9965 40137 9999 40171
rect 11529 40137 11563 40171
rect 19717 40137 19751 40171
rect 22845 40137 22879 40171
rect 26801 40137 26835 40171
rect 26985 40137 27019 40171
rect 28089 40137 28123 40171
rect 29193 40137 29227 40171
rect 6837 40069 6871 40103
rect 14197 40069 14231 40103
rect 16681 40069 16715 40103
rect 25421 40069 25455 40103
rect 30297 40069 30331 40103
rect 1676 40001 1710 40035
rect 3525 40001 3559 40035
rect 3801 40001 3835 40035
rect 3985 40001 4019 40035
rect 4445 40001 4479 40035
rect 4712 40001 4746 40035
rect 6561 40001 6595 40035
rect 6745 40001 6779 40035
rect 6929 40001 6963 40035
rect 7757 40001 7791 40035
rect 8033 40001 8067 40035
rect 8217 40001 8251 40035
rect 9045 40001 9079 40035
rect 9321 40001 9355 40035
rect 9505 40001 9539 40035
rect 10149 40001 10183 40035
rect 11713 40001 11747 40035
rect 11989 40001 12023 40035
rect 12173 40001 12207 40035
rect 12633 40001 12667 40035
rect 12817 40001 12851 40035
rect 13737 40001 13771 40035
rect 14381 40001 14415 40035
rect 14657 40001 14691 40035
rect 14841 40001 14875 40035
rect 15301 40001 15335 40035
rect 15485 40001 15519 40035
rect 16865 40001 16899 40035
rect 17141 40001 17175 40035
rect 17325 40001 17359 40035
rect 17969 40001 18003 40035
rect 18705 40001 18739 40035
rect 19901 40001 19935 40035
rect 21833 40001 21867 40035
rect 22017 40001 22051 40035
rect 23029 40001 23063 40035
rect 23305 40001 23339 40035
rect 23489 40001 23523 40035
rect 25605 40001 25639 40035
rect 25881 40001 25915 40035
rect 26065 40001 26099 40035
rect 26801 40001 26835 40035
rect 27169 40001 27203 40035
rect 27445 40001 27479 40035
rect 27629 40001 27663 40035
rect 28273 40001 28307 40035
rect 28549 40001 28583 40035
rect 28733 40001 28767 40035
rect 29377 40001 29411 40035
rect 29653 40001 29687 40035
rect 29837 40001 29871 40035
rect 30481 40001 30515 40035
rect 30757 40001 30791 40035
rect 30941 40001 30975 40035
rect 1409 39933 1443 39967
rect 10425 39933 10459 39967
rect 13093 39933 13127 39967
rect 15761 39933 15795 39967
rect 18429 39933 18463 39967
rect 20361 39933 20395 39967
rect 20637 39933 20671 39967
rect 22293 39933 22327 39967
rect 24133 39933 24167 39967
rect 24409 39933 24443 39967
rect 13553 39865 13587 39899
rect 17785 39865 17819 39899
rect 2789 39797 2823 39831
rect 7113 39797 7147 39831
rect 10333 39797 10367 39831
rect 13001 39797 13035 39831
rect 15669 39797 15703 39831
rect 22201 39797 22235 39831
rect 2605 39593 2639 39627
rect 4261 39593 4295 39627
rect 7757 39593 7791 39627
rect 12265 39593 12299 39627
rect 16773 39593 16807 39627
rect 18061 39593 18095 39627
rect 22845 39593 22879 39627
rect 24409 39593 24443 39627
rect 2973 39457 3007 39491
rect 7297 39525 7331 39559
rect 15761 39525 15795 39559
rect 17141 39525 17175 39559
rect 24777 39525 24811 39559
rect 28733 39525 28767 39559
rect 4629 39457 4663 39491
rect 9229 39457 9263 39491
rect 12817 39457 12851 39491
rect 14381 39457 14415 39491
rect 17233 39457 17267 39491
rect 19625 39457 19659 39491
rect 24869 39457 24903 39491
rect 27629 39457 27663 39491
rect 29929 39457 29963 39491
rect 2789 39389 2823 39423
rect 3065 39389 3099 39423
rect 4261 39389 4295 39423
rect 4353 39389 4387 39423
rect 5641 39389 5675 39423
rect 5917 39389 5951 39423
rect 6009 39389 6043 39423
rect 6745 39389 6779 39423
rect 7113 39389 7147 39423
rect 7941 39389 7975 39423
rect 8217 39389 8251 39423
rect 8401 39389 8435 39423
rect 8953 39389 8987 39423
rect 10609 39389 10643 39423
rect 10793 39389 10827 39423
rect 10885 39389 10919 39423
rect 12081 39389 12115 39423
rect 12357 39389 12391 39423
rect 13001 39389 13035 39423
rect 13277 39389 13311 39423
rect 13461 39389 13495 39423
rect 14105 39389 14139 39423
rect 15577 39389 15611 39423
rect 15853 39389 15887 39423
rect 16957 39389 16991 39423
rect 18245 39389 18279 39423
rect 18521 39389 18555 39423
rect 18705 39389 18739 39423
rect 19441 39389 19475 39423
rect 19717 39389 19751 39423
rect 23029 39389 23063 39423
rect 23305 39389 23339 39423
rect 23489 39389 23523 39423
rect 24593 39389 24627 39423
rect 25881 39389 25915 39423
rect 26249 39389 26283 39423
rect 27353 39389 27387 39423
rect 28641 39389 28675 39423
rect 1777 39321 1811 39355
rect 5825 39321 5859 39355
rect 6929 39321 6963 39355
rect 7021 39321 7055 39355
rect 20637 39321 20671 39355
rect 26065 39321 26099 39355
rect 26157 39321 26191 39355
rect 30196 39321 30230 39355
rect 1869 39253 1903 39287
rect 6193 39253 6227 39287
rect 10425 39253 10459 39287
rect 11897 39253 11931 39287
rect 15393 39253 15427 39287
rect 19257 39253 19291 39287
rect 21925 39253 21959 39287
rect 26433 39253 26467 39287
rect 31309 39253 31343 39287
rect 3157 39049 3191 39083
rect 6377 39049 6411 39083
rect 10333 39049 10367 39083
rect 16037 39049 16071 39083
rect 21833 39049 21867 39083
rect 22845 39049 22879 39083
rect 7021 38981 7055 39015
rect 14280 38981 14314 39015
rect 17509 38981 17543 39015
rect 17601 38981 17635 39015
rect 2421 38913 2455 38947
rect 3341 38913 3375 38947
rect 3617 38913 3651 38947
rect 3801 38913 3835 38947
rect 4445 38913 4479 38947
rect 5089 38913 5123 38947
rect 5182 38913 5216 38947
rect 5365 38913 5399 38947
rect 5457 38913 5491 38947
rect 5595 38913 5629 38947
rect 6561 38913 6595 38947
rect 7205 38913 7239 38947
rect 7481 38913 7515 38947
rect 7665 38913 7699 38947
rect 8309 38913 8343 38947
rect 8585 38913 8619 38947
rect 8769 38913 8803 38947
rect 9413 38913 9447 38947
rect 9689 38913 9723 38947
rect 10517 38913 10551 38947
rect 10793 38913 10827 38947
rect 10977 38913 11011 38947
rect 11897 38913 11931 38947
rect 12153 38913 12187 38947
rect 15945 38913 15979 38947
rect 17233 38913 17267 38947
rect 17325 38913 17359 38947
rect 17693 38913 17727 38947
rect 18245 38913 18279 38947
rect 18512 38913 18546 38947
rect 20177 38913 20211 38947
rect 20453 38913 20487 38947
rect 22017 38913 22051 38947
rect 22293 38913 22327 38947
rect 22477 38913 22511 38947
rect 22569 38913 22603 38947
rect 2697 38845 2731 38879
rect 14013 38845 14047 38879
rect 4629 38777 4663 38811
rect 9597 38777 9631 38811
rect 15393 38777 15427 38811
rect 22569 38777 22603 38811
rect 27169 39049 27203 39083
rect 30481 39049 30515 39083
rect 27445 38981 27479 39015
rect 27537 38981 27571 39015
rect 23121 38913 23155 38947
rect 23397 38913 23431 38947
rect 23581 38913 23615 38947
rect 24041 38913 24075 38947
rect 24225 38913 24259 38947
rect 24685 38913 24719 38947
rect 27169 38913 27203 38947
rect 27261 38913 27295 38947
rect 27629 38913 27663 38947
rect 28457 38913 28491 38947
rect 28641 38913 28675 38947
rect 30665 38913 30699 38947
rect 30849 38913 30883 38947
rect 28733 38845 28767 38879
rect 29193 38845 29227 38879
rect 29469 38845 29503 38879
rect 30941 38845 30975 38879
rect 22845 38777 22879 38811
rect 28273 38777 28307 38811
rect 2237 38709 2271 38743
rect 2605 38709 2639 38743
rect 5733 38709 5767 38743
rect 8125 38709 8159 38743
rect 9229 38709 9263 38743
rect 13277 38709 13311 38743
rect 17233 38709 17267 38743
rect 19625 38709 19659 38743
rect 22937 38709 22971 38743
rect 24041 38709 24075 38743
rect 25973 38709 26007 38743
rect 27813 38709 27847 38743
rect 3249 38505 3283 38539
rect 5457 38505 5491 38539
rect 8309 38505 8343 38539
rect 11897 38505 11931 38539
rect 14105 38505 14139 38539
rect 17785 38505 17819 38539
rect 18613 38505 18647 38539
rect 23029 38505 23063 38539
rect 28641 38505 28675 38539
rect 29561 38505 29595 38539
rect 31033 38505 31067 38539
rect 7665 38437 7699 38471
rect 9505 38437 9539 38471
rect 16313 38437 16347 38471
rect 17141 38437 17175 38471
rect 28181 38437 28215 38471
rect 28549 38437 28583 38471
rect 29009 38437 29043 38471
rect 6285 38369 6319 38403
rect 18705 38369 18739 38403
rect 26617 38369 26651 38403
rect 31125 38369 31159 38403
rect 1869 38301 1903 38335
rect 4077 38301 4111 38335
rect 4353 38301 4387 38335
rect 4445 38301 4479 38335
rect 5365 38301 5399 38335
rect 5549 38301 5583 38335
rect 6552 38301 6586 38335
rect 8953 38301 8987 38335
rect 9229 38301 9263 38335
rect 9321 38301 9355 38335
rect 10149 38301 10183 38335
rect 13001 38301 13035 38335
rect 13277 38301 13311 38335
rect 13461 38301 13495 38335
rect 14105 38301 14139 38335
rect 14197 38301 14231 38335
rect 17141 38301 17175 38335
rect 17233 38301 17267 38335
rect 17417 38301 17451 38335
rect 17509 38301 17543 38335
rect 17647 38301 17681 38335
rect 18429 38301 18463 38335
rect 19809 38301 19843 38335
rect 21649 38301 21683 38335
rect 23673 38301 23707 38335
rect 24409 38301 24443 38335
rect 24502 38301 24536 38335
rect 24777 38301 24811 38335
rect 24874 38301 24908 38335
rect 25697 38301 25731 38335
rect 26157 38301 26191 38335
rect 26801 38301 26835 38335
rect 26893 38301 26927 38335
rect 27077 38301 27111 38335
rect 27169 38301 27203 38335
rect 27629 38301 27663 38335
rect 27813 38301 27847 38335
rect 27997 38301 28031 38335
rect 28549 38301 28583 38335
rect 28641 38301 28675 38335
rect 28733 38301 28767 38335
rect 29745 38301 29779 38335
rect 30021 38301 30055 38335
rect 30205 38301 30239 38335
rect 30849 38301 30883 38335
rect 2136 38233 2170 38267
rect 4261 38233 4295 38267
rect 8217 38233 8251 38267
rect 9137 38233 9171 38267
rect 10609 38233 10643 38267
rect 15025 38233 15059 38267
rect 20076 38233 20110 38267
rect 21916 38233 21950 38267
rect 24685 38233 24719 38267
rect 25789 38233 25823 38267
rect 25881 38233 25915 38267
rect 26019 38233 26053 38267
rect 27905 38233 27939 38267
rect 4629 38165 4663 38199
rect 5733 38165 5767 38199
rect 9965 38165 9999 38199
rect 12817 38165 12851 38199
rect 14473 38165 14507 38199
rect 18245 38165 18279 38199
rect 21189 38165 21223 38199
rect 23765 38165 23799 38199
rect 25053 38165 25087 38199
rect 25513 38165 25547 38199
rect 30665 38165 30699 38199
rect 2697 37961 2731 37995
rect 5733 37961 5767 37995
rect 8401 37961 8435 37995
rect 10885 37961 10919 37995
rect 18889 37961 18923 37995
rect 21189 37961 21223 37995
rect 22109 37961 22143 37995
rect 23489 37961 23523 37995
rect 25329 37961 25363 37995
rect 27629 37961 27663 37995
rect 15485 37893 15519 37927
rect 17316 37893 17350 37927
rect 23121 37893 23155 37927
rect 23337 37893 23371 37927
rect 30196 37893 30230 37927
rect 1869 37825 1903 37859
rect 2881 37825 2915 37859
rect 3157 37825 3191 37859
rect 3341 37825 3375 37859
rect 4077 37825 4111 37859
rect 5549 37825 5583 37859
rect 6561 37825 6595 37859
rect 7288 37825 7322 37859
rect 9505 37825 9539 37859
rect 9772 37825 9806 37859
rect 11897 37825 11931 37859
rect 12633 37825 12667 37859
rect 14013 37825 14047 37859
rect 14105 37825 14139 37859
rect 14289 37825 14323 37859
rect 14381 37825 14415 37859
rect 14473 37825 14507 37859
rect 15117 37825 15151 37859
rect 15210 37825 15244 37859
rect 15393 37825 15427 37859
rect 15582 37825 15616 37859
rect 19073 37825 19107 37859
rect 19349 37825 19383 37859
rect 19809 37825 19843 37859
rect 20076 37825 20110 37859
rect 22293 37825 22327 37859
rect 22477 37825 22511 37859
rect 24225 37825 24259 37859
rect 24317 37825 24351 37859
rect 24501 37825 24535 37859
rect 24593 37825 24627 37859
rect 24685 37825 24719 37859
rect 25513 37825 25547 37859
rect 25789 37825 25823 37859
rect 25973 37825 26007 37859
rect 26985 37825 27019 37859
rect 27078 37825 27112 37859
rect 27261 37825 27295 37859
rect 27361 37825 27395 37859
rect 27491 37825 27525 37859
rect 28089 37825 28123 37859
rect 28356 37825 28390 37859
rect 4353 37757 4387 37791
rect 7021 37757 7055 37791
rect 12173 37757 12207 37791
rect 12541 37757 12575 37791
rect 12909 37757 12943 37791
rect 2145 37621 2179 37655
rect 6377 37621 6411 37655
rect 11713 37621 11747 37655
rect 12081 37621 12115 37655
rect 12541 37621 12575 37655
rect 17049 37757 17083 37791
rect 19257 37757 19291 37791
rect 22569 37757 22603 37791
rect 24041 37757 24075 37791
rect 14657 37689 14691 37723
rect 29929 37757 29963 37791
rect 14013 37621 14047 37655
rect 15761 37621 15795 37655
rect 18429 37621 18463 37655
rect 23305 37621 23339 37655
rect 24685 37621 24719 37655
rect 29469 37621 29503 37655
rect 31309 37621 31343 37655
rect 2789 37417 2823 37451
rect 7573 37417 7607 37451
rect 8585 37417 8619 37451
rect 11621 37417 11655 37451
rect 16681 37417 16715 37451
rect 20637 37417 20671 37451
rect 22937 37417 22971 37451
rect 23673 37417 23707 37451
rect 23857 37417 23891 37451
rect 25789 37417 25823 37451
rect 27905 37417 27939 37451
rect 6101 37281 6135 37315
rect 7113 37281 7147 37315
rect 8033 37281 8067 37315
rect 1409 37213 1443 37247
rect 4353 37213 4387 37247
rect 4446 37213 4480 37247
rect 4629 37213 4663 37247
rect 4859 37213 4893 37247
rect 5825 37213 5859 37247
rect 6837 37213 6871 37247
rect 7021 37213 7055 37247
rect 7757 37213 7791 37247
rect 7941 37213 7975 37247
rect 13553 37349 13587 37383
rect 21833 37349 21867 37383
rect 25053 37349 25087 37383
rect 26709 37349 26743 37383
rect 10885 37281 10919 37315
rect 12173 37281 12207 37315
rect 15669 37281 15703 37315
rect 19349 37281 19383 37315
rect 21097 37281 21131 37315
rect 9045 37213 9079 37247
rect 9229 37213 9263 37247
rect 10517 37213 10551 37247
rect 10609 37213 10643 37247
rect 10977 37213 11011 37247
rect 14565 37213 14599 37247
rect 14658 37213 14692 37247
rect 14933 37213 14967 37247
rect 15071 37213 15105 37247
rect 15853 37213 15887 37247
rect 17785 37213 17819 37247
rect 17969 37213 18003 37247
rect 18245 37213 18279 37247
rect 18441 37213 18475 37247
rect 19625 37213 19659 37247
rect 20821 37213 20855 37247
rect 21005 37213 21039 37247
rect 21649 37213 21683 37247
rect 22845 37213 22879 37247
rect 23029 37213 23063 37247
rect 24409 37213 24443 37247
rect 24593 37213 24627 37247
rect 24961 37213 24995 37247
rect 25053 37213 25087 37247
rect 25973 37213 26007 37247
rect 26157 37213 26191 37247
rect 26249 37213 26283 37247
rect 26709 37213 26743 37247
rect 26893 37213 26927 37247
rect 27353 37213 27387 37247
rect 27721 37213 27755 37247
rect 28549 37213 28583 37247
rect 28825 37213 28859 37247
rect 29021 37213 29055 37247
rect 1654 37145 1688 37179
rect 4721 37145 4755 37179
rect 5917 37145 5951 37179
rect 8585 37145 8619 37179
rect 11529 37145 11563 37179
rect 12418 37145 12452 37179
rect 14841 37145 14875 37179
rect 16037 37145 16071 37179
rect 16589 37145 16623 37179
rect 23489 37145 23523 37179
rect 27537 37145 27571 37179
rect 27629 37145 27663 37179
rect 29561 37145 29595 37179
rect 4997 37077 5031 37111
rect 5457 37077 5491 37111
rect 6653 37077 6687 37111
rect 9137 37077 9171 37111
rect 10333 37077 10367 37111
rect 15209 37077 15243 37111
rect 23699 37077 23733 37111
rect 24869 37077 24903 37111
rect 28365 37077 28399 37111
rect 30849 37077 30883 37111
rect 1409 36873 1443 36907
rect 5273 36873 5307 36907
rect 8033 36873 8067 36907
rect 9045 36873 9079 36907
rect 11805 36873 11839 36907
rect 14657 36873 14691 36907
rect 15761 36873 15795 36907
rect 15853 36873 15887 36907
rect 16865 36873 16899 36907
rect 18521 36873 18555 36907
rect 18613 36873 18647 36907
rect 19717 36873 19751 36907
rect 20453 36873 20487 36907
rect 30205 36873 30239 36907
rect 4997 36805 5031 36839
rect 9781 36805 9815 36839
rect 11161 36805 11195 36839
rect 11897 36805 11931 36839
rect 12173 36805 12207 36839
rect 1593 36737 1627 36771
rect 2329 36737 2363 36771
rect 2513 36737 2547 36771
rect 2789 36737 2823 36771
rect 2973 36737 3007 36771
rect 3801 36737 3835 36771
rect 4077 36737 4111 36771
rect 4261 36737 4295 36771
rect 4721 36737 4755 36771
rect 4905 36737 4939 36771
rect 5089 36737 5123 36771
rect 6561 36737 6595 36771
rect 7849 36737 7883 36771
rect 8033 36737 8067 36771
rect 8677 36737 8711 36771
rect 8861 36737 8895 36771
rect 9045 36737 9079 36771
rect 9597 36737 9631 36771
rect 10149 36737 10183 36771
rect 10241 36737 10275 36771
rect 10517 36737 10551 36771
rect 1869 36669 1903 36703
rect 6837 36669 6871 36703
rect 9413 36669 9447 36703
rect 8861 36601 8895 36635
rect 10149 36601 10183 36635
rect 10517 36601 10551 36635
rect 11529 36737 11563 36771
rect 11713 36737 11747 36771
rect 12817 36737 12851 36771
rect 13093 36737 13127 36771
rect 13277 36737 13311 36771
rect 14105 36737 14139 36771
rect 14289 36737 14323 36771
rect 14381 36737 14415 36771
rect 14473 36737 14507 36771
rect 16681 36737 16715 36771
rect 16957 36737 16991 36771
rect 17601 36737 17635 36771
rect 16037 36669 16071 36703
rect 17877 36669 17911 36703
rect 23121 36805 23155 36839
rect 18797 36737 18831 36771
rect 19073 36737 19107 36771
rect 19257 36737 19291 36771
rect 19901 36737 19935 36771
rect 20177 36737 20211 36771
rect 20361 36737 20395 36771
rect 20453 36737 20487 36771
rect 20915 36737 20949 36771
rect 21833 36737 21867 36771
rect 22937 36737 22971 36771
rect 24133 36737 24167 36771
rect 25237 36737 25271 36771
rect 25513 36737 25547 36771
rect 26157 36737 26191 36771
rect 26433 36737 26467 36771
rect 27261 36737 27295 36771
rect 27517 36737 27551 36771
rect 29285 36737 29319 36771
rect 30389 36737 30423 36771
rect 30665 36737 30699 36771
rect 30849 36737 30883 36771
rect 29561 36669 29595 36703
rect 18521 36601 18555 36635
rect 22293 36601 22327 36635
rect 24317 36601 24351 36635
rect 25973 36601 26007 36635
rect 29469 36601 29503 36635
rect 1777 36533 1811 36567
rect 3617 36533 3651 36567
rect 6377 36533 6411 36567
rect 6745 36533 6779 36567
rect 11161 36533 11195 36567
rect 12081 36533 12115 36567
rect 12173 36533 12207 36567
rect 12633 36533 12667 36567
rect 15393 36533 15427 36567
rect 16681 36533 16715 36567
rect 17417 36533 17451 36567
rect 17785 36533 17819 36567
rect 21005 36533 21039 36567
rect 21925 36533 21959 36567
rect 25053 36533 25087 36567
rect 25421 36533 25455 36567
rect 26341 36533 26375 36567
rect 28641 36533 28675 36567
rect 29101 36533 29135 36567
rect 7941 36329 7975 36363
rect 8033 36329 8067 36363
rect 8401 36329 8435 36363
rect 9689 36329 9723 36363
rect 10885 36329 10919 36363
rect 11529 36329 11563 36363
rect 23673 36329 23707 36363
rect 27629 36329 27663 36363
rect 28917 36329 28951 36363
rect 1593 36261 1627 36295
rect 7389 36261 7423 36295
rect 5549 36193 5583 36227
rect 1409 36125 1443 36159
rect 2513 36125 2547 36159
rect 2789 36125 2823 36159
rect 2973 36125 3007 36159
rect 3985 36125 4019 36159
rect 4261 36125 4295 36159
rect 4445 36125 4479 36159
rect 5816 36125 5850 36159
rect 7573 36125 7607 36159
rect 13553 36261 13587 36295
rect 14841 36261 14875 36295
rect 16497 36261 16531 36295
rect 17785 36261 17819 36295
rect 27169 36261 27203 36295
rect 9321 36193 9355 36227
rect 10977 36193 11011 36227
rect 25789 36193 25823 36227
rect 29561 36193 29595 36227
rect 8033 36125 8067 36159
rect 8217 36125 8251 36159
rect 9505 36125 9539 36159
rect 10701 36125 10735 36159
rect 11437 36125 11471 36159
rect 11621 36125 11655 36159
rect 12173 36125 12207 36159
rect 14565 36125 14599 36159
rect 14749 36125 14783 36159
rect 15761 36125 15795 36159
rect 16037 36125 16071 36159
rect 16681 36125 16715 36159
rect 16773 36125 16807 36159
rect 16957 36125 16991 36159
rect 17049 36125 17083 36159
rect 17969 36125 18003 36159
rect 18245 36125 18279 36159
rect 18429 36125 18463 36159
rect 19441 36125 19475 36159
rect 19717 36125 19751 36159
rect 19901 36125 19935 36159
rect 20821 36125 20855 36159
rect 22661 36125 22695 36159
rect 23581 36125 23615 36159
rect 23765 36125 23799 36159
rect 24593 36125 24627 36159
rect 24869 36125 24903 36159
rect 25053 36125 25087 36159
rect 27813 36125 27847 36159
rect 28089 36125 28123 36159
rect 28273 36125 28307 36159
rect 29817 36125 29851 36159
rect 12440 36057 12474 36091
rect 15945 36057 15979 36091
rect 21088 36057 21122 36091
rect 22937 36057 22971 36091
rect 24409 36057 24443 36091
rect 26056 36057 26090 36091
rect 28825 36057 28859 36091
rect 2329 35989 2363 36023
rect 3801 35989 3835 36023
rect 6929 35989 6963 36023
rect 7941 35989 7975 36023
rect 10517 35989 10551 36023
rect 15577 35989 15611 36023
rect 19257 35989 19291 36023
rect 22201 35989 22235 36023
rect 30941 35989 30975 36023
rect 2789 35785 2823 35819
rect 14933 35785 14967 35819
rect 3433 35717 3467 35751
rect 6377 35717 6411 35751
rect 13369 35717 13403 35751
rect 14565 35717 14599 35751
rect 14765 35717 14799 35751
rect 15853 35717 15887 35751
rect 30174 35717 30208 35751
rect 1409 35649 1443 35683
rect 1676 35649 1710 35683
rect 6561 35649 6595 35683
rect 6837 35649 6871 35683
rect 7021 35649 7055 35683
rect 7665 35649 7699 35683
rect 7932 35649 7966 35683
rect 10793 35649 10827 35683
rect 10977 35649 11011 35683
rect 11785 35649 11819 35683
rect 13553 35649 13587 35683
rect 13737 35649 13771 35683
rect 15761 35649 15795 35683
rect 16865 35649 16899 35683
rect 17132 35649 17166 35683
rect 18705 35649 18739 35683
rect 18972 35649 19006 35683
rect 20913 35649 20947 35683
rect 21005 35649 21039 35683
rect 21097 35649 21131 35683
rect 21833 35649 21867 35683
rect 22744 35649 22778 35683
rect 24409 35649 24443 35683
rect 24676 35649 24710 35683
rect 26433 35649 26467 35683
rect 27169 35649 27203 35683
rect 27445 35649 27479 35683
rect 27629 35649 27663 35683
rect 28181 35649 28215 35683
rect 29009 35649 29043 35683
rect 29285 35649 29319 35683
rect 29469 35649 29503 35683
rect 9505 35581 9539 35615
rect 9781 35581 9815 35615
rect 11529 35581 11563 35615
rect 13829 35581 13863 35615
rect 15945 35581 15979 35615
rect 22477 35581 22511 35615
rect 29929 35581 29963 35615
rect 10885 35513 10919 35547
rect 21925 35513 21959 35547
rect 23857 35513 23891 35547
rect 26249 35513 26283 35547
rect 4721 35445 4755 35479
rect 9045 35445 9079 35479
rect 12909 35445 12943 35479
rect 14749 35445 14783 35479
rect 15393 35445 15427 35479
rect 18245 35445 18279 35479
rect 20085 35445 20119 35479
rect 21281 35445 21315 35479
rect 25789 35445 25823 35479
rect 26985 35445 27019 35479
rect 28273 35445 28307 35479
rect 28825 35445 28859 35479
rect 31309 35445 31343 35479
rect 1869 35241 1903 35275
rect 2237 35241 2271 35275
rect 3157 35241 3191 35275
rect 6469 35241 6503 35275
rect 8953 35241 8987 35275
rect 12081 35241 12115 35275
rect 14933 35241 14967 35275
rect 15577 35241 15611 35275
rect 17141 35241 17175 35275
rect 17601 35241 17635 35275
rect 18061 35241 18095 35275
rect 19257 35241 19291 35275
rect 23029 35241 23063 35275
rect 24961 35241 24995 35275
rect 26065 35241 26099 35275
rect 26433 35241 26467 35275
rect 29009 35241 29043 35275
rect 5181 35173 5215 35207
rect 9321 35173 9355 35207
rect 11713 35173 11747 35207
rect 13553 35173 13587 35207
rect 17417 35173 17451 35207
rect 2329 35105 2363 35139
rect 3801 35105 3835 35139
rect 9413 35105 9447 35139
rect 14565 35105 14599 35139
rect 2053 35037 2087 35071
rect 2973 35037 3007 35071
rect 3249 35037 3283 35071
rect 6653 35037 6687 35071
rect 6929 35037 6963 35071
rect 7113 35037 7147 35071
rect 7757 35037 7791 35071
rect 8033 35037 8067 35071
rect 8217 35037 8251 35071
rect 9137 35037 9171 35071
rect 9873 35037 9907 35071
rect 14749 35037 14783 35071
rect 15393 35037 15427 35071
rect 16589 35037 16623 35071
rect 16773 35037 16807 35071
rect 16957 35037 16991 35071
rect 17785 35037 17819 35071
rect 4046 34969 4080 35003
rect 10140 34969 10174 35003
rect 13369 34969 13403 35003
rect 16865 34969 16899 35003
rect 17417 34969 17451 35003
rect 19625 35173 19659 35207
rect 23397 35173 23431 35207
rect 29101 35173 29135 35207
rect 21925 35105 21959 35139
rect 30297 35105 30331 35139
rect 18705 35037 18739 35071
rect 19441 35037 19475 35071
rect 19717 35037 19751 35071
rect 20177 35037 20211 35071
rect 20821 35037 20855 35071
rect 21189 35037 21223 35071
rect 21557 35037 21591 35071
rect 22109 35037 22143 35071
rect 23213 35037 23247 35071
rect 23489 35037 23523 35071
rect 25145 35037 25179 35071
rect 25421 35037 25455 35071
rect 25605 35037 25639 35071
rect 26249 35037 26283 35071
rect 26525 35037 26559 35071
rect 27169 35037 27203 35071
rect 27629 35037 27663 35071
rect 29101 35037 29135 35071
rect 29837 35037 29871 35071
rect 30481 35037 30515 35071
rect 30757 35037 30791 35071
rect 30941 35037 30975 35071
rect 18061 34969 18095 35003
rect 27874 34969 27908 35003
rect 29653 34969 29687 35003
rect 2789 34901 2823 34935
rect 7573 34901 7607 34935
rect 11253 34901 11287 34935
rect 12081 34901 12115 34935
rect 12265 34901 12299 34935
rect 18521 34901 18555 34935
rect 20269 34901 20303 34935
rect 26985 34901 27019 34935
rect 3709 34697 3743 34731
rect 5181 34697 5215 34731
rect 5641 34697 5675 34731
rect 7757 34697 7791 34731
rect 8401 34697 8435 34731
rect 11805 34697 11839 34731
rect 11897 34697 11931 34731
rect 14197 34697 14231 34731
rect 14749 34697 14783 34731
rect 17417 34697 17451 34731
rect 18429 34697 18463 34731
rect 22109 34697 22143 34731
rect 1409 34561 1443 34595
rect 3065 34561 3099 34595
rect 4046 34629 4080 34663
rect 6622 34629 6656 34663
rect 8309 34629 8343 34663
rect 11713 34629 11747 34663
rect 12081 34629 12115 34663
rect 19533 34629 19567 34663
rect 22661 34629 22695 34663
rect 25973 34629 26007 34663
rect 5825 34561 5859 34595
rect 8953 34561 8987 34595
rect 9220 34561 9254 34595
rect 13185 34561 13219 34595
rect 14013 34561 14047 34595
rect 14197 34561 14231 34595
rect 14657 34561 14691 34595
rect 14841 34561 14875 34595
rect 15485 34561 15519 34595
rect 16773 34561 16807 34595
rect 17601 34561 17635 34595
rect 18245 34561 18279 34595
rect 18521 34561 18555 34595
rect 22293 34561 22327 34595
rect 3341 34493 3375 34527
rect 3709 34493 3743 34527
rect 3801 34493 3835 34527
rect 6377 34493 6411 34527
rect 11529 34493 11563 34527
rect 13369 34493 13403 34527
rect 13461 34493 13495 34527
rect 15669 34493 15703 34527
rect 15761 34493 15795 34527
rect 22937 34561 22971 34595
rect 23121 34561 23155 34595
rect 23673 34561 23707 34595
rect 24869 34561 24903 34595
rect 25145 34561 25179 34595
rect 25329 34561 25363 34595
rect 26157 34561 26191 34595
rect 27445 34561 27479 34595
rect 28365 34561 28399 34595
rect 28549 34561 28583 34595
rect 29469 34561 29503 34595
rect 30665 34561 30699 34595
rect 30941 34561 30975 34595
rect 31125 34561 31159 34595
rect 23213 34493 23247 34527
rect 26341 34493 26375 34527
rect 26433 34493 26467 34527
rect 27169 34493 27203 34527
rect 13001 34425 13035 34459
rect 16957 34425 16991 34459
rect 22661 34425 22695 34459
rect 29193 34493 29227 34527
rect 30481 34493 30515 34527
rect 28365 34425 28399 34459
rect 28733 34425 28767 34459
rect 1593 34357 1627 34391
rect 2881 34357 2915 34391
rect 3249 34357 3283 34391
rect 10333 34357 10367 34391
rect 15301 34357 15335 34391
rect 18245 34357 18279 34391
rect 20821 34357 20855 34391
rect 22753 34357 22787 34391
rect 23765 34357 23799 34391
rect 24685 34357 24719 34391
rect 1869 34153 1903 34187
rect 2237 34153 2271 34187
rect 5917 34153 5951 34187
rect 8953 34153 8987 34187
rect 10057 34153 10091 34187
rect 11713 34153 11747 34187
rect 14657 34153 14691 34187
rect 15209 34153 15243 34187
rect 18613 34153 18647 34187
rect 20729 34153 20763 34187
rect 23489 34153 23523 34187
rect 25789 34153 25823 34187
rect 31033 34153 31067 34187
rect 17693 34085 17727 34119
rect 21557 34085 21591 34119
rect 28549 34085 28583 34119
rect 28917 34085 28951 34119
rect 2329 34017 2363 34051
rect 3157 34017 3191 34051
rect 6929 34017 6963 34051
rect 10425 34017 10459 34051
rect 14749 34017 14783 34051
rect 16313 34017 16347 34051
rect 18705 34017 18739 34051
rect 21649 34017 21683 34051
rect 26341 34017 26375 34051
rect 2053 33949 2087 33983
rect 2973 33949 3007 33983
rect 3249 33949 3283 33983
rect 4537 33949 4571 33983
rect 9137 33949 9171 33983
rect 9413 33949 9447 33983
rect 9597 33949 9631 33983
rect 10241 33949 10275 33983
rect 10517 33949 10551 33983
rect 11069 33949 11103 33983
rect 11161 33949 11195 33983
rect 11897 33949 11931 33983
rect 11989 33949 12023 33983
rect 13001 33949 13035 33983
rect 14473 33949 14507 33983
rect 15393 33949 15427 33983
rect 15669 33949 15703 33983
rect 15853 33949 15887 33983
rect 16497 33949 16531 33983
rect 18429 33949 18463 33983
rect 19349 33949 19383 33983
rect 21373 33949 21407 33983
rect 22109 33949 22143 33983
rect 22376 33949 22410 33983
rect 24409 33949 24443 33983
rect 26597 33949 26631 33983
rect 28733 33949 28767 33983
rect 29009 33949 29043 33983
rect 29745 33949 29779 33983
rect 30021 33949 30055 33983
rect 30205 33949 30239 33983
rect 30849 33949 30883 33983
rect 31125 33949 31159 33983
rect 4782 33881 4816 33915
rect 7196 33881 7230 33915
rect 11713 33881 11747 33915
rect 13185 33881 13219 33915
rect 17509 33881 17543 33915
rect 19616 33881 19650 33915
rect 21189 33881 21223 33915
rect 24676 33881 24710 33915
rect 2789 33813 2823 33847
rect 8309 33813 8343 33847
rect 14289 33813 14323 33847
rect 16681 33813 16715 33847
rect 18245 33813 18279 33847
rect 27721 33813 27755 33847
rect 29561 33813 29595 33847
rect 30665 33813 30699 33847
rect 5089 33609 5123 33643
rect 7573 33609 7607 33643
rect 8769 33609 8803 33643
rect 12817 33609 12851 33643
rect 15393 33609 15427 33643
rect 15761 33609 15795 33643
rect 20085 33609 20119 33643
rect 21925 33609 21959 33643
rect 24593 33609 24627 33643
rect 25713 33609 25747 33643
rect 29653 33609 29687 33643
rect 30297 33609 30331 33643
rect 7021 33541 7055 33575
rect 11529 33541 11563 33575
rect 13452 33541 13486 33575
rect 20729 33541 20763 33575
rect 22201 33541 22235 33575
rect 23719 33541 23753 33575
rect 25513 33541 25547 33575
rect 1409 33473 1443 33507
rect 1676 33473 1710 33507
rect 3249 33473 3283 33507
rect 3505 33473 3539 33507
rect 5273 33473 5307 33507
rect 5549 33473 5583 33507
rect 5733 33473 5767 33507
rect 6837 33473 6871 33507
rect 7113 33473 7147 33507
rect 7757 33473 7791 33507
rect 8033 33473 8067 33507
rect 8953 33473 8987 33507
rect 9229 33473 9263 33507
rect 9413 33473 9447 33507
rect 10333 33473 10367 33507
rect 10977 33473 11011 33507
rect 11713 33473 11747 33507
rect 11805 33473 11839 33507
rect 12541 33473 12575 33507
rect 12725 33473 12759 33507
rect 12817 33473 12851 33507
rect 15853 33473 15887 33507
rect 16865 33473 16899 33507
rect 17132 33473 17166 33507
rect 18705 33473 18739 33507
rect 18961 33473 18995 33507
rect 20545 33473 20579 33507
rect 20821 33473 20855 33507
rect 21833 33473 21867 33507
rect 22845 33473 22879 33507
rect 23305 33473 23339 33507
rect 24777 33473 24811 33507
rect 25053 33473 25087 33507
rect 27169 33473 27203 33507
rect 27445 33473 27479 33507
rect 27629 33473 27663 33507
rect 28273 33473 28307 33507
rect 28540 33473 28574 33507
rect 30481 33473 30515 33507
rect 30757 33473 30791 33507
rect 30941 33473 30975 33507
rect 7941 33405 7975 33439
rect 13185 33405 13219 33439
rect 15945 33405 15979 33439
rect 11529 33337 11563 33371
rect 20545 33337 20579 33371
rect 24961 33337 24995 33371
rect 25881 33337 25915 33371
rect 2789 33269 2823 33303
rect 4629 33269 4663 33303
rect 6653 33269 6687 33303
rect 10149 33269 10183 33303
rect 10793 33269 10827 33303
rect 12541 33269 12575 33303
rect 14565 33269 14599 33303
rect 18245 33269 18279 33303
rect 22017 33269 22051 33303
rect 22109 33269 22143 33303
rect 22661 33269 22695 33303
rect 23673 33269 23707 33303
rect 23857 33269 23891 33303
rect 25697 33269 25731 33303
rect 26985 33269 27019 33303
rect 1685 33065 1719 33099
rect 3341 33065 3375 33099
rect 9137 33065 9171 33099
rect 13461 33065 13495 33099
rect 14473 33065 14507 33099
rect 16497 33065 16531 33099
rect 17417 33065 17451 33099
rect 22845 33065 22879 33099
rect 23213 33065 23247 33099
rect 25697 33065 25731 33099
rect 28549 33065 28583 33099
rect 31309 33065 31343 33099
rect 2053 32997 2087 33031
rect 3801 32997 3835 33031
rect 5549 32997 5583 33031
rect 10333 32997 10367 33031
rect 18613 32997 18647 33031
rect 22017 32997 22051 33031
rect 1869 32861 1903 32895
rect 2145 32861 2179 32895
rect 2789 32861 2823 32895
rect 3065 32861 3099 32895
rect 3249 32861 3283 32895
rect 3341 32861 3375 32895
rect 3985 32861 4019 32895
rect 4445 32861 4479 32895
rect 4721 32861 4755 32895
rect 6193 32929 6227 32963
rect 10425 32929 10459 32963
rect 15117 32929 15151 32963
rect 20637 32929 20671 32963
rect 22477 32929 22511 32963
rect 5917 32861 5951 32895
rect 6101 32861 6135 32895
rect 6745 32861 6779 32895
rect 7021 32861 7055 32895
rect 7113 32861 7147 32895
rect 7941 32861 7975 32895
rect 8217 32861 8251 32895
rect 10149 32861 10183 32895
rect 10885 32861 10919 32895
rect 12725 32861 12759 32895
rect 13369 32861 13403 32895
rect 14289 32861 14323 32895
rect 14565 32861 14599 32895
rect 15384 32861 15418 32895
rect 18521 32861 18555 32895
rect 18705 32861 18739 32895
rect 19349 32861 19383 32895
rect 19993 32861 20027 32895
rect 22661 32861 22695 32895
rect 28917 32997 28951 33031
rect 23581 32929 23615 32963
rect 23673 32929 23707 32963
rect 25237 32929 25271 32963
rect 26617 32929 26651 32963
rect 29929 32929 29963 32963
rect 23489 32861 23523 32895
rect 23765 32861 23799 32895
rect 24961 32861 24995 32895
rect 25145 32861 25179 32895
rect 25881 32861 25915 32895
rect 26065 32861 26099 32895
rect 26157 32861 26191 32895
rect 26801 32861 26835 32895
rect 27077 32861 27111 32895
rect 27261 32861 27295 32895
rect 28733 32861 28767 32895
rect 29009 32861 29043 32895
rect 30196 32861 30230 32895
rect 2605 32793 2639 32827
rect 5457 32793 5491 32827
rect 6929 32793 6963 32827
rect 8953 32793 8987 32827
rect 9169 32793 9203 32827
rect 9965 32793 9999 32827
rect 11130 32793 11164 32827
rect 17693 32793 17727 32827
rect 17969 32793 18003 32827
rect 20904 32793 20938 32827
rect 23213 32793 23247 32827
rect 27905 32793 27939 32827
rect 5733 32725 5767 32759
rect 7297 32725 7331 32759
rect 7757 32725 7791 32759
rect 8125 32725 8159 32759
rect 9321 32725 9355 32759
rect 12265 32725 12299 32759
rect 12817 32725 12851 32759
rect 14105 32725 14139 32759
rect 17877 32725 17911 32759
rect 19441 32725 19475 32759
rect 20085 32725 20119 32759
rect 23305 32725 23339 32759
rect 24777 32725 24811 32759
rect 27997 32725 28031 32759
rect 5825 32521 5859 32555
rect 6377 32521 6411 32555
rect 8677 32521 8711 32555
rect 11897 32521 11931 32555
rect 14473 32521 14507 32555
rect 16129 32521 16163 32555
rect 16681 32521 16715 32555
rect 17877 32521 17911 32555
rect 20453 32521 20487 32555
rect 31309 32521 31343 32555
rect 4712 32453 4746 32487
rect 7665 32453 7699 32487
rect 7849 32453 7883 32487
rect 8769 32453 8803 32487
rect 12541 32453 12575 32487
rect 12900 32453 12934 32487
rect 21189 32453 21223 32487
rect 22017 32453 22051 32487
rect 22836 32453 22870 32487
rect 1409 32385 1443 32419
rect 1676 32385 1710 32419
rect 3433 32385 3467 32419
rect 3709 32385 3743 32419
rect 3893 32385 3927 32419
rect 4445 32385 4479 32419
rect 6561 32385 6595 32419
rect 6837 32385 6871 32419
rect 7021 32385 7055 32419
rect 8585 32385 8619 32419
rect 9505 32385 9539 32419
rect 9761 32385 9795 32419
rect 9045 32317 9079 32351
rect 2789 32249 2823 32283
rect 8309 32249 8343 32283
rect 11529 32249 11563 32283
rect 14657 32385 14691 32419
rect 14933 32385 14967 32419
rect 15117 32385 15151 32419
rect 15945 32385 15979 32419
rect 17049 32385 17083 32419
rect 18061 32385 18095 32419
rect 18337 32385 18371 32419
rect 19349 32385 19383 32419
rect 19625 32385 19659 32419
rect 20361 32385 20395 32419
rect 21005 32385 21039 32419
rect 21281 32385 21315 32419
rect 21649 32385 21683 32419
rect 21833 32385 21867 32419
rect 22109 32385 22143 32419
rect 22569 32385 22603 32419
rect 24409 32385 24443 32419
rect 24676 32385 24710 32419
rect 26433 32385 26467 32419
rect 27169 32385 27203 32419
rect 28227 32385 28261 32419
rect 29469 32385 29503 32419
rect 12633 32317 12667 32351
rect 15761 32317 15795 32351
rect 17141 32317 17175 32351
rect 17233 32317 17267 32351
rect 14013 32249 14047 32283
rect 18245 32249 18279 32283
rect 19533 32249 19567 32283
rect 22201 32317 22235 32351
rect 27353 32317 27387 32351
rect 28089 32317 28123 32351
rect 28365 32317 28399 32351
rect 29653 32317 29687 32351
rect 30389 32317 30423 32351
rect 30506 32317 30540 32351
rect 30665 32317 30699 32351
rect 21833 32249 21867 32283
rect 3249 32181 3283 32215
rect 8953 32181 8987 32215
rect 10885 32181 10919 32215
rect 11897 32181 11931 32215
rect 12081 32181 12115 32215
rect 12541 32181 12575 32215
rect 19165 32181 19199 32215
rect 21005 32181 21039 32215
rect 21649 32181 21683 32215
rect 23949 32249 23983 32283
rect 27813 32249 27847 32283
rect 30113 32249 30147 32283
rect 22201 32181 22235 32215
rect 25789 32181 25823 32215
rect 26249 32181 26283 32215
rect 29009 32181 29043 32215
rect 2421 31977 2455 32011
rect 3801 31977 3835 32011
rect 7573 31977 7607 32011
rect 9597 31977 9631 32011
rect 10885 31977 10919 32011
rect 13461 31977 13495 32011
rect 21005 31977 21039 32011
rect 23213 31977 23247 32011
rect 25421 31977 25455 32011
rect 27905 31977 27939 32011
rect 28549 31977 28583 32011
rect 2789 31909 2823 31943
rect 7113 31909 7147 31943
rect 9045 31909 9079 31943
rect 4997 31841 5031 31875
rect 5273 31841 5307 31875
rect 7849 31841 7883 31875
rect 8033 31841 8067 31875
rect 9229 31841 9263 31875
rect 10701 31841 10735 31875
rect 12449 31909 12483 31943
rect 12541 31909 12575 31943
rect 14197 31909 14231 31943
rect 17233 31909 17267 31943
rect 18429 31909 18463 31943
rect 12173 31841 12207 31875
rect 15853 31841 15887 31875
rect 16773 31841 16807 31875
rect 17785 31841 17819 31875
rect 1961 31773 1995 31807
rect 2605 31773 2639 31807
rect 2881 31773 2915 31807
rect 3985 31773 4019 31807
rect 4261 31773 4295 31807
rect 4445 31773 4479 31807
rect 6469 31773 6503 31807
rect 6562 31773 6596 31807
rect 6745 31773 6779 31807
rect 6837 31773 6871 31807
rect 6975 31773 7009 31807
rect 7757 31773 7791 31807
rect 7941 31773 7975 31807
rect 8217 31773 8251 31807
rect 9505 31773 9539 31807
rect 9781 31773 9815 31807
rect 10333 31773 10367 31807
rect 10517 31773 10551 31807
rect 10885 31773 10919 31807
rect 11345 31773 11379 31807
rect 11621 31773 11655 31807
rect 12357 31773 12391 31807
rect 12632 31773 12666 31807
rect 12829 31773 12863 31807
rect 13369 31773 13403 31807
rect 14381 31773 14415 31807
rect 14657 31773 14691 31807
rect 14841 31773 14875 31807
rect 15669 31773 15703 31807
rect 15945 31773 15979 31807
rect 16589 31773 16623 31807
rect 18429 31773 18463 31807
rect 18705 31773 18739 31807
rect 19257 31773 19291 31807
rect 19524 31773 19558 31807
rect 1777 31705 1811 31739
rect 9321 31705 9355 31739
rect 22201 31909 22235 31943
rect 24869 31909 24903 31943
rect 30481 31909 30515 31943
rect 21097 31841 21131 31875
rect 22477 31841 22511 31875
rect 22661 31841 22695 31875
rect 26525 31841 26559 31875
rect 29009 31841 29043 31875
rect 30573 31841 30607 31875
rect 21373 31773 21407 31807
rect 21465 31773 21499 31807
rect 21557 31773 21591 31807
rect 21741 31773 21775 31807
rect 22385 31773 22419 31807
rect 22560 31773 22594 31807
rect 23213 31773 23247 31807
rect 23489 31773 23523 31807
rect 24777 31773 24811 31807
rect 25605 31773 25639 31807
rect 25881 31773 25915 31807
rect 26065 31773 26099 31807
rect 26792 31773 26826 31807
rect 28733 31773 28767 31807
rect 28917 31773 28951 31807
rect 30297 31773 30331 31807
rect 31125 31773 31159 31807
rect 11437 31637 11471 31671
rect 15485 31637 15519 31671
rect 17601 31637 17635 31671
rect 17693 31637 17727 31671
rect 18613 31637 18647 31671
rect 20637 31637 20671 31671
rect 21005 31637 21039 31671
rect 23397 31637 23431 31671
rect 30113 31637 30147 31671
rect 31217 31637 31251 31671
rect 7297 31433 7331 31467
rect 8309 31433 8343 31467
rect 9965 31433 9999 31467
rect 13277 31433 13311 31467
rect 14289 31433 14323 31467
rect 15301 31433 15335 31467
rect 17233 31433 17267 31467
rect 6745 31365 6779 31399
rect 7113 31365 7147 31399
rect 8125 31365 8159 31399
rect 9321 31365 9355 31399
rect 11989 31365 12023 31399
rect 13093 31365 13127 31399
rect 2605 31297 2639 31331
rect 3893 31297 3927 31331
rect 4537 31297 4571 31331
rect 5825 31297 5859 31331
rect 6929 31297 6963 31331
rect 7021 31297 7055 31331
rect 2881 31229 2915 31263
rect 4813 31229 4847 31263
rect 2789 31161 2823 31195
rect 4721 31161 4755 31195
rect 8309 31297 8343 31331
rect 8585 31297 8619 31331
rect 9781 31297 9815 31331
rect 10609 31297 10643 31331
rect 10885 31297 10919 31331
rect 14473 31297 14507 31331
rect 15485 31297 15519 31331
rect 15761 31297 15795 31331
rect 15945 31297 15979 31331
rect 16865 31297 16899 31331
rect 8677 31229 8711 31263
rect 9689 31229 9723 31263
rect 14105 31229 14139 31263
rect 17141 31229 17175 31263
rect 18429 31433 18463 31467
rect 18981 31433 19015 31467
rect 20913 31433 20947 31467
rect 21833 31433 21867 31467
rect 24317 31433 24351 31467
rect 28365 31433 28399 31467
rect 31309 31433 31343 31467
rect 20729 31365 20763 31399
rect 17601 31297 17635 31331
rect 17785 31297 17819 31331
rect 18061 31297 18095 31331
rect 18245 31297 18279 31331
rect 18429 31297 18463 31331
rect 19165 31297 19199 31331
rect 19441 31297 19475 31331
rect 19625 31297 19659 31331
rect 20545 31297 20579 31331
rect 22017 31297 22051 31331
rect 22293 31297 22327 31331
rect 23489 31297 23523 31331
rect 24133 31297 24167 31331
rect 25237 31297 25271 31331
rect 26065 31297 26099 31331
rect 26985 31297 27019 31331
rect 28549 31297 28583 31331
rect 28825 31297 28859 31331
rect 29469 31297 29503 31331
rect 30196 31297 30230 31331
rect 23305 31229 23339 31263
rect 25513 31229 25547 31263
rect 27261 31229 27295 31263
rect 28733 31229 28767 31263
rect 29929 31229 29963 31263
rect 12725 31161 12759 31195
rect 17233 31161 17267 31195
rect 25421 31161 25455 31195
rect 26249 31161 26283 31195
rect 2421 31093 2455 31127
rect 3709 31093 3743 31127
rect 4353 31093 4387 31127
rect 5641 31093 5675 31127
rect 8125 31093 8159 31127
rect 9413 31093 9447 31127
rect 10425 31093 10459 31127
rect 10793 31093 10827 31127
rect 12081 31093 12115 31127
rect 13093 31093 13127 31127
rect 14473 31093 14507 31127
rect 16681 31093 16715 31127
rect 17049 31093 17083 31127
rect 22201 31093 22235 31127
rect 23673 31093 23707 31127
rect 25053 31093 25087 31127
rect 29285 31093 29319 31127
rect 4261 30889 4295 30923
rect 6745 30889 6779 30923
rect 7849 30889 7883 30923
rect 9229 30889 9263 30923
rect 11161 30889 11195 30923
rect 12909 30889 12943 30923
rect 14105 30889 14139 30923
rect 16589 30889 16623 30923
rect 19257 30889 19291 30923
rect 23581 30889 23615 30923
rect 26249 30889 26283 30923
rect 30665 30889 30699 30923
rect 2881 30821 2915 30855
rect 6193 30821 6227 30855
rect 12449 30821 12483 30855
rect 13461 30821 13495 30855
rect 14565 30821 14599 30855
rect 21741 30821 21775 30855
rect 11989 30753 12023 30787
rect 1501 30685 1535 30719
rect 1768 30685 1802 30719
rect 4445 30685 4479 30719
rect 4721 30685 4755 30719
rect 4905 30685 4939 30719
rect 5733 30685 5767 30719
rect 7389 30685 7423 30719
rect 8033 30685 8067 30719
rect 8125 30685 8159 30719
rect 8309 30685 8343 30719
rect 8401 30685 8435 30719
rect 9137 30685 9171 30719
rect 9781 30685 9815 30719
rect 10048 30685 10082 30719
rect 11897 30685 11931 30719
rect 12081 30685 12115 30719
rect 6469 30617 6503 30651
rect 14749 30753 14783 30787
rect 20361 30753 20395 30787
rect 22201 30753 22235 30787
rect 29561 30753 29595 30787
rect 12725 30685 12759 30719
rect 13369 30685 13403 30719
rect 14289 30685 14323 30719
rect 14381 30685 14415 30719
rect 14657 30685 14691 30719
rect 12541 30617 12575 30651
rect 5549 30549 5583 30583
rect 6377 30549 6411 30583
rect 6561 30549 6595 30583
rect 7205 30549 7239 30583
rect 12449 30549 12483 30583
rect 15209 30685 15243 30719
rect 15476 30685 15510 30719
rect 17049 30685 17083 30719
rect 19441 30685 19475 30719
rect 19717 30685 19751 30719
rect 19901 30685 19935 30719
rect 24409 30685 24443 30719
rect 24676 30685 24710 30719
rect 26433 30685 26467 30719
rect 26709 30685 26743 30719
rect 26893 30685 26927 30719
rect 27905 30685 27939 30719
rect 28733 30685 28767 30719
rect 28917 30685 28951 30719
rect 29009 30685 29043 30719
rect 29745 30685 29779 30719
rect 30021 30685 30055 30719
rect 30205 30685 30239 30719
rect 30849 30685 30883 30719
rect 31125 30685 31159 30719
rect 31309 30685 31343 30719
rect 17294 30617 17328 30651
rect 20628 30617 20662 30651
rect 22446 30617 22480 30651
rect 28089 30617 28123 30651
rect 14749 30549 14783 30583
rect 18429 30549 18463 30583
rect 25789 30549 25823 30583
rect 28549 30549 28583 30583
rect 1869 30345 1903 30379
rect 8585 30345 8619 30379
rect 9321 30345 9355 30379
rect 14841 30345 14875 30379
rect 17509 30345 17543 30379
rect 20085 30345 20119 30379
rect 20637 30345 20671 30379
rect 22109 30345 22143 30379
rect 4506 30277 4540 30311
rect 11529 30277 11563 30311
rect 13553 30277 13587 30311
rect 16773 30277 16807 30311
rect 17417 30277 17451 30311
rect 23121 30277 23155 30311
rect 28273 30277 28307 30311
rect 2053 30209 2087 30243
rect 2329 30209 2363 30243
rect 2513 30209 2547 30243
rect 3157 30209 3191 30243
rect 3433 30209 3467 30243
rect 3617 30209 3651 30243
rect 7021 30209 7055 30243
rect 7205 30209 7239 30243
rect 7389 30209 7423 30243
rect 8401 30209 8435 30243
rect 8493 30209 8527 30243
rect 9505 30209 9539 30243
rect 11713 30209 11747 30243
rect 12541 30209 12575 30243
rect 12725 30209 12759 30243
rect 15853 30209 15887 30243
rect 4261 30141 4295 30175
rect 7297 30141 7331 30175
rect 9965 30141 9999 30175
rect 10241 30141 10275 30175
rect 11989 30141 12023 30175
rect 8217 30073 8251 30107
rect 16957 30073 16991 30107
rect 17693 30209 17727 30243
rect 17969 30209 18003 30243
rect 18153 30209 18187 30243
rect 18889 30209 18923 30243
rect 19809 30209 19843 30243
rect 19901 30209 19935 30243
rect 20821 30209 20855 30243
rect 22293 30209 22327 30243
rect 22477 30209 22511 30243
rect 23029 30209 23063 30243
rect 23673 30209 23707 30243
rect 25053 30209 25087 30243
rect 25789 30209 25823 30243
rect 25973 30209 26007 30243
rect 26249 30209 26283 30243
rect 26433 30209 26467 30243
rect 27261 30209 27295 30243
rect 30665 30209 30699 30243
rect 30941 30209 30975 30243
rect 31125 30209 31159 30243
rect 18245 30141 18279 30175
rect 18613 30141 18647 30175
rect 21097 30141 21131 30175
rect 22569 30141 22603 30175
rect 23857 30141 23891 30175
rect 25329 30141 25363 30175
rect 26985 30141 27019 30175
rect 18429 30073 18463 30107
rect 19809 30073 19843 30107
rect 24869 30073 24903 30107
rect 30481 30073 30515 30107
rect 2973 30005 3007 30039
rect 5641 30005 5675 30039
rect 8769 30005 8803 30039
rect 11897 30005 11931 30039
rect 15945 30005 15979 30039
rect 17417 30005 17451 30039
rect 21005 30005 21039 30039
rect 25237 30005 25271 30039
rect 29561 30005 29595 30039
rect 2789 29801 2823 29835
rect 6469 29801 6503 29835
rect 6653 29801 6687 29835
rect 13553 29801 13587 29835
rect 19993 29801 20027 29835
rect 20821 29801 20855 29835
rect 24961 29801 24995 29835
rect 31309 29801 31343 29835
rect 11713 29733 11747 29767
rect 14565 29733 14599 29767
rect 16681 29733 16715 29767
rect 17141 29733 17175 29767
rect 23213 29733 23247 29767
rect 5181 29665 5215 29699
rect 7389 29665 7423 29699
rect 9229 29665 9263 29699
rect 9597 29665 9631 29699
rect 21833 29665 21867 29699
rect 25513 29665 25547 29699
rect 25697 29665 25731 29699
rect 25881 29665 25915 29699
rect 26525 29665 26559 29699
rect 29929 29665 29963 29699
rect 1409 29597 1443 29631
rect 3985 29597 4019 29631
rect 4261 29597 4295 29631
rect 4445 29597 4479 29631
rect 4905 29597 4939 29631
rect 7113 29597 7147 29631
rect 9125 29597 9159 29631
rect 10333 29597 10367 29631
rect 12173 29597 12207 29631
rect 14381 29597 14415 29631
rect 14657 29597 14691 29631
rect 15393 29597 15427 29631
rect 15669 29597 15703 29631
rect 16957 29597 16991 29631
rect 17141 29597 17175 29631
rect 17693 29597 17727 29631
rect 17969 29597 18003 29631
rect 18153 29597 18187 29631
rect 21005 29597 21039 29631
rect 21097 29597 21131 29631
rect 23673 29597 23707 29631
rect 25789 29597 25823 29631
rect 25973 29597 26007 29631
rect 28733 29597 28767 29631
rect 28917 29597 28951 29631
rect 29009 29597 29043 29631
rect 30185 29597 30219 29631
rect 1676 29529 1710 29563
rect 6285 29529 6319 29563
rect 8953 29529 8987 29563
rect 10600 29529 10634 29563
rect 12440 29529 12474 29563
rect 14197 29529 14231 29563
rect 16681 29529 16715 29563
rect 19901 29529 19935 29563
rect 20821 29529 20855 29563
rect 22078 29529 22112 29563
rect 24869 29529 24903 29563
rect 26770 29529 26804 29563
rect 3801 29461 3835 29495
rect 6485 29461 6519 29495
rect 9321 29461 9355 29495
rect 9505 29461 9539 29495
rect 16865 29461 16899 29495
rect 17509 29461 17543 29495
rect 23765 29461 23799 29495
rect 27905 29461 27939 29495
rect 28549 29461 28583 29495
rect 1685 29257 1719 29291
rect 5825 29257 5859 29291
rect 7113 29257 7147 29291
rect 10701 29257 10735 29291
rect 13001 29257 13035 29291
rect 21097 29257 21131 29291
rect 21833 29257 21867 29291
rect 22477 29257 22511 29291
rect 28549 29257 28583 29291
rect 1593 29189 1627 29223
rect 6653 29189 6687 29223
rect 2421 29121 2455 29155
rect 3157 29121 3191 29155
rect 3341 29121 3375 29155
rect 3617 29121 3651 29155
rect 3801 29121 3835 29155
rect 4445 29121 4479 29155
rect 4701 29121 4735 29155
rect 6929 29121 6963 29155
rect 7297 29121 7331 29155
rect 7941 29121 7975 29155
rect 8033 29121 8067 29155
rect 8217 29121 8251 29155
rect 8319 29121 8353 29155
rect 9321 29121 9355 29155
rect 9588 29121 9622 29155
rect 11529 29121 11563 29155
rect 13185 29121 13219 29155
rect 13461 29121 13495 29155
rect 14197 29121 14231 29155
rect 14933 29121 14967 29155
rect 15117 29121 15151 29155
rect 15393 29121 15427 29155
rect 15577 29121 15611 29155
rect 17141 29121 17175 29155
rect 17325 29121 17359 29155
rect 18613 29121 18647 29155
rect 21005 29121 21039 29155
rect 22017 29121 22051 29155
rect 22201 29121 22235 29155
rect 2697 29053 2731 29087
rect 6837 29053 6871 29087
rect 7205 29053 7239 29087
rect 11805 29053 11839 29087
rect 14381 29053 14415 29087
rect 14473 29053 14507 29087
rect 17509 29053 17543 29087
rect 17601 29053 17635 29087
rect 22293 29053 22327 29087
rect 2605 28985 2639 29019
rect 13369 28985 13403 29019
rect 14013 28985 14047 29019
rect 19901 28985 19935 29019
rect 25789 29189 25823 29223
rect 22753 29121 22787 29155
rect 22845 29121 22879 29155
rect 23121 29121 23155 29155
rect 24133 29121 24167 29155
rect 24409 29121 24443 29155
rect 24501 29121 24535 29155
rect 24593 29121 24627 29155
rect 24777 29121 24811 29155
rect 28365 29121 28399 29155
rect 29377 29121 29411 29155
rect 30113 29121 30147 29155
rect 30389 29121 30423 29155
rect 22937 29053 22971 29087
rect 24869 29053 24903 29087
rect 25421 29053 25455 29087
rect 27077 29053 27111 29087
rect 27353 29053 27387 29087
rect 29193 29053 29227 29087
rect 30230 29053 30264 29087
rect 23121 28985 23155 29019
rect 29837 28985 29871 29019
rect 2237 28917 2271 28951
rect 7757 28917 7791 28951
rect 22477 28917 22511 28951
rect 25789 28917 25823 28951
rect 25973 28917 26007 28951
rect 31033 28917 31067 28951
rect 4169 28713 4203 28747
rect 6929 28713 6963 28747
rect 8953 28713 8987 28747
rect 10057 28713 10091 28747
rect 11161 28713 11195 28747
rect 11529 28713 11563 28747
rect 12081 28713 12115 28747
rect 13277 28713 13311 28747
rect 15577 28713 15611 28747
rect 17877 28713 17911 28747
rect 20637 28713 20671 28747
rect 21465 28713 21499 28747
rect 21741 28713 21775 28747
rect 22661 28713 22695 28747
rect 25973 28713 26007 28747
rect 26893 28713 26927 28747
rect 29009 28713 29043 28747
rect 3249 28645 3283 28679
rect 6377 28645 6411 28679
rect 18705 28645 18739 28679
rect 4537 28577 4571 28611
rect 5365 28577 5399 28611
rect 11621 28577 11655 28611
rect 24777 28577 24811 28611
rect 27629 28577 27663 28611
rect 1869 28509 1903 28543
rect 4353 28509 4387 28543
rect 4629 28509 4663 28543
rect 5089 28509 5123 28543
rect 6561 28509 6595 28543
rect 6653 28509 6687 28543
rect 7941 28509 7975 28543
rect 8217 28509 8251 28543
rect 8401 28509 8435 28543
rect 9137 28509 9171 28543
rect 9229 28509 9263 28543
rect 9413 28509 9447 28543
rect 9505 28509 9539 28543
rect 10241 28509 10275 28543
rect 10517 28509 10551 28543
rect 10701 28509 10735 28543
rect 10793 28509 10827 28543
rect 11345 28509 11379 28543
rect 12265 28509 12299 28543
rect 12541 28509 12575 28543
rect 12725 28509 12759 28543
rect 13553 28509 13587 28543
rect 14289 28509 14323 28543
rect 14565 28509 14599 28543
rect 14749 28509 14783 28543
rect 15761 28509 15795 28543
rect 16037 28509 16071 28543
rect 16497 28509 16531 28543
rect 19257 28509 19291 28543
rect 19513 28509 19547 28543
rect 21097 28509 21131 28543
rect 21741 28509 21775 28543
rect 22937 28509 22971 28543
rect 23029 28509 23063 28543
rect 23142 28509 23176 28543
rect 23305 28509 23339 28543
rect 24409 28509 24443 28543
rect 24593 28509 24627 28543
rect 24685 28509 24719 28543
rect 24961 28509 24995 28543
rect 25605 28509 25639 28543
rect 25789 28509 25823 28543
rect 26525 28509 26559 28543
rect 29929 28509 29963 28543
rect 30185 28509 30219 28543
rect 2136 28441 2170 28475
rect 6745 28441 6779 28475
rect 13277 28441 13311 28475
rect 15945 28441 15979 28475
rect 16764 28441 16798 28475
rect 18521 28441 18555 28475
rect 21465 28441 21499 28475
rect 22385 28441 22419 28475
rect 27896 28441 27930 28475
rect 7757 28373 7791 28407
rect 10793 28373 10827 28407
rect 13461 28373 13495 28407
rect 14105 28373 14139 28407
rect 21649 28373 21683 28407
rect 22569 28373 22603 28407
rect 25145 28373 25179 28407
rect 26893 28373 26927 28407
rect 27077 28373 27111 28407
rect 31309 28373 31343 28407
rect 9689 28169 9723 28203
rect 14933 28169 14967 28203
rect 16129 28169 16163 28203
rect 17233 28169 17267 28203
rect 19625 28169 19659 28203
rect 21649 28169 21683 28203
rect 2973 28101 3007 28135
rect 17509 28101 17543 28135
rect 17601 28101 17635 28135
rect 18337 28101 18371 28135
rect 18521 28101 18555 28135
rect 20637 28101 20671 28135
rect 23857 28169 23891 28203
rect 24225 28169 24259 28203
rect 24869 28169 24903 28203
rect 25881 28169 25915 28203
rect 27537 28169 27571 28203
rect 27905 28169 27939 28203
rect 28273 28169 28307 28203
rect 28825 28169 28859 28203
rect 1409 28033 1443 28067
rect 2513 28033 2547 28067
rect 5365 28033 5399 28067
rect 6644 28033 6678 28067
rect 8401 28033 8435 28067
rect 8677 28033 8711 28067
rect 8861 28033 8895 28067
rect 8953 28033 8987 28067
rect 9873 28033 9907 28067
rect 10149 28033 10183 28067
rect 10333 28033 10367 28067
rect 10793 28033 10827 28067
rect 10977 28033 11011 28067
rect 11969 28033 12003 28067
rect 13809 28033 13843 28067
rect 15393 28033 15427 28067
rect 15577 28033 15611 28067
rect 15669 28033 15703 28067
rect 15945 28033 15979 28067
rect 17417 28033 17451 28067
rect 17693 28033 17727 28067
rect 17877 28033 17911 28067
rect 18613 28033 18647 28067
rect 19717 28033 19751 28067
rect 20913 28033 20947 28067
rect 21005 28033 21039 28067
rect 21097 28033 21131 28067
rect 21281 28033 21315 28067
rect 21649 28033 21683 28067
rect 21925 28033 21959 28067
rect 22911 28033 22945 28067
rect 23213 28033 23247 28067
rect 5641 27965 5675 27999
rect 6377 27965 6411 27999
rect 5549 27897 5583 27931
rect 7757 27897 7791 27931
rect 11713 27965 11747 27999
rect 13553 27965 13587 27999
rect 15761 27965 15795 27999
rect 18409 27965 18443 27999
rect 19809 27965 19843 27999
rect 23029 27965 23063 27999
rect 23121 27965 23155 27999
rect 19257 27897 19291 27931
rect 22109 27897 22143 27931
rect 22753 27897 22787 27931
rect 24593 28033 24627 28067
rect 24685 28033 24719 28067
rect 24961 28033 24995 28067
rect 26157 28033 26191 28067
rect 26341 28033 26375 28067
rect 27169 28033 27203 28067
rect 26065 27965 26099 27999
rect 26249 27965 26283 27999
rect 27445 27965 27479 27999
rect 26985 27897 27019 27931
rect 28365 28101 28399 28135
rect 28825 28033 28859 28067
rect 29285 28033 29319 28067
rect 29561 28033 29595 28067
rect 29745 28033 29779 28067
rect 30205 28033 30239 28067
rect 30481 28033 30515 28067
rect 30757 28033 30791 28067
rect 30941 28033 30975 28067
rect 28457 27965 28491 27999
rect 1593 27829 1627 27863
rect 2329 27829 2363 27863
rect 4261 27829 4295 27863
rect 5181 27829 5215 27863
rect 8217 27829 8251 27863
rect 8953 27829 8987 27863
rect 10885 27829 10919 27863
rect 13093 27829 13127 27863
rect 23857 27829 23891 27863
rect 24501 27829 24535 27863
rect 27353 27829 27387 27863
rect 27537 27829 27571 27863
rect 29101 27829 29135 27863
rect 30205 27829 30239 27863
rect 30297 27829 30331 27863
rect 11529 27625 11563 27659
rect 16037 27625 16071 27659
rect 20913 27625 20947 27659
rect 21465 27625 21499 27659
rect 24501 27625 24535 27659
rect 26157 27625 26191 27659
rect 28549 27625 28583 27659
rect 31309 27625 31343 27659
rect 2605 27557 2639 27591
rect 2973 27557 3007 27591
rect 4353 27557 4387 27591
rect 6285 27557 6319 27591
rect 7205 27557 7239 27591
rect 9321 27557 9355 27591
rect 11897 27557 11931 27591
rect 22017 27557 22051 27591
rect 25513 27557 25547 27591
rect 28089 27557 28123 27591
rect 2053 27489 2087 27523
rect 2145 27489 2179 27523
rect 3065 27489 3099 27523
rect 4905 27489 4939 27523
rect 8493 27489 8527 27523
rect 9413 27489 9447 27523
rect 18889 27489 18923 27523
rect 23029 27489 23063 27523
rect 24685 27489 24719 27523
rect 29009 27489 29043 27523
rect 29929 27489 29963 27523
rect 1869 27421 1903 27455
rect 2789 27421 2823 27455
rect 4169 27421 4203 27455
rect 4445 27421 4479 27455
rect 5172 27421 5206 27455
rect 7021 27421 7055 27455
rect 7297 27421 7331 27455
rect 7941 27421 7975 27455
rect 8217 27421 8251 27455
rect 8401 27421 8435 27455
rect 7757 27353 7791 27387
rect 9137 27421 9171 27455
rect 9873 27421 9907 27455
rect 10149 27421 10183 27455
rect 11713 27421 11747 27455
rect 11989 27421 12023 27455
rect 12633 27421 12667 27455
rect 12909 27421 12943 27455
rect 13093 27421 13127 27455
rect 14657 27421 14691 27455
rect 14913 27421 14947 27455
rect 16589 27421 16623 27455
rect 17325 27421 17359 27455
rect 12449 27353 12483 27387
rect 17592 27353 17626 27387
rect 19533 27421 19567 27455
rect 19622 27421 19656 27455
rect 19717 27421 19751 27455
rect 19901 27421 19935 27455
rect 20729 27421 20763 27455
rect 21373 27421 21407 27455
rect 22293 27421 22327 27455
rect 22753 27421 22787 27455
rect 24409 27421 24443 27455
rect 25329 27421 25363 27455
rect 26709 27421 26743 27455
rect 28733 27421 28767 27455
rect 28917 27421 28951 27455
rect 20545 27353 20579 27387
rect 22017 27353 22051 27387
rect 26065 27353 26099 27387
rect 26954 27353 26988 27387
rect 30196 27353 30230 27387
rect 1685 27285 1719 27319
rect 3985 27285 4019 27319
rect 6837 27285 6871 27319
rect 8493 27285 8527 27319
rect 8953 27285 8987 27319
rect 16773 27285 16807 27319
rect 18705 27285 18739 27319
rect 18889 27285 18923 27319
rect 19257 27285 19291 27319
rect 22201 27285 22235 27319
rect 24685 27285 24719 27319
rect 7205 27081 7239 27115
rect 10977 27081 11011 27115
rect 11529 27081 11563 27115
rect 13553 27081 13587 27115
rect 14105 27081 14139 27115
rect 17693 27081 17727 27115
rect 18613 27081 18647 27115
rect 23213 27081 23247 27115
rect 25513 27081 25547 27115
rect 25973 27081 26007 27115
rect 30389 27081 30423 27115
rect 8392 27013 8426 27047
rect 10793 27013 10827 27047
rect 11161 27013 11195 27047
rect 12633 27013 12667 27047
rect 1676 26945 1710 26979
rect 3801 26945 3835 26979
rect 4068 26945 4102 26979
rect 5825 26945 5859 26979
rect 6561 26945 6595 26979
rect 6745 26945 6779 26979
rect 7389 26945 7423 26979
rect 7573 26945 7607 26979
rect 7665 26945 7699 26979
rect 1409 26877 1443 26911
rect 8125 26877 8159 26911
rect 10425 26877 10459 26911
rect 5181 26809 5215 26843
rect 9505 26809 9539 26843
rect 11805 26945 11839 26979
rect 11897 26945 11931 26979
rect 12010 26945 12044 26979
rect 12173 26945 12207 26979
rect 12541 26945 12575 26979
rect 12817 26945 12851 26979
rect 13737 26945 13771 26979
rect 14013 26945 14047 26979
rect 2789 26741 2823 26775
rect 5641 26741 5675 26775
rect 6561 26741 6595 26775
rect 10793 26741 10827 26775
rect 11161 26741 11195 26775
rect 20821 27013 20855 27047
rect 22078 27013 22112 27047
rect 23581 27013 23615 27047
rect 14473 26945 14507 26979
rect 14657 26945 14691 26979
rect 14749 26945 14783 26979
rect 15761 26945 15795 26979
rect 15945 26945 15979 26979
rect 16957 26945 16991 26979
rect 17877 26945 17911 26979
rect 18153 26945 18187 26979
rect 18889 26945 18923 26979
rect 19073 26945 19107 26979
rect 20085 26945 20119 26979
rect 20361 26945 20395 26979
rect 21005 26945 21039 26979
rect 21833 26945 21867 26979
rect 14105 26877 14139 26911
rect 18797 26877 18831 26911
rect 18981 26877 19015 26911
rect 21281 26877 21315 26911
rect 13001 26809 13035 26843
rect 20269 26809 20303 26843
rect 24389 26945 24423 26979
rect 26157 26945 26191 26979
rect 26985 26945 27019 26979
rect 27169 26945 27203 26979
rect 27445 26945 27479 26979
rect 27629 26945 27663 26979
rect 28273 26945 28307 26979
rect 29193 26945 29227 26979
rect 29377 26945 29411 26979
rect 30573 26945 30607 26979
rect 24133 26877 24167 26911
rect 26433 26877 26467 26911
rect 28549 26877 28583 26911
rect 29469 26877 29503 26911
rect 30849 26877 30883 26911
rect 26341 26809 26375 26843
rect 30757 26809 30791 26843
rect 12541 26741 12575 26775
rect 13921 26741 13955 26775
rect 14473 26741 14507 26775
rect 16129 26741 16163 26775
rect 17141 26741 17175 26775
rect 18061 26741 18095 26775
rect 19901 26741 19935 26775
rect 21189 26741 21223 26775
rect 23581 26741 23615 26775
rect 28089 26741 28123 26775
rect 28457 26741 28491 26775
rect 29009 26741 29043 26775
rect 4445 26537 4479 26571
rect 5549 26537 5583 26571
rect 8125 26537 8159 26571
rect 9137 26537 9171 26571
rect 11897 26537 11931 26571
rect 12817 26537 12851 26571
rect 13093 26537 13127 26571
rect 13461 26537 13495 26571
rect 21649 26537 21683 26571
rect 22845 26537 22879 26571
rect 23397 26537 23431 26571
rect 29929 26537 29963 26571
rect 30849 26537 30883 26571
rect 3065 26469 3099 26503
rect 11989 26401 12023 26435
rect 12909 26401 12943 26435
rect 2145 26333 2179 26367
rect 2421 26333 2455 26367
rect 2605 26333 2639 26367
rect 3249 26333 3283 26367
rect 3985 26333 4019 26367
rect 4629 26333 4663 26367
rect 4905 26333 4939 26367
rect 5089 26333 5123 26367
rect 5733 26333 5767 26367
rect 6009 26333 6043 26367
rect 6193 26333 6227 26367
rect 6745 26333 6779 26367
rect 7012 26333 7046 26367
rect 9689 26333 9723 26367
rect 11713 26333 11747 26367
rect 12633 26333 12667 26367
rect 18521 26469 18555 26503
rect 22569 26469 22603 26503
rect 23765 26469 23799 26503
rect 18153 26401 18187 26435
rect 13369 26333 13403 26367
rect 14657 26333 14691 26367
rect 15301 26333 15335 26367
rect 15577 26333 15611 26367
rect 15761 26333 15795 26367
rect 16773 26333 16807 26367
rect 17693 26333 17727 26367
rect 9045 26265 9079 26299
rect 9956 26265 9990 26299
rect 12449 26265 12483 26299
rect 13093 26265 13127 26299
rect 14473 26265 14507 26299
rect 15117 26265 15151 26299
rect 18061 26265 18095 26299
rect 18521 26333 18555 26367
rect 18705 26333 18739 26367
rect 19809 26333 19843 26367
rect 21833 26333 21867 26367
rect 22109 26333 22143 26367
rect 22293 26333 22327 26367
rect 30021 26401 30055 26435
rect 30941 26401 30975 26435
rect 22753 26333 22787 26367
rect 22937 26333 22971 26367
rect 23581 26333 23615 26367
rect 23857 26333 23891 26367
rect 24593 26333 24627 26367
rect 24869 26333 24903 26367
rect 25053 26333 25087 26367
rect 25513 26333 25547 26367
rect 27629 26333 27663 26367
rect 29745 26333 29779 26367
rect 30665 26333 30699 26367
rect 20054 26265 20088 26299
rect 22569 26265 22603 26299
rect 24409 26265 24443 26299
rect 25780 26265 25814 26299
rect 27896 26265 27930 26299
rect 29561 26265 29595 26299
rect 30481 26265 30515 26299
rect 1961 26197 1995 26231
rect 3801 26197 3835 26231
rect 11069 26197 11103 26231
rect 11529 26197 11563 26231
rect 16865 26197 16899 26231
rect 18153 26197 18187 26231
rect 21189 26197 21223 26231
rect 26893 26197 26927 26231
rect 29009 26197 29043 26231
rect 1593 25993 1627 26027
rect 6745 25993 6779 26027
rect 12909 25993 12943 26027
rect 20177 25993 20211 26027
rect 23489 25993 23523 26027
rect 25789 25993 25823 26027
rect 2780 25925 2814 25959
rect 4353 25925 4387 25959
rect 5733 25925 5767 25959
rect 9505 25925 9539 25959
rect 19349 25925 19383 25959
rect 22201 25925 22235 25959
rect 24654 25925 24688 25959
rect 29920 25925 29954 25959
rect 1777 25857 1811 25891
rect 4537 25857 4571 25891
rect 4813 25857 4847 25891
rect 4997 25857 5031 25891
rect 5641 25857 5675 25891
rect 5825 25857 5859 25891
rect 7757 25857 7791 25891
rect 10517 25857 10551 25891
rect 10793 25857 10827 25891
rect 10977 25857 11011 25891
rect 11529 25857 11563 25891
rect 11785 25857 11819 25891
rect 13553 25857 13587 25891
rect 14565 25857 14599 25891
rect 14832 25857 14866 25891
rect 16773 25857 16807 25891
rect 17684 25857 17718 25891
rect 19533 25857 19567 25891
rect 20361 25857 20395 25891
rect 20637 25857 20671 25891
rect 20821 25857 20855 25891
rect 24409 25857 24443 25891
rect 26985 25857 27019 25891
rect 27629 25857 27663 25891
rect 27896 25857 27930 25891
rect 29653 25857 29687 25891
rect 2053 25789 2087 25823
rect 2513 25789 2547 25823
rect 6837 25789 6871 25823
rect 7021 25789 7055 25823
rect 13829 25789 13863 25823
rect 17417 25789 17451 25823
rect 1961 25653 1995 25687
rect 3893 25653 3927 25687
rect 6377 25653 6411 25687
rect 10333 25653 10367 25687
rect 13369 25653 13403 25687
rect 13737 25653 13771 25687
rect 15945 25653 15979 25687
rect 16865 25653 16899 25687
rect 18797 25653 18831 25687
rect 27077 25653 27111 25687
rect 29009 25653 29043 25687
rect 31033 25653 31067 25687
rect 3893 25449 3927 25483
rect 6101 25449 6135 25483
rect 8309 25449 8343 25483
rect 13001 25449 13035 25483
rect 13921 25449 13955 25483
rect 15209 25449 15243 25483
rect 18061 25449 18095 25483
rect 22385 25449 22419 25483
rect 24777 25449 24811 25483
rect 31309 25449 31343 25483
rect 2329 25381 2363 25415
rect 5733 25381 5767 25415
rect 2881 25313 2915 25347
rect 1409 25245 1443 25279
rect 4077 25245 4111 25279
rect 4721 25245 4755 25279
rect 4997 25245 5031 25279
rect 5181 25245 5215 25279
rect 5917 25245 5951 25279
rect 6009 25245 6043 25279
rect 6101 25245 6135 25279
rect 6193 25381 6227 25415
rect 7941 25381 7975 25415
rect 8953 25381 8987 25415
rect 7297 25313 7331 25347
rect 6193 25245 6227 25279
rect 6469 25245 6503 25279
rect 7205 25245 7239 25279
rect 9137 25313 9171 25347
rect 9229 25313 9263 25347
rect 13277 25313 13311 25347
rect 13461 25313 13495 25347
rect 15577 25381 15611 25415
rect 17509 25381 17543 25415
rect 14105 25313 14139 25347
rect 15669 25313 15703 25347
rect 19257 25313 19291 25347
rect 22753 25313 22787 25347
rect 8217 25245 8251 25279
rect 9321 25245 9355 25279
rect 9413 25245 9447 25279
rect 9965 25245 9999 25279
rect 10977 25245 11011 25279
rect 11253 25245 11287 25279
rect 11437 25245 11471 25279
rect 12081 25245 12115 25279
rect 12357 25245 12391 25279
rect 12541 25245 12575 25279
rect 13185 25245 13219 25279
rect 13369 25245 13403 25279
rect 13921 25245 13955 25279
rect 14381 25245 14415 25279
rect 14473 25245 14507 25279
rect 14565 25245 14599 25279
rect 14749 25245 14783 25279
rect 15393 25245 15427 25279
rect 17233 25245 17267 25279
rect 18245 25245 18279 25279
rect 18429 25245 18463 25279
rect 18521 25245 18555 25279
rect 19441 25245 19475 25279
rect 19717 25245 19751 25279
rect 19901 25245 19935 25279
rect 21097 25245 21131 25279
rect 21373 25245 21407 25279
rect 21557 25245 21591 25279
rect 22569 25245 22603 25279
rect 22845 25245 22879 25279
rect 23857 25245 23891 25279
rect 25053 25245 25087 25279
rect 25973 25245 26007 25279
rect 26249 25245 26283 25279
rect 26433 25245 26467 25279
rect 27169 25245 27203 25279
rect 29929 25245 29963 25279
rect 2789 25177 2823 25211
rect 5733 25177 5767 25211
rect 7941 25177 7975 25211
rect 10057 25177 10091 25211
rect 16313 25177 16347 25211
rect 23489 25177 23523 25211
rect 24409 25177 24443 25211
rect 30196 25177 30230 25211
rect 1593 25109 1627 25143
rect 2697 25109 2731 25143
rect 4537 25109 4571 25143
rect 6561 25109 6595 25143
rect 10793 25109 10827 25143
rect 11897 25109 11931 25143
rect 16589 25109 16623 25143
rect 20913 25109 20947 25143
rect 23397 25109 23431 25143
rect 23581 25109 23615 25143
rect 23673 25109 23707 25143
rect 24786 25109 24820 25143
rect 25789 25109 25823 25143
rect 28457 25109 28491 25143
rect 2145 24905 2179 24939
rect 5457 24905 5491 24939
rect 22191 24905 22225 24939
rect 1685 24837 1719 24871
rect 10333 24837 10367 24871
rect 13084 24837 13118 24871
rect 14933 24837 14967 24871
rect 16129 24837 16163 24871
rect 16221 24837 16255 24871
rect 22661 24837 22695 24871
rect 24133 24837 24167 24871
rect 2973 24769 3007 24803
rect 3157 24769 3191 24803
rect 4344 24769 4378 24803
rect 6377 24769 6411 24803
rect 6561 24769 6595 24803
rect 6653 24769 6687 24803
rect 7113 24769 7147 24803
rect 7380 24769 7414 24803
rect 8953 24769 8987 24803
rect 9321 24769 9355 24803
rect 9689 24769 9723 24803
rect 10057 24769 10091 24803
rect 11805 24769 11839 24803
rect 14749 24769 14783 24803
rect 15945 24769 15979 24803
rect 16865 24769 16899 24803
rect 18521 24769 18555 24803
rect 18705 24769 18739 24803
rect 18797 24769 18831 24803
rect 18889 24769 18923 24803
rect 19441 24769 19475 24803
rect 19717 24769 19751 24803
rect 19901 24769 19935 24803
rect 21005 24769 21039 24803
rect 21189 24769 21223 24803
rect 22753 24769 22787 24803
rect 23305 24769 23339 24803
rect 23489 24769 23523 24803
rect 24317 24769 24351 24803
rect 25053 24769 25087 24803
rect 25237 24769 25271 24803
rect 25513 24769 25547 24803
rect 25697 24769 25731 24803
rect 26249 24769 26283 24803
rect 26985 24769 27019 24803
rect 27169 24769 27203 24803
rect 27445 24769 27479 24803
rect 28089 24769 28123 24803
rect 29101 24769 29135 24803
rect 29285 24769 29319 24803
rect 29561 24769 29595 24803
rect 29745 24769 29779 24803
rect 30389 24769 30423 24803
rect 30665 24769 30699 24803
rect 30849 24769 30883 24803
rect 2881 24701 2915 24735
rect 3617 24701 3651 24735
rect 4077 24701 4111 24735
rect 11529 24701 11563 24735
rect 12817 24701 12851 24735
rect 16221 24701 16255 24735
rect 17141 24701 17175 24735
rect 1961 24633 1995 24667
rect 18337 24633 18371 24667
rect 21281 24701 21315 24735
rect 22661 24701 22695 24735
rect 24593 24701 24627 24735
rect 26433 24701 26467 24735
rect 27353 24701 27387 24735
rect 28365 24701 28399 24735
rect 30205 24701 30239 24735
rect 23673 24633 23707 24667
rect 6377 24565 6411 24599
rect 8493 24565 8527 24599
rect 14197 24565 14231 24599
rect 18889 24565 18923 24599
rect 19257 24565 19291 24599
rect 20821 24565 20855 24599
rect 24501 24565 24535 24599
rect 27905 24565 27939 24599
rect 28273 24565 28307 24599
rect 2329 24361 2363 24395
rect 3801 24361 3835 24395
rect 4997 24361 5031 24395
rect 5365 24361 5399 24395
rect 6469 24361 6503 24395
rect 8125 24361 8159 24395
rect 9137 24361 9171 24395
rect 9689 24361 9723 24395
rect 13737 24361 13771 24395
rect 22201 24361 22235 24395
rect 25881 24361 25915 24395
rect 28181 24361 28215 24395
rect 1777 24157 1811 24191
rect 6653 24293 6687 24327
rect 2421 24225 2455 24259
rect 4353 24225 4387 24259
rect 5457 24225 5491 24259
rect 6101 24225 6135 24259
rect 11161 24293 11195 24327
rect 11253 24225 11287 24259
rect 15301 24293 15335 24327
rect 20269 24293 20303 24327
rect 22661 24293 22695 24327
rect 27721 24293 27755 24327
rect 16865 24225 16899 24259
rect 19625 24225 19659 24259
rect 20821 24225 20855 24259
rect 23305 24225 23339 24259
rect 2697 24157 2731 24191
rect 5181 24157 5215 24191
rect 7757 24157 7791 24191
rect 8125 24157 8159 24191
rect 8217 24157 8251 24191
rect 8401 24157 8435 24191
rect 9045 24157 9079 24191
rect 9965 24157 9999 24191
rect 10057 24157 10091 24191
rect 10149 24157 10183 24191
rect 10333 24157 10367 24191
rect 10977 24157 11011 24191
rect 13645 24157 13679 24191
rect 14105 24157 14139 24191
rect 14289 24157 14323 24191
rect 15117 24157 15151 24191
rect 15393 24157 15427 24191
rect 15853 24157 15887 24191
rect 16037 24157 16071 24191
rect 19441 24157 19475 24191
rect 19717 24157 19751 24191
rect 20177 24157 20211 24191
rect 21077 24157 21111 24191
rect 23029 24157 23063 24191
rect 24501 24157 24535 24191
rect 24768 24157 24802 24191
rect 26341 24157 26375 24191
rect 28365 24157 28399 24191
rect 28641 24157 28675 24191
rect 28825 24157 28859 24191
rect 30297 24157 30331 24191
rect 30573 24157 30607 24191
rect 30757 24157 30791 24191
rect 2329 24089 2363 24123
rect 4169 24089 4203 24123
rect 8309 24089 8343 24123
rect 11805 24089 11839 24123
rect 14473 24089 14507 24123
rect 17132 24089 17166 24123
rect 26608 24089 26642 24123
rect 1869 24021 1903 24055
rect 4261 24021 4295 24055
rect 6469 24021 6503 24055
rect 7573 24021 7607 24055
rect 10793 24021 10827 24055
rect 13093 24021 13127 24055
rect 14933 24021 14967 24055
rect 16221 24021 16255 24055
rect 18245 24021 18279 24055
rect 19257 24021 19291 24055
rect 23121 24021 23155 24055
rect 30113 24021 30147 24055
rect 2789 23817 2823 23851
rect 6377 23817 6411 23851
rect 6745 23817 6779 23851
rect 8953 23817 8987 23851
rect 11805 23817 11839 23851
rect 12173 23817 12207 23851
rect 12265 23817 12299 23851
rect 13185 23817 13219 23851
rect 13553 23817 13587 23851
rect 17141 23817 17175 23851
rect 30665 23817 30699 23851
rect 3617 23749 3651 23783
rect 7840 23749 7874 23783
rect 14648 23749 14682 23783
rect 17049 23749 17083 23783
rect 19993 23749 20027 23783
rect 21833 23749 21867 23783
rect 22033 23749 22067 23783
rect 1409 23681 1443 23715
rect 1665 23681 1699 23715
rect 4445 23681 4479 23715
rect 4721 23681 4755 23715
rect 4905 23681 4939 23715
rect 5457 23681 5491 23715
rect 7573 23681 7607 23715
rect 10057 23681 10091 23715
rect 10333 23681 10367 23715
rect 10517 23681 10551 23715
rect 13645 23681 13679 23715
rect 18061 23681 18095 23715
rect 18245 23681 18279 23715
rect 20637 23681 20671 23715
rect 23112 23681 23146 23715
rect 25237 23681 25271 23715
rect 25513 23681 25547 23715
rect 25697 23681 25731 23715
rect 26249 23681 26283 23715
rect 27169 23681 27203 23715
rect 27445 23681 27479 23715
rect 27629 23681 27663 23715
rect 28089 23681 28123 23715
rect 29377 23681 29411 23715
rect 30849 23681 30883 23715
rect 31033 23681 31067 23715
rect 6837 23613 6871 23647
rect 6929 23613 6963 23647
rect 12357 23613 12391 23647
rect 13737 23613 13771 23647
rect 14381 23613 14415 23647
rect 17233 23613 17267 23647
rect 3249 23545 3283 23579
rect 20913 23613 20947 23647
rect 22845 23613 22879 23647
rect 26985 23613 27019 23647
rect 28365 23613 28399 23647
rect 29653 23613 29687 23647
rect 31125 23613 31159 23647
rect 24225 23545 24259 23579
rect 3617 23477 3651 23511
rect 3801 23477 3835 23511
rect 4261 23477 4295 23511
rect 5549 23477 5583 23511
rect 9873 23477 9907 23511
rect 15761 23477 15795 23511
rect 16681 23477 16715 23511
rect 18061 23477 18095 23511
rect 20453 23477 20487 23511
rect 20821 23477 20855 23511
rect 22017 23477 22051 23511
rect 22201 23477 22235 23511
rect 25053 23477 25087 23511
rect 26341 23477 26375 23511
rect 2605 23273 2639 23307
rect 4353 23273 4387 23307
rect 8033 23273 8067 23307
rect 10057 23273 10091 23307
rect 12449 23273 12483 23307
rect 23673 23273 23707 23307
rect 25053 23273 25087 23307
rect 27997 23273 28031 23307
rect 15393 23205 15427 23239
rect 16497 23205 16531 23239
rect 25237 23205 25271 23239
rect 4445 23137 4479 23171
rect 6929 23137 6963 23171
rect 9505 23137 9539 23171
rect 10517 23137 10551 23171
rect 12909 23137 12943 23171
rect 15853 23137 15887 23171
rect 21097 23137 21131 23171
rect 25973 23137 26007 23171
rect 29929 23137 29963 23171
rect 2789 23069 2823 23103
rect 3065 23069 3099 23103
rect 4169 23069 4203 23103
rect 5089 23069 5123 23103
rect 5733 23069 5767 23103
rect 6009 23069 6043 23103
rect 6193 23069 6227 23103
rect 6653 23069 6687 23103
rect 7941 23069 7975 23103
rect 9321 23069 9355 23103
rect 9597 23069 9631 23103
rect 10241 23069 10275 23103
rect 10425 23069 10459 23103
rect 11069 23069 11103 23103
rect 13093 23069 13127 23103
rect 13369 23069 13403 23103
rect 13553 23069 13587 23103
rect 14289 23069 14323 23103
rect 14473 23069 14507 23103
rect 14565 23069 14599 23103
rect 16497 23069 16531 23103
rect 16681 23069 16715 23103
rect 16773 23069 16807 23103
rect 17877 23069 17911 23103
rect 18153 23069 18187 23103
rect 18337 23069 18371 23103
rect 19257 23069 19291 23103
rect 19513 23069 19547 23103
rect 26801 23069 26835 23103
rect 27077 23069 27111 23103
rect 27261 23069 27295 23103
rect 28181 23069 28215 23103
rect 28457 23069 28491 23103
rect 28641 23069 28675 23103
rect 1869 23001 1903 23035
rect 2053 23001 2087 23035
rect 2973 23001 3007 23035
rect 11336 23001 11370 23035
rect 15945 23001 15979 23035
rect 21342 23001 21376 23035
rect 23489 23001 23523 23035
rect 23705 23001 23739 23035
rect 24869 23001 24903 23035
rect 25789 23001 25823 23035
rect 30174 23001 30208 23035
rect 3985 22933 4019 22967
rect 4905 22933 4939 22967
rect 5549 22933 5583 22967
rect 8401 22933 8435 22967
rect 9137 22933 9171 22967
rect 14105 22933 14139 22967
rect 15853 22933 15887 22967
rect 17693 22933 17727 22967
rect 20637 22933 20671 22967
rect 22477 22933 22511 22967
rect 23857 22933 23891 22967
rect 25069 22933 25103 22967
rect 26617 22933 26651 22967
rect 31309 22933 31343 22967
rect 1501 22729 1535 22763
rect 2421 22729 2455 22763
rect 7757 22729 7791 22763
rect 10057 22729 10091 22763
rect 11345 22729 11379 22763
rect 14197 22729 14231 22763
rect 15117 22729 15151 22763
rect 17693 22729 17727 22763
rect 18797 22729 18831 22763
rect 20729 22729 20763 22763
rect 27169 22729 27203 22763
rect 29193 22729 29227 22763
rect 29929 22729 29963 22763
rect 2789 22661 2823 22695
rect 4813 22661 4847 22695
rect 8484 22661 8518 22695
rect 1685 22593 1719 22627
rect 1869 22593 1903 22627
rect 3801 22593 3835 22627
rect 4077 22593 4111 22627
rect 4629 22593 4663 22627
rect 5457 22593 5491 22627
rect 5641 22593 5675 22627
rect 6377 22593 6411 22627
rect 6633 22593 6667 22627
rect 8217 22593 8251 22627
rect 10241 22593 10275 22627
rect 10517 22593 10551 22627
rect 10701 22593 10735 22627
rect 1961 22525 1995 22559
rect 2881 22525 2915 22559
rect 3065 22525 3099 22559
rect 5733 22525 5767 22559
rect 13084 22661 13118 22695
rect 19257 22661 19291 22695
rect 26341 22661 26375 22695
rect 27077 22661 27111 22695
rect 28080 22661 28114 22695
rect 31125 22661 31159 22695
rect 15301 22593 15335 22627
rect 15577 22593 15611 22627
rect 15761 22593 15795 22627
rect 16773 22593 16807 22627
rect 16957 22593 16991 22627
rect 17141 22593 17175 22627
rect 17877 22593 17911 22627
rect 18153 22593 18187 22627
rect 18613 22593 18647 22627
rect 18797 22593 18831 22627
rect 19441 22593 19475 22627
rect 19533 22593 19567 22627
rect 19809 22593 19843 22627
rect 20913 22593 20947 22627
rect 21925 22593 21959 22627
rect 22181 22593 22215 22627
rect 24225 22593 24259 22627
rect 24492 22593 24526 22627
rect 26157 22593 26191 22627
rect 27813 22593 27847 22627
rect 30113 22593 30147 22627
rect 30389 22593 30423 22627
rect 30573 22593 30607 22627
rect 11529 22525 11563 22559
rect 11805 22525 11839 22559
rect 12817 22525 12851 22559
rect 17233 22525 17267 22559
rect 19717 22525 19751 22559
rect 21189 22525 21223 22559
rect 3985 22457 4019 22491
rect 5273 22457 5307 22491
rect 9597 22457 9631 22491
rect 11345 22457 11379 22491
rect 3617 22389 3651 22423
rect 18061 22389 18095 22423
rect 21097 22389 21131 22423
rect 23305 22389 23339 22423
rect 25605 22389 25639 22423
rect 31217 22389 31251 22423
rect 1961 22185 1995 22219
rect 3801 22185 3835 22219
rect 5917 22185 5951 22219
rect 4905 22117 4939 22151
rect 2145 21981 2179 22015
rect 2421 21981 2455 22015
rect 2605 21981 2639 22015
rect 3249 21981 3283 22015
rect 3985 21981 4019 22015
rect 4261 21981 4295 22015
rect 4445 21981 4479 22015
rect 5089 21981 5123 22015
rect 5365 21981 5399 22015
rect 5549 21981 5583 22015
rect 7481 22185 7515 22219
rect 8217 22185 8251 22219
rect 12173 22185 12207 22219
rect 15669 22185 15703 22219
rect 20269 22185 20303 22219
rect 11805 22117 11839 22151
rect 13369 22117 13403 22151
rect 6285 22049 6319 22083
rect 7481 22049 7515 22083
rect 11713 22049 11747 22083
rect 7113 21981 7147 22015
rect 7389 21981 7423 22015
rect 7849 21981 7883 22015
rect 9413 21981 9447 22015
rect 11437 21981 11471 22015
rect 11621 21981 11655 22015
rect 5917 21913 5951 21947
rect 6101 21913 6135 21947
rect 6929 21913 6963 21947
rect 9680 21913 9714 21947
rect 11253 21913 11287 21947
rect 19257 22117 19291 22151
rect 23121 22117 23155 22151
rect 26985 22117 27019 22151
rect 12541 22049 12575 22083
rect 12633 22049 12667 22083
rect 15669 22049 15703 22083
rect 19625 22049 19659 22083
rect 19717 22049 19751 22083
rect 21373 22049 21407 22083
rect 27721 22049 27755 22083
rect 12357 21981 12391 22015
rect 13185 21981 13219 22015
rect 14105 21981 14139 22015
rect 15117 21981 15151 22015
rect 15393 21981 15427 22015
rect 15577 21981 15611 22015
rect 19441 21981 19475 22015
rect 20177 21981 20211 22015
rect 20361 21981 20395 22015
rect 22017 21981 22051 22015
rect 22201 21981 22235 22015
rect 22477 21981 22511 22015
rect 22661 21981 22695 22015
rect 23305 21981 23339 22015
rect 23581 21981 23615 22015
rect 23765 21981 23799 22015
rect 24593 21981 24627 22015
rect 24777 21981 24811 22015
rect 24869 21981 24903 22015
rect 25605 21981 25639 22015
rect 27445 21981 27479 22015
rect 28825 21981 28859 22015
rect 29929 21981 29963 22015
rect 16037 21913 16071 21947
rect 16313 21913 16347 21947
rect 16407 21913 16441 21947
rect 17969 21913 18003 21947
rect 25872 21913 25906 21947
rect 29009 21913 29043 21947
rect 30196 21913 30230 21947
rect 3065 21845 3099 21879
rect 7297 21845 7331 21879
rect 8217 21845 8251 21879
rect 8401 21845 8435 21879
rect 10793 21845 10827 21879
rect 11805 21845 11839 21879
rect 14289 21845 14323 21879
rect 14933 21845 14967 21879
rect 15669 21845 15703 21879
rect 20821 21845 20855 21879
rect 21189 21845 21223 21879
rect 21281 21845 21315 21879
rect 24409 21845 24443 21879
rect 31309 21845 31343 21879
rect 5641 21641 5675 21675
rect 7665 21641 7699 21675
rect 9873 21641 9907 21675
rect 11989 21641 12023 21675
rect 20729 21641 20763 21675
rect 21925 21641 21959 21675
rect 22477 21641 22511 21675
rect 3148 21573 3182 21607
rect 9413 21573 9447 21607
rect 1409 21505 1443 21539
rect 2421 21505 2455 21539
rect 4905 21505 4939 21539
rect 5825 21505 5859 21539
rect 6561 21505 6595 21539
rect 7849 21505 7883 21539
rect 8125 21505 8159 21539
rect 9229 21505 9263 21539
rect 10057 21505 10091 21539
rect 10333 21505 10367 21539
rect 10517 21505 10551 21539
rect 10609 21505 10643 21539
rect 2881 21437 2915 21471
rect 5181 21437 5215 21471
rect 7941 21437 7975 21471
rect 8033 21437 8067 21471
rect 12817 21573 12851 21607
rect 16926 21573 16960 21607
rect 19616 21573 19650 21607
rect 12081 21505 12115 21539
rect 12265 21505 12299 21539
rect 11989 21437 12023 21471
rect 12541 21437 12575 21471
rect 4261 21369 4295 21403
rect 6745 21369 6779 21403
rect 10609 21369 10643 21403
rect 13001 21505 13035 21539
rect 13185 21505 13219 21539
rect 14381 21505 14415 21539
rect 15301 21505 15335 21539
rect 15577 21505 15611 21539
rect 18153 21505 18187 21539
rect 18521 21505 18555 21539
rect 18705 21505 18739 21539
rect 18797 21505 18831 21539
rect 22109 21505 22143 21539
rect 14657 21437 14691 21471
rect 15117 21437 15151 21471
rect 15485 21437 15519 21471
rect 16681 21437 16715 21471
rect 19349 21437 19383 21471
rect 22385 21437 22419 21471
rect 12817 21369 12851 21403
rect 14565 21369 14599 21403
rect 18061 21369 18095 21403
rect 18153 21369 18187 21403
rect 22753 21641 22787 21675
rect 22845 21641 22879 21675
rect 23213 21641 23247 21675
rect 24593 21641 24627 21675
rect 25973 21641 26007 21675
rect 23305 21573 23339 21607
rect 29193 21573 29227 21607
rect 29285 21573 29319 21607
rect 22753 21505 22787 21539
rect 24777 21505 24811 21539
rect 24961 21505 24995 21539
rect 26157 21505 26191 21539
rect 26341 21505 26375 21539
rect 27169 21505 27203 21539
rect 27445 21505 27479 21539
rect 27629 21505 27663 21539
rect 28273 21505 28307 21539
rect 29009 21505 29043 21539
rect 29377 21505 29411 21539
rect 30205 21505 30239 21539
rect 30481 21505 30515 21539
rect 30665 21505 30699 21539
rect 31125 21505 31159 21539
rect 23397 21437 23431 21471
rect 25053 21437 25087 21471
rect 26433 21437 26467 21471
rect 28549 21437 28583 21471
rect 31217 21369 31251 21403
rect 1593 21301 1627 21335
rect 2237 21301 2271 21335
rect 4721 21301 4755 21335
rect 5089 21301 5123 21335
rect 12449 21301 12483 21335
rect 13369 21301 13403 21335
rect 14197 21301 14231 21335
rect 18521 21301 18555 21335
rect 22293 21301 22327 21335
rect 22477 21301 22511 21335
rect 26985 21301 27019 21335
rect 28089 21301 28123 21335
rect 28457 21301 28491 21335
rect 29561 21301 29595 21335
rect 30021 21301 30055 21335
rect 2789 21097 2823 21131
rect 6285 21097 6319 21131
rect 8125 21097 8159 21131
rect 11437 21097 11471 21131
rect 17785 21097 17819 21131
rect 19257 21097 19291 21131
rect 25789 21097 25823 21131
rect 26709 21097 26743 21131
rect 29009 21097 29043 21131
rect 30757 21097 30791 21131
rect 7665 21029 7699 21063
rect 10057 21029 10091 21063
rect 1409 20893 1443 20927
rect 4169 20893 4203 20927
rect 6469 20893 6503 20927
rect 6561 20893 6595 20927
rect 6745 20893 6779 20927
rect 6837 20893 6871 20927
rect 12541 20961 12575 20995
rect 14749 20961 14783 20995
rect 7757 20893 7791 20927
rect 7941 20893 7975 20927
rect 9321 20893 9355 20927
rect 10701 20893 10735 20927
rect 10885 20893 10919 20927
rect 11345 20893 11379 20927
rect 12081 20893 12115 20927
rect 12265 20893 12299 20927
rect 12725 20893 12759 20927
rect 14105 20893 14139 20927
rect 14289 20893 14323 20927
rect 15016 20893 15050 20927
rect 17141 20893 17175 20927
rect 17410 20893 17444 20927
rect 17601 20893 17635 20927
rect 1676 20825 1710 20859
rect 4436 20825 4470 20859
rect 7665 20825 7699 20859
rect 9781 20825 9815 20859
rect 10793 20825 10827 20859
rect 28181 21029 28215 21063
rect 30297 21029 30331 21063
rect 22569 20961 22603 20995
rect 23121 20961 23155 20995
rect 23213 20961 23247 20995
rect 25053 20961 25087 20995
rect 26801 20961 26835 20995
rect 31217 20961 31251 20995
rect 18061 20893 18095 20927
rect 18245 20893 18279 20927
rect 18521 20893 18555 20927
rect 18705 20893 18739 20927
rect 19441 20893 19475 20927
rect 19717 20893 19751 20927
rect 19901 20893 19935 20927
rect 20453 20825 20487 20859
rect 24777 20893 24811 20927
rect 24961 20893 24995 20927
rect 25605 20893 25639 20927
rect 26525 20893 26559 20927
rect 27537 20893 27571 20927
rect 27630 20893 27664 20927
rect 28002 20893 28036 20927
rect 28641 20893 28675 20927
rect 28825 20893 28859 20927
rect 29653 20893 29687 20927
rect 29801 20893 29835 20927
rect 30118 20893 30152 20927
rect 30941 20893 30975 20927
rect 31125 20893 31159 20927
rect 23029 20825 23063 20859
rect 25145 20825 25179 20859
rect 27813 20825 27847 20859
rect 27905 20825 27939 20859
rect 29929 20825 29963 20859
rect 30021 20825 30055 20859
rect 5549 20757 5583 20791
rect 9137 20757 9171 20791
rect 10241 20757 10275 20791
rect 14197 20757 14231 20791
rect 16129 20757 16163 20791
rect 16957 20757 16991 20791
rect 17785 20757 17819 20791
rect 21741 20757 21775 20791
rect 22569 20757 22603 20791
rect 22661 20757 22695 20791
rect 26341 20757 26375 20791
rect 1869 20553 1903 20587
rect 5089 20553 5123 20587
rect 5549 20553 5583 20587
rect 9941 20553 9975 20587
rect 10057 20553 10091 20587
rect 10885 20553 10919 20587
rect 13001 20553 13035 20587
rect 23489 20553 23523 20587
rect 23673 20553 23707 20587
rect 27261 20553 27295 20587
rect 27629 20553 27663 20587
rect 27721 20553 27755 20587
rect 29837 20553 29871 20587
rect 30205 20553 30239 20587
rect 4629 20485 4663 20519
rect 9413 20485 9447 20519
rect 9597 20485 9631 20519
rect 12909 20485 12943 20519
rect 13820 20485 13854 20519
rect 16497 20485 16531 20519
rect 2053 20417 2087 20451
rect 3341 20417 3375 20451
rect 4445 20417 4479 20451
rect 5457 20417 5491 20451
rect 6929 20417 6963 20451
rect 7941 20417 7975 20451
rect 8033 20417 8067 20451
rect 8217 20417 8251 20451
rect 8309 20417 8343 20451
rect 8769 20417 8803 20451
rect 9853 20417 9887 20451
rect 10149 20417 10183 20451
rect 10793 20417 10827 20451
rect 11345 20417 11379 20451
rect 11621 20417 11655 20451
rect 11804 20417 11838 20451
rect 12173 20417 12207 20451
rect 15393 20417 15427 20451
rect 15577 20417 15611 20451
rect 2329 20349 2363 20383
rect 3065 20349 3099 20383
rect 5641 20349 5675 20383
rect 7021 20349 7055 20383
rect 7113 20349 7147 20383
rect 8861 20349 8895 20383
rect 11897 20349 11931 20383
rect 11989 20349 12023 20383
rect 13553 20349 13587 20383
rect 17877 20485 17911 20519
rect 18225 20485 18259 20519
rect 19441 20485 19475 20519
rect 16865 20417 16899 20451
rect 16957 20417 16991 20451
rect 17233 20417 17267 20451
rect 6561 20281 6595 20315
rect 11529 20281 11563 20315
rect 14933 20281 14967 20315
rect 16497 20281 16531 20315
rect 17141 20281 17175 20315
rect 17969 20417 18003 20451
rect 21097 20417 21131 20451
rect 21281 20417 21315 20451
rect 22017 20417 22051 20451
rect 22201 20417 22235 20451
rect 23121 20417 23155 20451
rect 24133 20417 24167 20451
rect 25329 20417 25363 20451
rect 26157 20417 26191 20451
rect 29101 20417 29135 20451
rect 29193 20417 29227 20451
rect 30021 20417 30055 20451
rect 30297 20417 30331 20451
rect 30941 20417 30975 20451
rect 19809 20349 19843 20383
rect 20085 20349 20119 20383
rect 22293 20349 22327 20383
rect 24317 20349 24351 20383
rect 25145 20349 25179 20383
rect 26433 20349 26467 20383
rect 27813 20349 27847 20383
rect 29009 20349 29043 20383
rect 29285 20349 29319 20383
rect 31217 20349 31251 20383
rect 21189 20281 21223 20315
rect 2237 20213 2271 20247
rect 7757 20213 7791 20247
rect 12265 20213 12299 20247
rect 15761 20213 15795 20247
rect 16681 20213 16715 20247
rect 17877 20213 17911 20247
rect 19349 20213 19383 20247
rect 19441 20213 19475 20247
rect 21833 20213 21867 20247
rect 23489 20213 23523 20247
rect 25513 20213 25547 20247
rect 25973 20213 26007 20247
rect 26341 20213 26375 20247
rect 28825 20213 28859 20247
rect 30757 20213 30791 20247
rect 31125 20213 31159 20247
rect 2145 20009 2179 20043
rect 5181 20009 5215 20043
rect 7021 20009 7055 20043
rect 13645 20009 13679 20043
rect 17417 20009 17451 20043
rect 17785 20009 17819 20043
rect 19625 20009 19659 20043
rect 23857 20009 23891 20043
rect 24225 20009 24259 20043
rect 24777 20009 24811 20043
rect 25053 20009 25087 20043
rect 27261 20009 27295 20043
rect 28365 20009 28399 20043
rect 1593 19941 1627 19975
rect 7665 19941 7699 19975
rect 9413 19941 9447 19975
rect 5641 19873 5675 19907
rect 8309 19873 8343 19907
rect 11713 19873 11747 19907
rect 15117 19941 15151 19975
rect 14105 19873 14139 19907
rect 15761 19873 15795 19907
rect 16865 19873 16899 19907
rect 17233 19873 17267 19907
rect 1409 19805 1443 19839
rect 2329 19805 2363 19839
rect 2605 19805 2639 19839
rect 2789 19805 2823 19839
rect 3801 19805 3835 19839
rect 9413 19805 9447 19839
rect 9965 19805 9999 19839
rect 10057 19805 10091 19839
rect 10517 19805 10551 19839
rect 11253 19805 11287 19839
rect 11897 19805 11931 19839
rect 12081 19805 12115 19839
rect 12909 19805 12943 19839
rect 13093 19805 13127 19839
rect 13185 19805 13219 19839
rect 13311 19805 13345 19839
rect 13553 19805 13587 19839
rect 13645 19805 13679 19839
rect 14289 19805 14323 19839
rect 14565 19805 14599 19839
rect 15485 19805 15519 19839
rect 4046 19737 4080 19771
rect 5908 19737 5942 19771
rect 21557 19941 21591 19975
rect 22477 19873 22511 19907
rect 27721 19941 27755 19975
rect 29929 19873 29963 19907
rect 17969 19805 18003 19839
rect 22733 19805 22767 19839
rect 24225 19805 24259 19839
rect 24409 19805 24443 19839
rect 24593 19805 24627 19839
rect 25053 19805 25087 19839
rect 25237 19805 25271 19839
rect 25421 19805 25455 19839
rect 25881 19805 25915 19839
rect 26148 19805 26182 19839
rect 27721 19805 27755 19839
rect 27905 19805 27939 19839
rect 28549 19805 28583 19839
rect 28641 19805 28675 19839
rect 28825 19805 28859 19839
rect 28917 19805 28951 19839
rect 30196 19805 30230 19839
rect 18153 19737 18187 19771
rect 19441 19737 19475 19771
rect 20269 19737 20303 19771
rect 949 19669 983 19703
rect 8033 19669 8067 19703
rect 8125 19669 8159 19703
rect 14473 19669 14507 19703
rect 15577 19669 15611 19703
rect 17049 19669 17083 19703
rect 17693 19669 17727 19703
rect 19641 19669 19675 19703
rect 19809 19669 19843 19703
rect 25329 19669 25363 19703
rect 31309 19669 31343 19703
rect 4353 19465 4387 19499
rect 7021 19465 7055 19499
rect 7205 19465 7239 19499
rect 12909 19465 12943 19499
rect 13369 19465 13403 19499
rect 14289 19465 14323 19499
rect 15393 19465 15427 19499
rect 15761 19465 15795 19499
rect 16497 19465 16531 19499
rect 16865 19465 16899 19499
rect 17141 19465 17175 19499
rect 10885 19397 10919 19431
rect 11774 19397 11808 19431
rect 1409 19329 1443 19363
rect 1676 19329 1710 19363
rect 3433 19329 3467 19363
rect 3709 19329 3743 19363
rect 3893 19329 3927 19363
rect 4537 19329 4571 19363
rect 4997 19329 5031 19363
rect 5273 19329 5307 19363
rect 7665 19329 7699 19363
rect 7932 19329 7966 19363
rect 9505 19329 9539 19363
rect 9689 19329 9723 19363
rect 10517 19329 10551 19363
rect 11529 19329 11563 19363
rect 13553 19329 13587 19363
rect 13737 19329 13771 19363
rect 14473 19329 14507 19363
rect 14749 19329 14783 19363
rect 14933 19329 14967 19363
rect 15853 19329 15887 19363
rect 6653 19261 6687 19295
rect 9597 19261 9631 19295
rect 10701 19261 10735 19295
rect 13829 19261 13863 19295
rect 15945 19261 15979 19295
rect 10793 19193 10827 19227
rect 11345 19193 11379 19227
rect 2789 19125 2823 19159
rect 3249 19125 3283 19159
rect 7021 19125 7055 19159
rect 9045 19125 9079 19159
rect 10977 19125 11011 19159
rect 16681 19329 16715 19363
rect 16865 19329 16899 19363
rect 17049 19329 17083 19363
rect 16497 19125 16531 19159
rect 18245 19465 18279 19499
rect 17509 19329 17543 19363
rect 17785 19329 17819 19363
rect 17969 19329 18003 19363
rect 18061 19329 18095 19363
rect 17141 19193 17175 19227
rect 17049 19125 17083 19159
rect 17325 19125 17359 19159
rect 18153 19125 18187 19159
rect 19165 19465 19199 19499
rect 21833 19465 21867 19499
rect 23213 19465 23247 19499
rect 25605 19465 25639 19499
rect 27997 19465 28031 19499
rect 28549 19465 28583 19499
rect 30113 19465 30147 19499
rect 18613 19329 18647 19363
rect 18889 19329 18923 19363
rect 19073 19329 19107 19363
rect 19165 19329 19199 19363
rect 19809 19329 19843 19363
rect 21005 19329 21039 19363
rect 21189 19329 21223 19363
rect 22017 19329 22051 19363
rect 22293 19329 22327 19363
rect 22477 19329 22511 19363
rect 24225 19329 24259 19363
rect 24481 19329 24515 19363
rect 26065 19329 26099 19363
rect 26249 19329 26283 19363
rect 27445 19329 27479 19363
rect 19533 19261 19567 19295
rect 20821 19261 20855 19295
rect 23397 19261 23431 19295
rect 23489 19261 23523 19295
rect 23581 19261 23615 19295
rect 23673 19261 23707 19295
rect 27721 19261 27755 19295
rect 18429 19193 18463 19227
rect 28641 19397 28675 19431
rect 30573 19397 30607 19431
rect 29561 19329 29595 19363
rect 29745 19329 29779 19363
rect 29833 19329 29867 19363
rect 29929 19329 29963 19363
rect 30757 19329 30791 19363
rect 30849 19329 30883 19363
rect 31033 19329 31067 19363
rect 31125 19329 31159 19363
rect 28733 19261 28767 19295
rect 18245 19125 18279 19159
rect 26157 19125 26191 19159
rect 27261 19125 27295 19159
rect 27629 19125 27663 19159
rect 27997 19125 28031 19159
rect 28181 19125 28215 19159
rect 6653 18921 6687 18955
rect 9689 18921 9723 18955
rect 9781 18921 9815 18955
rect 13829 18921 13863 18955
rect 14289 18921 14323 18955
rect 17693 18921 17727 18955
rect 21189 18921 21223 18955
rect 22293 18921 22327 18955
rect 23857 18921 23891 18955
rect 1409 18853 1443 18887
rect 8125 18853 8159 18887
rect 8953 18853 8987 18887
rect 6285 18785 6319 18819
rect 1593 18717 1627 18751
rect 2237 18717 2271 18751
rect 2513 18717 2547 18751
rect 2697 18717 2731 18751
rect 4537 18717 4571 18751
rect 4813 18717 4847 18751
rect 7389 18717 7423 18751
rect 7481 18717 7515 18751
rect 8309 18717 8343 18751
rect 8401 18717 8435 18751
rect 9229 18717 9263 18751
rect 3893 18649 3927 18683
rect 4077 18649 4111 18683
rect 8125 18649 8159 18683
rect 8953 18649 8987 18683
rect 12725 18853 12759 18887
rect 17325 18853 17359 18887
rect 11989 18785 12023 18819
rect 13737 18785 13771 18819
rect 13829 18785 13863 18819
rect 28917 18853 28951 18887
rect 29561 18853 29595 18887
rect 30205 18853 30239 18887
rect 17693 18785 17727 18819
rect 18245 18785 18279 18819
rect 19809 18785 19843 18819
rect 24501 18785 24535 18819
rect 27261 18785 27295 18819
rect 28181 18785 28215 18819
rect 9965 18717 9999 18751
rect 10238 18727 10272 18761
rect 10977 18717 11011 18751
rect 11621 18717 11655 18751
rect 11805 18717 11839 18751
rect 13185 18717 13219 18751
rect 10149 18649 10183 18683
rect 11161 18649 11195 18683
rect 12541 18649 12575 18683
rect 14105 18717 14139 18751
rect 15301 18717 15335 18751
rect 15577 18717 15611 18751
rect 16957 18717 16991 18751
rect 17141 18717 17175 18751
rect 17417 18717 17451 18751
rect 18429 18717 18463 18751
rect 18705 18717 18739 18751
rect 21925 18717 21959 18751
rect 23213 18717 23247 18751
rect 23489 18717 23523 18751
rect 24777 18717 24811 18751
rect 25789 18717 25823 18751
rect 26056 18717 26090 18751
rect 28089 18717 28123 18751
rect 28825 18717 28859 18751
rect 29745 18717 29779 18751
rect 30389 18717 30423 18751
rect 30665 18717 30699 18751
rect 30849 18717 30883 18751
rect 20054 18649 20088 18683
rect 23698 18649 23732 18683
rect 27261 18649 27295 18683
rect 27997 18649 28031 18683
rect 2053 18581 2087 18615
rect 6653 18581 6687 18615
rect 6837 18581 6871 18615
rect 9137 18581 9171 18615
rect 9689 18581 9723 18615
rect 13369 18581 13403 18615
rect 13737 18581 13771 18615
rect 18613 18581 18647 18615
rect 22293 18581 22327 18615
rect 22477 18581 22511 18615
rect 23581 18581 23615 18615
rect 27169 18581 27203 18615
rect 27629 18581 27663 18615
rect 1777 18377 1811 18411
rect 3709 18377 3743 18411
rect 6377 18377 6411 18411
rect 6929 18377 6963 18411
rect 7481 18377 7515 18411
rect 18061 18377 18095 18411
rect 19533 18377 19567 18411
rect 22017 18377 22051 18411
rect 24317 18377 24351 18411
rect 1961 18241 1995 18275
rect 2973 18241 3007 18275
rect 3157 18241 3191 18275
rect 4160 18309 4194 18343
rect 8677 18309 8711 18343
rect 8861 18309 8895 18343
rect 18521 18309 18555 18343
rect 21833 18309 21867 18343
rect 6621 18241 6655 18275
rect 6929 18241 6963 18275
rect 7665 18241 7699 18275
rect 7757 18241 7791 18275
rect 7941 18241 7975 18275
rect 8033 18241 8067 18275
rect 9505 18241 9539 18275
rect 10241 18241 10275 18275
rect 10425 18241 10459 18275
rect 10701 18241 10735 18275
rect 10885 18241 10919 18275
rect 11805 18241 11839 18275
rect 12081 18241 12115 18275
rect 13001 18241 13035 18275
rect 13737 18241 13771 18275
rect 14004 18241 14038 18275
rect 15577 18241 15611 18275
rect 15761 18241 15795 18275
rect 16037 18241 16071 18275
rect 16681 18241 16715 18275
rect 16937 18241 16971 18275
rect 18706 18241 18740 18275
rect 18797 18241 18831 18275
rect 19073 18241 19107 18275
rect 19717 18241 19751 18275
rect 20453 18241 20487 18275
rect 20637 18241 20671 18275
rect 20913 18241 20947 18275
rect 21097 18241 21131 18275
rect 22109 18241 22143 18275
rect 22836 18241 22870 18275
rect 2237 18173 2271 18207
rect 3249 18173 3283 18207
rect 3709 18173 3743 18207
rect 3893 18173 3927 18207
rect 6745 18173 6779 18207
rect 6837 18173 6871 18207
rect 9781 18173 9815 18207
rect 15945 18173 15979 18207
rect 19993 18173 20027 18207
rect 22569 18173 22603 18207
rect 2145 18105 2179 18139
rect 11621 18105 11655 18139
rect 13185 18105 13219 18139
rect 23949 18105 23983 18139
rect 26801 18377 26835 18411
rect 26985 18377 27019 18411
rect 28289 18377 28323 18411
rect 28917 18377 28951 18411
rect 29653 18377 29687 18411
rect 30021 18377 30055 18411
rect 24409 18309 24443 18343
rect 24625 18309 24659 18343
rect 25237 18241 25271 18275
rect 25513 18241 25547 18275
rect 24777 18105 24811 18139
rect 28089 18309 28123 18343
rect 27169 18241 27203 18275
rect 27445 18241 27479 18275
rect 27629 18241 27663 18275
rect 29101 18241 29135 18275
rect 29377 18241 29411 18275
rect 29515 18241 29549 18275
rect 30205 18241 30239 18275
rect 30849 18241 30883 18275
rect 31125 18241 31159 18275
rect 31309 18241 31343 18275
rect 29653 18173 29687 18207
rect 28457 18105 28491 18139
rect 2789 18037 2823 18071
rect 5273 18037 5307 18071
rect 9321 18037 9355 18071
rect 9689 18037 9723 18071
rect 11989 18037 12023 18071
rect 15117 18037 15151 18071
rect 18981 18037 19015 18071
rect 19901 18037 19935 18071
rect 21833 18037 21867 18071
rect 24317 18037 24351 18071
rect 24593 18037 24627 18071
rect 26801 18037 26835 18071
rect 28273 18037 28307 18071
rect 30665 18037 30699 18071
rect 2789 17833 2823 17867
rect 3157 17833 3191 17867
rect 5181 17833 5215 17867
rect 7573 17833 7607 17867
rect 14289 17833 14323 17867
rect 18153 17833 18187 17867
rect 22109 17833 22143 17867
rect 23213 17833 23247 17867
rect 23765 17833 23799 17867
rect 27813 17833 27847 17867
rect 31309 17833 31343 17867
rect 2053 17765 2087 17799
rect 11437 17765 11471 17799
rect 1685 17697 1719 17731
rect 3249 17697 3283 17731
rect 5733 17697 5767 17731
rect 8125 17697 8159 17731
rect 11345 17697 11379 17731
rect 2973 17629 3007 17663
rect 3985 17629 4019 17663
rect 4261 17629 4295 17663
rect 4445 17629 4479 17663
rect 8033 17629 8067 17663
rect 3801 17561 3835 17595
rect 5089 17561 5123 17595
rect 6000 17561 6034 17595
rect 9321 17561 9355 17595
rect 11345 17561 11379 17595
rect 12265 17765 12299 17799
rect 11713 17629 11747 17663
rect 11989 17629 12023 17663
rect 12173 17629 12207 17663
rect 12357 17765 12391 17799
rect 16497 17697 16531 17731
rect 17785 17697 17819 17731
rect 20269 17697 20303 17731
rect 22845 17697 22879 17731
rect 23029 17697 23063 17731
rect 27997 17697 28031 17731
rect 29929 17697 29963 17731
rect 12357 17629 12391 17663
rect 12541 17629 12575 17663
rect 12817 17629 12851 17663
rect 13093 17629 13127 17663
rect 13277 17629 13311 17663
rect 15025 17629 15059 17663
rect 15301 17629 15335 17663
rect 15485 17629 15519 17663
rect 16773 17629 16807 17663
rect 17969 17629 18003 17663
rect 18245 17629 18279 17663
rect 19993 17629 20027 17663
rect 20177 17629 20211 17663
rect 20729 17629 20763 17663
rect 22753 17629 22787 17663
rect 22937 17629 22971 17663
rect 23213 17629 23247 17663
rect 23581 17629 23615 17663
rect 24593 17629 24627 17663
rect 24869 17629 24903 17663
rect 25053 17629 25087 17663
rect 27721 17629 27755 17663
rect 12265 17561 12299 17595
rect 14197 17561 14231 17595
rect 14841 17561 14875 17595
rect 19809 17561 19843 17595
rect 20974 17561 21008 17595
rect 25513 17561 25547 17595
rect 28825 17561 28859 17595
rect 29009 17561 29043 17595
rect 30196 17561 30230 17595
rect 2145 17493 2179 17527
rect 7113 17493 7147 17527
rect 7941 17493 7975 17527
rect 10609 17493 10643 17527
rect 11437 17493 11471 17527
rect 11529 17493 11563 17527
rect 12541 17493 12575 17527
rect 12633 17493 12667 17527
rect 17601 17493 17635 17527
rect 17693 17493 17727 17527
rect 22569 17493 22603 17527
rect 24409 17493 24443 17527
rect 26801 17493 26835 17527
rect 28273 17493 28307 17527
rect 4077 17289 4111 17323
rect 5457 17289 5491 17323
rect 7113 17289 7147 17323
rect 7297 17289 7331 17323
rect 8125 17289 8159 17323
rect 10885 17289 10919 17323
rect 11529 17289 11563 17323
rect 17233 17289 17267 17323
rect 18981 17289 19015 17323
rect 20177 17289 20211 17323
rect 22385 17289 22419 17323
rect 23121 17289 23155 17323
rect 24041 17289 24075 17323
rect 26985 17289 27019 17323
rect 2789 17221 2823 17255
rect 4997 17221 5031 17255
rect 1501 17153 1535 17187
rect 1685 17153 1719 17187
rect 2145 17153 2179 17187
rect 2329 17153 2363 17187
rect 8217 17153 8251 17187
rect 8953 17153 8987 17187
rect 9220 17153 9254 17187
rect 10793 17153 10827 17187
rect 11713 17153 11747 17187
rect 12541 17153 12575 17187
rect 12808 17153 12842 17187
rect 14381 17153 14415 17187
rect 14565 17153 14599 17187
rect 14841 17153 14875 17187
rect 15669 17153 15703 17187
rect 15945 17153 15979 17187
rect 16129 17153 16163 17187
rect 16865 17153 16899 17187
rect 17049 17153 17083 17187
rect 8401 17085 8435 17119
rect 11989 17085 12023 17119
rect 15485 17085 15519 17119
rect 17141 17085 17175 17119
rect 17233 17085 17267 17119
rect 17509 17221 17543 17255
rect 17868 17221 17902 17255
rect 19717 17221 19751 17255
rect 27874 17221 27908 17255
rect 17608 17153 17642 17187
rect 19533 17153 19567 17187
rect 20361 17153 20395 17187
rect 20637 17153 20671 17187
rect 20821 17153 20855 17187
rect 22017 17153 22051 17187
rect 22201 17153 22235 17187
rect 23305 17153 23339 17187
rect 24225 17153 24259 17187
rect 24501 17153 24535 17187
rect 25217 17153 25251 17187
rect 27169 17153 27203 17187
rect 27629 17153 27663 17187
rect 29653 17153 29687 17187
rect 30297 17153 30331 17187
rect 30573 17153 30607 17187
rect 30757 17153 30791 17187
rect 23581 17085 23615 17119
rect 24961 17085 24995 17119
rect 5273 17017 5307 17051
rect 6745 17017 6779 17051
rect 7757 17017 7791 17051
rect 14749 17017 14783 17051
rect 16681 17017 16715 17051
rect 17509 17017 17543 17051
rect 1501 16949 1535 16983
rect 2145 16949 2179 16983
rect 7113 16949 7147 16983
rect 10333 16949 10367 16983
rect 11897 16949 11931 16983
rect 13921 16949 13955 16983
rect 23489 16949 23523 16983
rect 24409 16949 24443 16983
rect 26341 16949 26375 16983
rect 29009 16949 29043 16983
rect 29469 16949 29503 16983
rect 30113 16949 30147 16983
rect 7941 16745 7975 16779
rect 8309 16745 8343 16779
rect 12633 16745 12667 16779
rect 22109 16745 22143 16779
rect 24409 16745 24443 16779
rect 25973 16745 26007 16779
rect 26709 16745 26743 16779
rect 6101 16677 6135 16711
rect 17509 16677 17543 16711
rect 3801 16609 3835 16643
rect 6929 16609 6963 16643
rect 8401 16609 8435 16643
rect 9413 16609 9447 16643
rect 11253 16609 11287 16643
rect 14105 16609 14139 16643
rect 16773 16609 16807 16643
rect 19349 16609 19383 16643
rect 19809 16609 19843 16643
rect 20821 16609 20855 16643
rect 30849 16677 30883 16711
rect 2145 16541 2179 16575
rect 2237 16541 2271 16575
rect 3985 16541 4019 16575
rect 5089 16541 5123 16575
rect 7113 16541 7147 16575
rect 7205 16541 7239 16575
rect 7389 16541 7423 16575
rect 7481 16541 7515 16575
rect 8125 16541 8159 16575
rect 11520 16541 11554 16575
rect 14372 16541 14406 16575
rect 16129 16541 16163 16575
rect 16589 16541 16623 16575
rect 16681 16541 16715 16575
rect 17785 16541 17819 16575
rect 18061 16541 18095 16575
rect 19533 16541 19567 16575
rect 19717 16541 19751 16575
rect 21005 16541 21039 16575
rect 21281 16541 21315 16575
rect 21557 16541 21591 16575
rect 22569 16541 22603 16575
rect 22845 16541 22879 16575
rect 23029 16541 23063 16575
rect 23581 16541 23615 16575
rect 2605 16473 2639 16507
rect 2973 16473 3007 16507
rect 4169 16473 4203 16507
rect 5181 16473 5215 16507
rect 5549 16473 5583 16507
rect 5917 16473 5951 16507
rect 9658 16473 9692 16507
rect 13277 16473 13311 16507
rect 24869 16541 24903 16575
rect 25145 16541 25179 16575
rect 25329 16541 25363 16575
rect 26617 16541 26651 16575
rect 26893 16541 26927 16575
rect 27721 16541 27755 16575
rect 28273 16541 28307 16575
rect 29561 16541 29595 16575
rect 25881 16473 25915 16507
rect 28457 16473 28491 16507
rect 1869 16405 1903 16439
rect 3157 16405 3191 16439
rect 4813 16405 4847 16439
rect 10793 16405 10827 16439
rect 13369 16405 13403 16439
rect 15485 16405 15519 16439
rect 16129 16405 16163 16439
rect 16221 16405 16255 16439
rect 17969 16405 18003 16439
rect 21189 16405 21223 16439
rect 21649 16405 21683 16439
rect 22385 16405 22419 16439
rect 23765 16405 23799 16439
rect 23949 16405 23983 16439
rect 24685 16405 24719 16439
rect 27169 16405 27203 16439
rect 5089 16201 5123 16235
rect 5917 16201 5951 16235
rect 7297 16201 7331 16235
rect 7481 16201 7515 16235
rect 8309 16201 8343 16235
rect 9229 16201 9263 16235
rect 11805 16201 11839 16235
rect 18429 16201 18463 16235
rect 20269 16201 20303 16235
rect 23673 16201 23707 16235
rect 24961 16201 24995 16235
rect 2136 16133 2170 16167
rect 16129 16133 16163 16167
rect 4077 16065 4111 16099
rect 5457 16065 5491 16099
rect 5549 16065 5583 16099
rect 5917 16065 5951 16099
rect 8125 16065 8159 16099
rect 9413 16065 9447 16099
rect 10149 16065 10183 16099
rect 10333 16065 10367 16099
rect 10609 16065 10643 16099
rect 10793 16065 10827 16099
rect 11989 16065 12023 16099
rect 12265 16065 12299 16099
rect 12449 16065 12483 16099
rect 13553 16065 13587 16099
rect 15126 16065 15160 16099
rect 15393 16065 15427 16099
rect 15577 16065 15611 16099
rect 1869 15997 1903 16031
rect 3801 15997 3835 16031
rect 5641 15997 5675 16031
rect 6929 15997 6963 16031
rect 7941 15997 7975 16031
rect 9689 15997 9723 16031
rect 13277 15997 13311 16031
rect 16129 15997 16163 16031
rect 16681 16133 16715 16167
rect 17294 16133 17328 16167
rect 19156 16133 19190 16167
rect 21097 16133 21131 16167
rect 18889 16065 18923 16099
rect 20729 16065 20763 16099
rect 21833 16065 21867 16099
rect 22100 16065 22134 16099
rect 23857 16065 23891 16099
rect 24501 16065 24535 16099
rect 17049 15997 17083 16031
rect 24317 15997 24351 16031
rect 24869 15997 24903 16031
rect 24961 15997 24995 16031
rect 25789 16201 25823 16235
rect 31217 16201 31251 16235
rect 26341 16133 26375 16167
rect 29377 16133 29411 16167
rect 26065 16065 26099 16099
rect 27077 16065 27111 16099
rect 28273 16065 28307 16099
rect 29193 16065 29227 16099
rect 29837 16065 29871 16099
rect 30104 16065 30138 16099
rect 25789 15997 25823 16031
rect 25881 15997 25915 16031
rect 26433 15997 26467 16031
rect 27353 15997 27387 16031
rect 28089 15997 28123 16031
rect 28641 15997 28675 16031
rect 3249 15929 3283 15963
rect 9597 15929 9631 15963
rect 16681 15929 16715 15963
rect 24777 15929 24811 15963
rect 27629 15929 27663 15963
rect 28549 15929 28583 15963
rect 949 15861 983 15895
rect 7297 15861 7331 15895
rect 14933 15861 14967 15895
rect 21097 15861 21131 15895
rect 21281 15861 21315 15895
rect 23213 15861 23247 15895
rect 27445 15861 27479 15895
rect 1409 15657 1443 15691
rect 3801 15657 3835 15691
rect 4997 15657 5031 15691
rect 15761 15657 15795 15691
rect 18245 15657 18279 15691
rect 19533 15657 19567 15691
rect 24501 15657 24535 15691
rect 24961 15657 24995 15691
rect 29009 15657 29043 15691
rect 30665 15657 30699 15691
rect 2881 15589 2915 15623
rect 6285 15589 6319 15623
rect 7113 15589 7147 15623
rect 8309 15589 8343 15623
rect 13645 15589 13679 15623
rect 27997 15589 28031 15623
rect 31033 15589 31067 15623
rect 2053 15521 2087 15555
rect 4353 15521 4387 15555
rect 5457 15521 5491 15555
rect 5549 15521 5583 15555
rect 6837 15521 6871 15555
rect 1777 15453 1811 15487
rect 2605 15385 2639 15419
rect 4169 15385 4203 15419
rect 4261 15385 4295 15419
rect 5365 15385 5399 15419
rect 6653 15385 6687 15419
rect 7297 15521 7331 15555
rect 8953 15521 8987 15555
rect 17233 15521 17267 15555
rect 17877 15521 17911 15555
rect 23397 15521 23431 15555
rect 27537 15521 27571 15555
rect 8217 15453 8251 15487
rect 11161 15453 11195 15487
rect 11345 15453 11379 15487
rect 11437 15453 11471 15487
rect 11897 15453 11931 15487
rect 12173 15453 12207 15487
rect 13369 15453 13403 15487
rect 13645 15453 13679 15487
rect 13737 15453 13771 15487
rect 14473 15453 14507 15487
rect 17141 15453 17175 15487
rect 18061 15453 18095 15487
rect 19717 15453 19751 15487
rect 19993 15453 20027 15487
rect 20177 15453 20211 15487
rect 20821 15453 20855 15487
rect 23581 15453 23615 15487
rect 23765 15453 23799 15487
rect 23857 15453 23891 15487
rect 24041 15453 24075 15487
rect 24409 15453 24443 15487
rect 24777 15453 24811 15487
rect 25605 15453 25639 15487
rect 27721 15453 27755 15487
rect 28089 15453 28123 15487
rect 28641 15453 28675 15487
rect 28733 15453 28767 15487
rect 28825 15453 28859 15487
rect 29745 15453 29779 15487
rect 30021 15453 30055 15487
rect 30205 15453 30239 15487
rect 30849 15453 30883 15487
rect 31125 15453 31159 15487
rect 7297 15385 7331 15419
rect 7573 15385 7607 15419
rect 9220 15385 9254 15419
rect 13553 15385 13587 15419
rect 17049 15385 17083 15419
rect 25872 15385 25906 15419
rect 29561 15385 29595 15419
rect 1869 15317 1903 15351
rect 3065 15317 3099 15351
rect 6745 15317 6779 15351
rect 7113 15317 7147 15351
rect 7665 15317 7699 15351
rect 10333 15317 10367 15351
rect 10977 15317 11011 15351
rect 13645 15317 13679 15351
rect 14105 15317 14139 15351
rect 14289 15317 14323 15351
rect 16681 15317 16715 15351
rect 22109 15317 22143 15351
rect 24041 15317 24075 15351
rect 26985 15317 27019 15351
rect 2605 15113 2639 15147
rect 4353 15113 4387 15147
rect 5825 15113 5859 15147
rect 15393 15113 15427 15147
rect 16037 15113 16071 15147
rect 16497 15113 16531 15147
rect 17049 15113 17083 15147
rect 17877 15113 17911 15147
rect 22109 15113 22143 15147
rect 27629 15113 27663 15147
rect 29745 15113 29779 15147
rect 30665 15113 30699 15147
rect 1501 15045 1535 15079
rect 2513 14977 2547 15011
rect 3525 14977 3559 15011
rect 3801 14977 3835 15011
rect 3985 14977 4019 15011
rect 2789 14909 2823 14943
rect 6837 15045 6871 15079
rect 12164 15045 12198 15079
rect 15485 15045 15519 15079
rect 4712 14977 4746 15011
rect 7849 14977 7883 15011
rect 8105 14977 8139 15011
rect 10057 14977 10091 15011
rect 10333 14977 10367 15011
rect 10517 14977 10551 15011
rect 14013 14977 14047 15011
rect 14280 14977 14314 15011
rect 4445 14909 4479 14943
rect 11897 14909 11931 14943
rect 1685 14841 1719 14875
rect 3341 14841 3375 14875
rect 4353 14841 4387 14875
rect 19809 15045 19843 15079
rect 19993 15045 20027 15079
rect 15945 14977 15979 15011
rect 16497 14977 16531 15011
rect 16773 14977 16807 15011
rect 16865 14977 16899 15011
rect 17877 14977 17911 15011
rect 17969 14977 18003 15011
rect 18889 14977 18923 15011
rect 20913 14977 20947 15011
rect 21005 14977 21039 15011
rect 21097 14977 21131 15011
rect 22293 14977 22327 15011
rect 22477 14977 22511 15011
rect 23121 14977 23155 15011
rect 23388 14977 23422 15011
rect 24869 14977 24903 15011
rect 25053 14977 25087 15011
rect 25237 14977 25271 15011
rect 25973 14977 26007 15011
rect 26249 14977 26283 15011
rect 26433 14977 26467 15011
rect 27077 14977 27111 15011
rect 28365 14977 28399 15011
rect 28632 14977 28666 15011
rect 30849 14977 30883 15011
rect 31125 14977 31159 15011
rect 20177 14909 20211 14943
rect 20821 14909 20855 14943
rect 22569 14909 22603 14943
rect 27353 14909 27387 14943
rect 18337 14841 18371 14875
rect 20637 14841 20671 14875
rect 24869 14841 24903 14875
rect 31033 14841 31067 14875
rect 2145 14773 2179 14807
rect 6929 14773 6963 14807
rect 9229 14773 9263 14807
rect 9873 14773 9907 14807
rect 13277 14773 13311 14807
rect 15485 14773 15519 14807
rect 18429 14773 18463 14807
rect 19073 14773 19107 14807
rect 24501 14773 24535 14807
rect 25789 14773 25823 14807
rect 27169 14773 27203 14807
rect 8309 14569 8343 14603
rect 14105 14569 14139 14603
rect 15301 14569 15335 14603
rect 23397 14569 23431 14603
rect 25973 14569 26007 14603
rect 27445 14569 27479 14603
rect 27721 14569 27755 14603
rect 28549 14569 28583 14603
rect 9689 14501 9723 14535
rect 13553 14501 13587 14535
rect 4445 14433 4479 14467
rect 6285 14433 6319 14467
rect 10241 14433 10275 14467
rect 1409 14365 1443 14399
rect 4261 14365 4295 14399
rect 4997 14365 5031 14399
rect 5181 14365 5215 14399
rect 6009 14365 6043 14399
rect 7389 14365 7423 14399
rect 9505 14365 9539 14399
rect 9781 14365 9815 14399
rect 9873 14365 9907 14399
rect 12173 14365 12207 14399
rect 14289 14365 14323 14399
rect 14565 14365 14599 14399
rect 14749 14365 14783 14399
rect 1676 14297 1710 14331
rect 5089 14297 5123 14331
rect 7297 14297 7331 14331
rect 7757 14297 7791 14331
rect 9321 14297 9355 14331
rect 10486 14297 10520 14331
rect 12418 14297 12452 14331
rect 17693 14501 17727 14535
rect 19533 14501 19567 14535
rect 24409 14501 24443 14535
rect 18521 14433 18555 14467
rect 29837 14433 29871 14467
rect 15577 14365 15611 14399
rect 15853 14365 15887 14399
rect 16037 14365 16071 14399
rect 16957 14365 16991 14399
rect 17233 14365 17267 14399
rect 17693 14365 17727 14399
rect 18337 14365 18371 14399
rect 18429 14365 18463 14399
rect 19349 14365 19383 14399
rect 20085 14365 20119 14399
rect 22477 14365 22511 14399
rect 22753 14365 22787 14399
rect 22937 14365 22971 14399
rect 23581 14365 23615 14399
rect 23765 14365 23799 14399
rect 23857 14365 23891 14399
rect 24593 14365 24627 14399
rect 24902 14365 24936 14399
rect 25065 14365 25099 14399
rect 25605 14365 25639 14399
rect 25697 14365 25731 14399
rect 25789 14365 25823 14399
rect 27169 14365 27203 14399
rect 27445 14365 27479 14399
rect 28733 14365 28767 14399
rect 28917 14365 28951 14399
rect 29009 14365 29043 14399
rect 30093 14365 30127 14399
rect 26525 14297 26559 14331
rect 26709 14297 26743 14331
rect 2789 14229 2823 14263
rect 3801 14229 3835 14263
rect 4169 14229 4203 14263
rect 5641 14229 5675 14263
rect 6101 14229 6135 14263
rect 7021 14229 7055 14263
rect 8125 14229 8159 14263
rect 9873 14229 9907 14263
rect 11621 14229 11655 14263
rect 15301 14229 15335 14263
rect 15393 14229 15427 14263
rect 17969 14229 18003 14263
rect 21373 14229 21407 14263
rect 22293 14229 22327 14263
rect 31217 14229 31251 14263
rect 2789 14025 2823 14059
rect 3893 14025 3927 14059
rect 4077 14025 4111 14059
rect 8217 14025 8251 14059
rect 8953 14025 8987 14059
rect 10333 14025 10367 14059
rect 14657 14025 14691 14059
rect 16681 14025 16715 14059
rect 21189 14025 21223 14059
rect 23213 14025 23247 14059
rect 26249 14025 26283 14059
rect 28825 14025 28859 14059
rect 29653 14025 29687 14059
rect 2145 13957 2179 13991
rect 3065 13957 3099 13991
rect 3157 13957 3191 13991
rect 3525 13957 3559 13991
rect 7021 13957 7055 13991
rect 14105 13957 14139 13991
rect 15301 13957 15335 13991
rect 17049 13957 17083 13991
rect 22078 13957 22112 13991
rect 23949 13957 23983 13991
rect 28457 13957 28491 13991
rect 28673 13957 28707 13991
rect 29929 13957 29963 13991
rect 1961 13889 1995 13923
rect 4905 13889 4939 13923
rect 6929 13889 6963 13923
rect 8677 13889 8711 13923
rect 8861 13889 8895 13923
rect 8953 13889 8987 13923
rect 9505 13889 9539 13923
rect 9689 13889 9723 13923
rect 10517 13889 10551 13923
rect 10793 13889 10827 13923
rect 10977 13889 11011 13923
rect 11989 13889 12023 13923
rect 12173 13889 12207 13923
rect 12909 13889 12943 13923
rect 13093 13889 13127 13923
rect 13369 13889 13403 13923
rect 13553 13889 13587 13923
rect 14013 13889 14047 13923
rect 14197 13889 14231 13923
rect 14289 13889 14323 13923
rect 14841 13889 14875 13923
rect 15117 13889 15151 13923
rect 1777 13821 1811 13855
rect 4629 13821 4663 13855
rect 7205 13821 7239 13855
rect 7757 13821 7791 13855
rect 9781 13821 9815 13855
rect 12357 13821 12391 13855
rect 12449 13821 12483 13855
rect 6561 13753 6595 13787
rect 8033 13753 8067 13787
rect 9321 13753 9355 13787
rect 15761 13889 15795 13923
rect 15945 13889 15979 13923
rect 17969 13889 18003 13923
rect 18236 13889 18270 13923
rect 19809 13889 19843 13923
rect 20065 13889 20099 13923
rect 16037 13821 16071 13855
rect 17141 13821 17175 13855
rect 17233 13821 17267 13855
rect 21833 13821 21867 13855
rect 24409 13889 24443 13923
rect 25145 13889 25179 13923
rect 25329 13889 25363 13923
rect 25605 13889 25639 13923
rect 25789 13889 25823 13923
rect 26433 13889 26467 13923
rect 27169 13889 27203 13923
rect 27445 13889 27479 13923
rect 29285 13889 29319 13923
rect 24593 13821 24627 13855
rect 24685 13821 24719 13855
rect 31125 13889 31159 13923
rect 31309 13889 31343 13923
rect 30297 13821 30331 13855
rect 30849 13821 30883 13855
rect 26985 13753 27019 13787
rect 27353 13753 27387 13787
rect 29837 13753 29871 13787
rect 29929 13753 29963 13787
rect 8677 13685 8711 13719
rect 14289 13685 14323 13719
rect 15025 13685 15059 13719
rect 15301 13685 15335 13719
rect 15577 13685 15611 13719
rect 19349 13685 19383 13719
rect 23949 13685 23983 13719
rect 24225 13685 24259 13719
rect 28641 13685 28675 13719
rect 29653 13685 29687 13719
rect 2697 13481 2731 13515
rect 3065 13481 3099 13515
rect 7113 13481 7147 13515
rect 7665 13481 7699 13515
rect 16589 13481 16623 13515
rect 17325 13481 17359 13515
rect 18429 13481 18463 13515
rect 19441 13481 19475 13515
rect 21833 13481 21867 13515
rect 22201 13481 22235 13515
rect 26157 13481 26191 13515
rect 26985 13481 27019 13515
rect 27629 13481 27663 13515
rect 28549 13481 28583 13515
rect 28825 13481 28859 13515
rect 29009 13481 29043 13515
rect 29929 13481 29963 13515
rect 30941 13481 30975 13515
rect 31125 13481 31159 13515
rect 4353 13413 4387 13447
rect 14197 13413 14231 13447
rect 15393 13413 15427 13447
rect 1409 13345 1443 13379
rect 3157 13345 3191 13379
rect 8125 13345 8159 13379
rect 8309 13345 8343 13379
rect 9413 13345 9447 13379
rect 16221 13345 16255 13379
rect 1685 13277 1719 13311
rect 2881 13277 2915 13311
rect 5825 13277 5859 13311
rect 7021 13277 7055 13311
rect 9137 13277 9171 13311
rect 10517 13277 10551 13311
rect 12541 13277 12575 13311
rect 12817 13277 12851 13311
rect 13001 13277 13035 13311
rect 14105 13277 14139 13311
rect 14289 13277 14323 13311
rect 15393 13277 15427 13311
rect 15577 13277 15611 13311
rect 16405 13277 16439 13311
rect 3985 13209 4019 13243
rect 5365 13209 5399 13243
rect 5457 13209 5491 13243
rect 10784 13209 10818 13243
rect 14841 13209 14875 13243
rect 15025 13209 15059 13243
rect 15761 13209 15795 13243
rect 17233 13209 17267 13243
rect 17969 13209 18003 13243
rect 19993 13345 20027 13379
rect 22293 13345 22327 13379
rect 24777 13345 24811 13379
rect 27077 13345 27111 13379
rect 27813 13345 27847 13379
rect 19349 13277 19383 13311
rect 22017 13277 22051 13311
rect 23397 13277 23431 13311
rect 23673 13277 23707 13311
rect 23857 13277 23891 13311
rect 25033 13277 25067 13311
rect 26801 13277 26835 13311
rect 27537 13277 27571 13311
rect 28549 13277 28583 13311
rect 29745 13277 29779 13311
rect 30021 13277 30055 13311
rect 20238 13209 20272 13243
rect 28641 13209 28675 13243
rect 30573 13209 30607 13243
rect 30950 13209 30984 13243
rect 4445 13141 4479 13175
rect 5089 13141 5123 13175
rect 6193 13141 6227 13175
rect 6377 13141 6411 13175
rect 8033 13141 8067 13175
rect 11897 13141 11931 13175
rect 12357 13141 12391 13175
rect 18245 13141 18279 13175
rect 18429 13141 18463 13175
rect 21373 13141 21407 13175
rect 23213 13141 23247 13175
rect 26617 13141 26651 13175
rect 27813 13141 27847 13175
rect 28841 13141 28875 13175
rect 29561 13141 29595 13175
rect 2145 12937 2179 12971
rect 4629 12937 4663 12971
rect 4813 12937 4847 12971
rect 5181 12937 5215 12971
rect 8033 12937 8067 12971
rect 26985 12937 27019 12971
rect 29653 12937 29687 12971
rect 1501 12869 1535 12903
rect 5273 12869 5307 12903
rect 14289 12869 14323 12903
rect 15016 12869 15050 12903
rect 18797 12869 18831 12903
rect 19441 12869 19475 12903
rect 2329 12801 2363 12835
rect 2605 12801 2639 12835
rect 2789 12801 2823 12835
rect 3433 12801 3467 12835
rect 3709 12801 3743 12835
rect 4353 12801 4387 12835
rect 4629 12801 4663 12835
rect 6377 12801 6411 12835
rect 7835 12801 7869 12835
rect 8585 12801 8619 12835
rect 8769 12801 8803 12835
rect 9505 12801 9539 12835
rect 9781 12801 9815 12835
rect 10241 12801 10275 12835
rect 11713 12801 11747 12835
rect 12541 12801 12575 12835
rect 12725 12801 12759 12835
rect 13277 12801 13311 12835
rect 13921 12801 13955 12835
rect 14105 12801 14139 12835
rect 14749 12801 14783 12835
rect 16773 12801 16807 12835
rect 16957 12801 16991 12835
rect 17049 12801 17083 12835
rect 17693 12801 17727 12835
rect 17969 12801 18003 12835
rect 18153 12801 18187 12835
rect 19625 12801 19659 12835
rect 20545 12801 20579 12835
rect 22017 12801 22051 12835
rect 23469 12801 23503 12835
rect 25053 12801 25087 12835
rect 25973 12801 26007 12835
rect 26249 12801 26283 12835
rect 26433 12801 26467 12835
rect 27169 12801 27203 12835
rect 27445 12801 27479 12835
rect 27629 12801 27663 12835
rect 28273 12801 28307 12835
rect 28540 12801 28574 12835
rect 30573 12801 30607 12835
rect 30849 12801 30883 12835
rect 5365 12733 5399 12767
rect 6653 12733 6687 12767
rect 7665 12733 7699 12767
rect 10149 12733 10183 12767
rect 11897 12733 11931 12767
rect 11989 12733 12023 12767
rect 19901 12733 19935 12767
rect 20821 12733 20855 12767
rect 21833 12733 21867 12767
rect 23213 12733 23247 12767
rect 25329 12733 25363 12767
rect 30757 12733 30791 12767
rect 1685 12665 1719 12699
rect 4169 12665 4203 12699
rect 16129 12665 16163 12699
rect 16773 12665 16807 12699
rect 20729 12665 20763 12699
rect 25145 12665 25179 12699
rect 3249 12597 3283 12631
rect 3617 12597 3651 12631
rect 9321 12597 9355 12631
rect 9689 12597 9723 12631
rect 10149 12597 10183 12631
rect 10425 12597 10459 12631
rect 11529 12597 11563 12631
rect 13369 12597 13403 12631
rect 17509 12597 17543 12631
rect 18889 12597 18923 12631
rect 19809 12597 19843 12631
rect 20361 12597 20395 12631
rect 22201 12597 22235 12631
rect 24593 12597 24627 12631
rect 25237 12597 25271 12631
rect 25789 12597 25823 12631
rect 30389 12597 30423 12631
rect 2789 12393 2823 12427
rect 5917 12393 5951 12427
rect 6745 12393 6779 12427
rect 13461 12393 13495 12427
rect 17693 12393 17727 12427
rect 19625 12393 19659 12427
rect 21649 12393 21683 12427
rect 23397 12393 23431 12427
rect 26157 12393 26191 12427
rect 28733 12393 28767 12427
rect 31309 12393 31343 12427
rect 21005 12325 21039 12359
rect 23765 12325 23799 12359
rect 4077 12257 4111 12291
rect 8309 12257 8343 12291
rect 8953 12257 8987 12291
rect 18705 12257 18739 12291
rect 29929 12257 29963 12291
rect 1409 12189 1443 12223
rect 4537 12189 4571 12223
rect 6469 12189 6503 12223
rect 6561 12189 6595 12223
rect 8033 12189 8067 12223
rect 9220 12189 9254 12223
rect 10793 12189 10827 12223
rect 11069 12189 11103 12223
rect 12725 12189 12759 12223
rect 13369 12189 13403 12223
rect 13553 12189 13587 12223
rect 14105 12189 14139 12223
rect 16313 12189 16347 12223
rect 18521 12189 18555 12223
rect 19809 12189 19843 12223
rect 20085 12189 20119 12223
rect 20269 12189 20303 12223
rect 21465 12189 21499 12223
rect 22569 12189 22603 12223
rect 23581 12189 23615 12223
rect 23857 12189 23891 12223
rect 24961 12189 24995 12223
rect 25145 12189 25179 12223
rect 25237 12189 25271 12223
rect 25973 12189 26007 12223
rect 26249 12189 26283 12223
rect 26709 12189 26743 12223
rect 26976 12189 27010 12223
rect 30196 12189 30230 12223
rect 1676 12121 1710 12155
rect 3893 12121 3927 12155
rect 4804 12121 4838 12155
rect 8125 12121 8159 12155
rect 14350 12121 14384 12155
rect 16580 12121 16614 12155
rect 20821 12121 20855 12155
rect 28549 12121 28583 12155
rect 7665 12053 7699 12087
rect 10333 12053 10367 12087
rect 12817 12053 12851 12087
rect 15485 12053 15519 12087
rect 22661 12053 22695 12087
rect 24777 12053 24811 12087
rect 25789 12053 25823 12087
rect 28089 12053 28123 12087
rect 28749 12053 28783 12087
rect 28917 12053 28951 12087
rect 6745 11849 6779 11883
rect 7941 11849 7975 11883
rect 10885 11849 10919 11883
rect 13185 11849 13219 11883
rect 14013 11849 14047 11883
rect 15485 11849 15519 11883
rect 23673 11849 23707 11883
rect 24501 11849 24535 11883
rect 25253 11849 25287 11883
rect 27445 11849 27479 11883
rect 28917 11849 28951 11883
rect 30297 11849 30331 11883
rect 1777 11781 1811 11815
rect 2942 11781 2976 11815
rect 6837 11781 6871 11815
rect 8033 11781 8067 11815
rect 10793 11781 10827 11815
rect 16865 11781 16899 11815
rect 21925 11781 21959 11815
rect 25053 11781 25087 11815
rect 27813 11781 27847 11815
rect 1961 11713 1995 11747
rect 4445 11713 4479 11747
rect 4813 11713 4847 11747
rect 5089 11713 5123 11747
rect 5273 11713 5307 11747
rect 8769 11713 8803 11747
rect 9413 11713 9447 11747
rect 12072 11713 12106 11747
rect 15301 11713 15335 11747
rect 17049 11713 17083 11747
rect 17233 11713 17267 11747
rect 18429 11713 18463 11747
rect 18705 11713 18739 11747
rect 18889 11713 18923 11747
rect 19349 11713 19383 11747
rect 19616 11713 19650 11747
rect 22753 11713 22787 11747
rect 23581 11713 23615 11747
rect 23805 11713 23839 11747
rect 23949 11713 23983 11747
rect 24409 11713 24443 11747
rect 25973 11713 26007 11747
rect 27629 11713 27663 11747
rect 27905 11713 27939 11747
rect 29101 11713 29135 11747
rect 29377 11713 29411 11747
rect 29561 11713 29595 11747
rect 30481 11713 30515 11747
rect 30757 11713 30791 11747
rect 30941 11713 30975 11747
rect 2237 11645 2271 11679
rect 2697 11645 2731 11679
rect 7021 11645 7055 11679
rect 8217 11645 8251 11679
rect 9689 11645 9723 11679
rect 11805 11645 11839 11679
rect 14105 11645 14139 11679
rect 14289 11645 14323 11679
rect 17325 11645 17359 11679
rect 23397 11645 23431 11679
rect 4077 11577 4111 11611
rect 4445 11577 4479 11611
rect 22109 11577 22143 11611
rect 22937 11577 22971 11611
rect 25421 11577 25455 11611
rect 2145 11509 2179 11543
rect 4629 11509 4663 11543
rect 6377 11509 6411 11543
rect 7573 11509 7607 11543
rect 8861 11509 8895 11543
rect 13645 11509 13679 11543
rect 18245 11509 18279 11543
rect 20729 11509 20763 11543
rect 25237 11509 25271 11543
rect 26065 11509 26099 11543
rect 2329 11305 2363 11339
rect 5089 11305 5123 11339
rect 7481 11305 7515 11339
rect 13001 11305 13035 11339
rect 17233 11305 17267 11339
rect 19533 11305 19567 11339
rect 24961 11305 24995 11339
rect 28917 11305 28951 11339
rect 31033 11305 31067 11339
rect 1869 11237 1903 11271
rect 5457 11237 5491 11271
rect 8769 11237 8803 11271
rect 8953 11237 8987 11271
rect 12909 11237 12943 11271
rect 28089 11237 28123 11271
rect 29101 11237 29135 11271
rect 4077 11169 4111 11203
rect 5549 11169 5583 11203
rect 1685 11101 1719 11135
rect 2513 11101 2547 11135
rect 2789 11101 2823 11135
rect 2973 11101 3007 11135
rect 3801 11101 3835 11135
rect 5273 11101 5307 11135
rect 8033 11101 8067 11135
rect 8217 11101 8251 11135
rect 6193 11033 6227 11067
rect 6469 11033 6503 11067
rect 6561 11033 6595 11067
rect 6929 11033 6963 11067
rect 7297 11033 7331 11067
rect 8401 11033 8435 11067
rect 9689 11169 9723 11203
rect 20177 11169 20211 11203
rect 20821 11169 20855 11203
rect 9229 11101 9263 11135
rect 9873 11101 9907 11135
rect 10149 11101 10183 11135
rect 10333 11101 10367 11135
rect 11437 11101 11471 11135
rect 14473 11101 14507 11135
rect 14729 11101 14763 11135
rect 17049 11101 17083 11135
rect 17325 11101 17359 11135
rect 18061 11101 18095 11135
rect 18153 11101 18187 11135
rect 18245 11101 18279 11135
rect 18429 11101 18463 11135
rect 19901 11101 19935 11135
rect 19993 11101 20027 11135
rect 22845 11101 22879 11135
rect 23121 11101 23155 11135
rect 23305 11101 23339 11135
rect 24869 11101 24903 11135
rect 25697 11101 25731 11135
rect 25881 11101 25915 11135
rect 25973 11101 26007 11135
rect 26709 11101 26743 11135
rect 26965 11101 26999 11135
rect 28733 11101 28767 11135
rect 29009 11101 29043 11135
rect 29561 11169 29595 11203
rect 31125 11169 31159 11203
rect 29745 11101 29779 11135
rect 30021 11101 30055 11135
rect 30205 11101 30239 11135
rect 30849 11101 30883 11135
rect 8953 11033 8987 11067
rect 9137 11033 9171 11067
rect 11621 11033 11655 11067
rect 12541 11033 12575 11067
rect 21088 11033 21122 11067
rect 22661 11033 22695 11067
rect 25513 11033 25547 11067
rect 28549 11033 28583 11067
rect 29101 11033 29135 11067
rect 30665 11033 30699 11067
rect 8769 10965 8803 10999
rect 15853 10965 15887 10999
rect 16865 10965 16899 10999
rect 17785 10965 17819 10999
rect 22201 10965 22235 10999
rect 5641 10761 5675 10795
rect 6745 10761 6779 10795
rect 8125 10761 8159 10795
rect 14197 10761 14231 10795
rect 20269 10761 20303 10795
rect 20545 10761 20579 10795
rect 23765 10761 23799 10795
rect 25513 10761 25547 10795
rect 28089 10761 28123 10795
rect 30113 10761 30147 10795
rect 30573 10761 30607 10795
rect 7757 10693 7791 10727
rect 7931 10693 7965 10727
rect 8493 10693 8527 10727
rect 10241 10693 10275 10727
rect 13277 10693 13311 10727
rect 13737 10693 13771 10727
rect 15853 10693 15887 10727
rect 20085 10693 20119 10727
rect 1961 10625 1995 10659
rect 2237 10625 2271 10659
rect 3341 10625 3375 10659
rect 4721 10625 4755 10659
rect 4997 10625 5031 10659
rect 5181 10625 5215 10659
rect 5825 10625 5859 10659
rect 7113 10625 7147 10659
rect 8217 10625 8251 10659
rect 21097 10693 21131 10727
rect 23489 10693 23523 10727
rect 29000 10693 29034 10727
rect 8677 10625 8711 10659
rect 9321 10625 9355 10659
rect 9505 10625 9539 10659
rect 10425 10625 10459 10659
rect 10701 10625 10735 10659
rect 10885 10625 10919 10659
rect 10977 10625 11011 10659
rect 11713 10625 11747 10659
rect 13093 10625 13127 10659
rect 15025 10625 15059 10659
rect 15209 10625 15243 10659
rect 16037 10625 16071 10659
rect 16129 10625 16163 10659
rect 16865 10625 16899 10659
rect 17049 10625 17083 10659
rect 17141 10625 17175 10659
rect 18133 10625 18167 10659
rect 19717 10625 19751 10659
rect 20545 10625 20579 10659
rect 20913 10625 20947 10659
rect 21189 10625 21223 10659
rect 22017 10625 22051 10659
rect 22293 10625 22327 10659
rect 22477 10625 22511 10659
rect 24409 10625 24443 10659
rect 25697 10625 25731 10659
rect 25973 10625 26007 10659
rect 26157 10625 26191 10659
rect 27169 10625 27203 10659
rect 27445 10625 27479 10659
rect 27629 10625 27663 10659
rect 28273 10625 28307 10659
rect 30757 10625 30791 10659
rect 31033 10625 31067 10659
rect 31217 10625 31251 10659
rect 2145 10557 2179 10591
rect 3157 10557 3191 10591
rect 3249 10557 3283 10591
rect 3433 10557 3467 10591
rect 7205 10557 7239 10591
rect 7297 10557 7331 10591
rect 7849 10557 7883 10591
rect 8493 10557 8527 10591
rect 8953 10489 8987 10523
rect 11989 10557 12023 10591
rect 16681 10557 16715 10591
rect 17877 10557 17911 10591
rect 23121 10557 23155 10591
rect 23397 10557 23431 10591
rect 23606 10557 23640 10591
rect 24685 10557 24719 10591
rect 28733 10557 28767 10591
rect 14105 10489 14139 10523
rect 15393 10489 15427 10523
rect 15853 10489 15887 10523
rect 20729 10489 20763 10523
rect 1777 10421 1811 10455
rect 2973 10421 3007 10455
rect 4537 10421 4571 10455
rect 7941 10421 7975 10455
rect 10977 10421 11011 10455
rect 11529 10421 11563 10455
rect 11897 10421 11931 10455
rect 19257 10421 19291 10455
rect 20085 10421 20119 10455
rect 21833 10421 21867 10455
rect 24225 10421 24259 10455
rect 24593 10421 24627 10455
rect 26985 10421 27019 10455
rect 5549 10217 5583 10251
rect 6745 10217 6779 10251
rect 7205 10217 7239 10251
rect 8217 10217 8251 10251
rect 8401 10217 8435 10251
rect 11161 10217 11195 10251
rect 13185 10217 13219 10251
rect 18061 10217 18095 10251
rect 21281 10217 21315 10251
rect 27629 10217 27663 10251
rect 31217 10217 31251 10251
rect 6561 10149 6595 10183
rect 7849 10149 7883 10183
rect 18613 10149 18647 10183
rect 20269 10149 20303 10183
rect 16313 10081 16347 10115
rect 22017 10081 22051 10115
rect 1409 10013 1443 10047
rect 4169 10013 4203 10047
rect 7389 10013 7423 10047
rect 9781 10013 9815 10047
rect 11805 10013 11839 10047
rect 16681 10013 16715 10047
rect 16937 10013 16971 10047
rect 18521 10013 18555 10047
rect 20085 10013 20119 10047
rect 21281 10013 21315 10047
rect 21557 10013 21591 10047
rect 24409 10013 24443 10047
rect 26249 10013 26283 10047
rect 28825 10013 28859 10047
rect 29837 10013 29871 10047
rect 30104 10013 30138 10047
rect 1676 9945 1710 9979
rect 4436 9945 4470 9979
rect 6285 9945 6319 9979
rect 8217 9945 8251 9979
rect 9137 9945 9171 9979
rect 10048 9945 10082 9979
rect 12072 9945 12106 9979
rect 14473 9945 14507 9979
rect 16313 9945 16347 9979
rect 19349 9945 19383 9979
rect 21465 9945 21499 9979
rect 22284 9945 22318 9979
rect 24654 9945 24688 9979
rect 26494 9945 26528 9979
rect 2789 9877 2823 9911
rect 9229 9877 9263 9911
rect 15761 9877 15795 9911
rect 19441 9877 19475 9911
rect 23397 9877 23431 9911
rect 25789 9877 25823 9911
rect 28641 9877 28675 9911
rect 5549 9673 5583 9707
rect 9137 9673 9171 9707
rect 22753 9673 22787 9707
rect 26341 9673 26375 9707
rect 1501 9605 1535 9639
rect 4905 9605 4939 9639
rect 1409 9537 1443 9571
rect 2053 9537 2087 9571
rect 3525 9537 3559 9571
rect 4077 9537 4111 9571
rect 5089 9537 5123 9571
rect 5365 9537 5399 9571
rect 2329 9469 2363 9503
rect 4169 9469 4203 9503
rect 7205 9605 7239 9639
rect 8309 9605 8343 9639
rect 8769 9605 8803 9639
rect 7113 9537 7147 9571
rect 7389 9469 7423 9503
rect 8401 9469 8435 9503
rect 8585 9469 8619 9503
rect 3617 9401 3651 9435
rect 5549 9401 5583 9435
rect 6745 9401 6779 9435
rect 8861 9605 8895 9639
rect 14372 9605 14406 9639
rect 24501 9605 24535 9639
rect 25228 9605 25262 9639
rect 10701 9537 10735 9571
rect 10973 9537 11007 9571
rect 11529 9537 11563 9571
rect 11713 9537 11747 9571
rect 11989 9537 12023 9571
rect 12173 9537 12207 9571
rect 13277 9537 13311 9571
rect 14105 9537 14139 9571
rect 16129 9537 16163 9571
rect 16865 9537 16899 9571
rect 18245 9537 18279 9571
rect 18429 9537 18463 9571
rect 20361 9537 20395 9571
rect 20637 9537 20671 9571
rect 20821 9537 20855 9571
rect 22017 9537 22051 9571
rect 22293 9537 22327 9571
rect 22937 9537 22971 9571
rect 23213 9537 23247 9571
rect 24317 9537 24351 9571
rect 27169 9537 27203 9571
rect 27629 9537 27663 9571
rect 27885 9537 27919 9571
rect 29469 9537 29503 9571
rect 31309 9537 31343 9571
rect 8861 9469 8895 9503
rect 9321 9469 9355 9503
rect 9413 9469 9447 9503
rect 9505 9469 9539 9503
rect 9597 9469 9631 9503
rect 17141 9469 17175 9503
rect 18153 9469 18187 9503
rect 18337 9469 18371 9503
rect 18981 9469 19015 9503
rect 24869 9469 24903 9503
rect 24961 9469 24995 9503
rect 29745 9469 29779 9503
rect 13553 9401 13587 9435
rect 15945 9401 15979 9435
rect 19257 9401 19291 9435
rect 21833 9401 21867 9435
rect 24685 9401 24719 9435
rect 5273 9333 5307 9367
rect 7941 9333 7975 9367
rect 8769 9333 8803 9367
rect 10517 9333 10551 9367
rect 10885 9333 10919 9367
rect 15485 9333 15519 9367
rect 16681 9333 16715 9367
rect 17049 9333 17083 9367
rect 17969 9333 18003 9367
rect 19441 9333 19475 9367
rect 20177 9333 20211 9367
rect 22201 9333 22235 9367
rect 23121 9333 23155 9367
rect 26985 9333 27019 9367
rect 29009 9333 29043 9367
rect 31125 9333 31159 9367
rect 4169 9129 4203 9163
rect 4445 9129 4479 9163
rect 2513 8993 2547 9027
rect 2973 8993 3007 9027
rect 2329 8925 2363 8959
rect 3801 8925 3835 8959
rect 2421 8857 2455 8891
rect 2973 8857 3007 8891
rect 5549 9129 5583 9163
rect 8217 9129 8251 9163
rect 25145 9129 25179 9163
rect 26157 9129 26191 9163
rect 27445 9129 27479 9163
rect 27813 9129 27847 9163
rect 30481 9129 30515 9163
rect 11897 9061 11931 9095
rect 13001 9061 13035 9095
rect 17509 9061 17543 9095
rect 18429 9061 18463 9095
rect 21649 9061 21683 9095
rect 23121 9061 23155 9095
rect 26525 9061 26559 9095
rect 5549 8993 5583 9027
rect 6377 8993 6411 9027
rect 10517 8993 10551 9027
rect 12633 8993 12667 9027
rect 14657 8993 14691 9027
rect 16957 8993 16991 9027
rect 26617 8993 26651 9027
rect 28365 8993 28399 9027
rect 30021 8993 30055 9027
rect 4997 8925 5031 8959
rect 5273 8925 5307 8959
rect 5457 8925 5491 8959
rect 6101 8925 6135 8959
rect 6285 8925 6319 8959
rect 6929 8925 6963 8959
rect 7205 8925 7239 8959
rect 8401 8925 8435 8959
rect 8769 8925 8803 8959
rect 9229 8925 9263 8959
rect 9321 8925 9355 8959
rect 9505 8925 9539 8959
rect 9965 8925 9999 8959
rect 10773 8925 10807 8959
rect 14924 8925 14958 8959
rect 16681 8925 16715 8959
rect 16865 8925 16899 8959
rect 17417 8925 17451 8959
rect 17601 8925 17635 8959
rect 18245 8925 18279 8959
rect 18521 8925 18555 8959
rect 19533 8925 19567 8959
rect 19717 8925 19751 8959
rect 19809 8925 19843 8959
rect 20085 8925 20119 8959
rect 20269 8925 20303 8959
rect 23121 8925 23155 8959
rect 23397 8925 23431 8959
rect 26341 8925 26375 8959
rect 27629 8925 27663 8959
rect 27905 8925 27939 8959
rect 28549 8925 28583 8959
rect 28825 8925 28859 8959
rect 29009 8925 29043 8959
rect 29745 8925 29779 8959
rect 29929 8925 29963 8959
rect 30665 8925 30699 8959
rect 31309 8925 31343 8959
rect 4813 8857 4847 8891
rect 5917 8857 5951 8891
rect 1961 8789 1995 8823
rect 4169 8789 4203 8823
rect 4353 8789 4387 8823
rect 4445 8789 4479 8823
rect 19349 8857 19383 8891
rect 20514 8857 20548 8891
rect 22293 8857 22327 8891
rect 22661 8857 22695 8891
rect 22845 8857 22879 8891
rect 24961 8857 24995 8891
rect 8769 8789 8803 8823
rect 13093 8789 13127 8823
rect 16037 8789 16071 8823
rect 16497 8789 16531 8823
rect 18061 8789 18095 8823
rect 20085 8789 20119 8823
rect 23029 8789 23063 8823
rect 23305 8789 23339 8823
rect 25161 8789 25195 8823
rect 25329 8789 25363 8823
rect 29561 8789 29595 8823
rect 31125 8789 31159 8823
rect 5549 8585 5583 8619
rect 7757 8585 7791 8619
rect 8217 8585 8251 8619
rect 8585 8585 8619 8619
rect 1869 8517 1903 8551
rect 3065 8517 3099 8551
rect 3433 8517 3467 8551
rect 9781 8517 9815 8551
rect 11621 8517 11655 8551
rect 16926 8517 16960 8551
rect 21833 8517 21867 8551
rect 23949 8517 23983 8551
rect 24165 8517 24199 8551
rect 28641 8517 28675 8551
rect 2053 8449 2087 8483
rect 2145 8449 2179 8483
rect 2973 8449 3007 8483
rect 3249 8381 3283 8415
rect 4169 8449 4203 8483
rect 4436 8449 4470 8483
rect 6633 8449 6667 8483
rect 10609 8449 10643 8483
rect 12357 8449 12391 8483
rect 13001 8449 13035 8483
rect 13268 8449 13302 8483
rect 18981 8449 19015 8483
rect 19165 8449 19199 8483
rect 19441 8449 19475 8483
rect 19637 8449 19671 8483
rect 20269 8449 20303 8483
rect 20545 8449 20579 8483
rect 20729 8449 20763 8483
rect 22661 8449 22695 8483
rect 23305 8449 23339 8483
rect 24869 8449 24903 8483
rect 25237 8449 25271 8483
rect 25421 8449 25455 8483
rect 25697 8449 25731 8483
rect 26157 8449 26191 8483
rect 27077 8449 27111 8483
rect 27905 8449 27939 8483
rect 31033 8449 31067 8483
rect 6377 8381 6411 8415
rect 8677 8381 8711 8415
rect 8861 8381 8895 8415
rect 9413 8381 9447 8415
rect 10885 8381 10919 8415
rect 12541 8381 12575 8415
rect 15301 8381 15335 8415
rect 15577 8381 15611 8415
rect 16681 8381 16715 8415
rect 22385 8381 22419 8415
rect 22845 8381 22879 8415
rect 1869 8313 1903 8347
rect 3433 8313 3467 8347
rect 9965 8313 9999 8347
rect 10425 8313 10459 8347
rect 10793 8313 10827 8347
rect 11805 8313 11839 8347
rect 14381 8313 14415 8347
rect 18061 8313 18095 8347
rect 20085 8313 20119 8347
rect 23397 8313 23431 8347
rect 24317 8313 24351 8347
rect 24869 8313 24903 8347
rect 28181 8381 28215 8415
rect 31309 8381 31343 8415
rect 25697 8313 25731 8347
rect 26341 8313 26375 8347
rect 28089 8313 28123 8347
rect 30849 8313 30883 8347
rect 31217 8313 31251 8347
rect 2605 8245 2639 8279
rect 9781 8245 9815 8279
rect 24133 8245 24167 8279
rect 25605 8245 25639 8279
rect 27169 8245 27203 8279
rect 27721 8245 27755 8279
rect 29929 8245 29963 8279
rect 32137 8109 32171 8143
rect 3801 8041 3835 8075
rect 8217 8041 8251 8075
rect 8953 8041 8987 8075
rect 11161 8041 11195 8075
rect 13461 8041 13495 8075
rect 15393 8041 15427 8075
rect 18429 8041 18463 8075
rect 20729 8041 20763 8075
rect 21649 8041 21683 8075
rect 21833 8041 21867 8075
rect 27077 8041 27111 8075
rect 30941 8041 30975 8075
rect 8033 7973 8067 8007
rect 9965 7973 9999 8007
rect 4261 7905 4295 7939
rect 7757 7905 7791 7939
rect 11069 7973 11103 8007
rect 12725 7973 12759 8007
rect 26525 7973 26559 8007
rect 24777 7905 24811 7939
rect 25145 7905 25179 7939
rect 27813 7905 27847 7939
rect 28227 7905 28261 7939
rect 1593 7837 1627 7871
rect 2237 7837 2271 7871
rect 2513 7837 2547 7871
rect 2697 7837 2731 7871
rect 3985 7837 4019 7871
rect 4169 7837 4203 7871
rect 4905 7837 4939 7871
rect 5181 7837 5215 7871
rect 5365 7837 5399 7871
rect 6193 7837 6227 7871
rect 6469 7837 6503 7871
rect 6653 7837 6687 7871
rect 7297 7837 7331 7871
rect 9137 7837 9171 7871
rect 9413 7837 9447 7871
rect 9965 7837 9999 7871
rect 10241 7837 10275 7871
rect 10517 7837 10551 7871
rect 10701 7837 10735 7871
rect 11069 7837 11103 7871
rect 11345 7837 11379 7871
rect 11621 7837 11655 7871
rect 11805 7837 11839 7871
rect 12541 7837 12575 7871
rect 12817 7837 12851 7871
rect 13369 7837 13403 7871
rect 14105 7837 14139 7871
rect 14381 7837 14415 7871
rect 15577 7837 15611 7871
rect 15853 7837 15887 7871
rect 16037 7837 16071 7871
rect 17049 7837 17083 7871
rect 19349 7837 19383 7871
rect 21281 7837 21315 7871
rect 22385 7837 22419 7871
rect 24961 7837 24995 7871
rect 25605 7837 25639 7871
rect 25789 7837 25823 7871
rect 27077 7837 27111 7871
rect 27169 7837 27203 7871
rect 27353 7837 27387 7871
rect 28089 7837 28123 7871
rect 28365 7837 28399 7871
rect 29561 7837 29595 7871
rect 29828 7837 29862 7871
rect 6009 7769 6043 7803
rect 9321 7769 9355 7803
rect 17316 7769 17350 7803
rect 19594 7769 19628 7803
rect 22630 7769 22664 7803
rect 26249 7769 26283 7803
rect 1409 7701 1443 7735
rect 2053 7701 2087 7735
rect 4721 7701 4755 7735
rect 7113 7701 7147 7735
rect 9965 7701 9999 7735
rect 10057 7701 10091 7735
rect 12357 7701 12391 7735
rect 21658 7701 21692 7735
rect 23765 7701 23799 7735
rect 25697 7701 25731 7735
rect 26709 7701 26743 7735
rect 29009 7701 29043 7735
rect 2053 7497 2087 7531
rect 6193 7497 6227 7531
rect 6377 7497 6411 7531
rect 8769 7497 8803 7531
rect 10977 7497 11011 7531
rect 14565 7497 14599 7531
rect 15669 7497 15703 7531
rect 16681 7497 16715 7531
rect 21097 7497 21131 7531
rect 22201 7497 22235 7531
rect 22385 7497 22419 7531
rect 29285 7497 29319 7531
rect 31309 7497 31343 7531
rect 1593 7361 1627 7395
rect 2237 7361 2271 7395
rect 2513 7361 2547 7395
rect 2697 7361 2731 7395
rect 3709 7361 3743 7395
rect 3985 7361 4019 7395
rect 4169 7361 4203 7395
rect 5365 7361 5399 7395
rect 5641 7361 5675 7395
rect 5825 7361 5859 7395
rect 11888 7429 11922 7463
rect 26985 7429 27019 7463
rect 30196 7429 30230 7463
rect 6561 7361 6595 7395
rect 6745 7361 6779 7395
rect 6837 7361 6871 7395
rect 7389 7361 7423 7395
rect 7656 7361 7690 7395
rect 9597 7361 9631 7395
rect 9864 7361 9898 7395
rect 11621 7361 11655 7395
rect 13645 7361 13679 7395
rect 13921 7361 13955 7395
rect 14105 7361 14139 7395
rect 14749 7361 14783 7395
rect 15025 7361 15059 7395
rect 15209 7361 15243 7395
rect 15853 7361 15887 7395
rect 16037 7361 16071 7395
rect 16865 7361 16899 7395
rect 17141 7361 17175 7395
rect 17325 7361 17359 7395
rect 18061 7361 18095 7395
rect 18328 7361 18362 7395
rect 20269 7361 20303 7395
rect 21281 7361 21315 7395
rect 23673 7361 23707 7395
rect 23765 7361 23799 7395
rect 24409 7361 24443 7395
rect 26065 7361 26099 7395
rect 26157 7361 26191 7395
rect 27905 7361 27939 7395
rect 28161 7361 28195 7395
rect 16129 7293 16163 7327
rect 20361 7293 20395 7327
rect 20545 7293 20579 7327
rect 21833 7293 21867 7327
rect 24501 7293 24535 7327
rect 26249 7293 26283 7327
rect 29929 7293 29963 7327
rect 6193 7225 6227 7259
rect 13001 7225 13035 7259
rect 24777 7225 24811 7259
rect 27353 7225 27387 7259
rect 1409 7157 1443 7191
rect 3525 7157 3559 7191
rect 5181 7157 5215 7191
rect 13461 7157 13495 7191
rect 19441 7157 19475 7191
rect 19901 7157 19935 7191
rect 22201 7157 22235 7191
rect 25697 7157 25731 7191
rect 27445 7157 27479 7191
rect 8125 6953 8159 6987
rect 10241 6953 10275 6987
rect 19349 6953 19383 6987
rect 21649 6953 21683 6987
rect 22569 6953 22603 6987
rect 22753 6953 22787 6987
rect 23581 6953 23615 6987
rect 23765 6953 23799 6987
rect 2789 6885 2823 6919
rect 12725 6885 12759 6919
rect 32137 6885 32171 6919
rect 4169 6817 4203 6851
rect 4261 6817 4295 6851
rect 8953 6817 8987 6851
rect 9229 6817 9263 6851
rect 10701 6817 10735 6851
rect 11345 6817 11379 6851
rect 13461 6817 13495 6851
rect 14565 6817 14599 6851
rect 15025 6817 15059 6851
rect 15301 6817 15335 6851
rect 15418 6817 15452 6851
rect 15577 6817 15611 6851
rect 16773 6817 16807 6851
rect 18061 6817 18095 6851
rect 19717 6817 19751 6851
rect 25513 6817 25547 6851
rect 25605 6817 25639 6851
rect 27169 6817 27203 6851
rect 28365 6817 28399 6851
rect 29745 6817 29779 6851
rect 31309 6817 31343 6851
rect 1409 6749 1443 6783
rect 3985 6749 4019 6783
rect 5089 6749 5123 6783
rect 5365 6749 5399 6783
rect 10425 6749 10459 6783
rect 10609 6749 10643 6783
rect 14381 6749 14415 6783
rect 16221 6749 16255 6783
rect 16957 6749 16991 6783
rect 17141 6749 17175 6783
rect 17233 6749 17267 6783
rect 17877 6749 17911 6783
rect 18153 6749 18187 6783
rect 19533 6749 19567 6783
rect 19809 6749 19843 6783
rect 20269 6749 20303 6783
rect 23213 6749 23247 6783
rect 24593 6749 24627 6783
rect 28089 6749 28123 6783
rect 29929 6749 29963 6783
rect 30205 6749 30239 6783
rect 30389 6749 30423 6783
rect 31033 6749 31067 6783
rect 31217 6749 31251 6783
rect 1676 6681 1710 6715
rect 6653 6681 6687 6715
rect 11612 6681 11646 6715
rect 13277 6681 13311 6715
rect 20536 6681 20570 6715
rect 22385 6681 22419 6715
rect 22601 6681 22635 6715
rect 25421 6681 25455 6715
rect 26985 6681 27019 6715
rect 3801 6613 3835 6647
rect 17693 6613 17727 6647
rect 23590 6613 23624 6647
rect 24409 6613 24443 6647
rect 25053 6613 25087 6647
rect 26617 6613 26651 6647
rect 27077 6613 27111 6647
rect 30849 6613 30883 6647
rect 1777 6409 1811 6443
rect 4537 6409 4571 6443
rect 5641 6409 5675 6443
rect 10333 6409 10367 6443
rect 12265 6409 12299 6443
rect 14933 6409 14967 6443
rect 16681 6409 16715 6443
rect 19717 6409 19751 6443
rect 27721 6409 27755 6443
rect 30481 6409 30515 6443
rect 3249 6341 3283 6375
rect 9229 6341 9263 6375
rect 15853 6341 15887 6375
rect 1961 6273 1995 6307
rect 2237 6273 2271 6307
rect 5457 6273 5491 6307
rect 5733 6273 5767 6307
rect 7941 6273 7975 6307
rect 8217 6273 8251 6307
rect 9413 6273 9447 6307
rect 9689 6273 9723 6307
rect 9873 6273 9907 6307
rect 10517 6273 10551 6307
rect 10793 6273 10827 6307
rect 11621 6273 11655 6307
rect 12449 6273 12483 6307
rect 13829 6273 13863 6307
rect 14105 6273 14139 6307
rect 14289 6273 14323 6307
rect 14749 6273 14783 6307
rect 15577 6273 15611 6307
rect 15761 6273 15795 6307
rect 15945 6273 15979 6307
rect 16957 6273 16991 6307
rect 17049 6273 17083 6307
rect 17141 6273 17175 6307
rect 17325 6273 17359 6307
rect 17785 6273 17819 6307
rect 18429 6273 18463 6307
rect 22477 6273 22511 6307
rect 23673 6273 23707 6307
rect 24409 6273 24443 6307
rect 24593 6273 24627 6307
rect 24869 6273 24903 6307
rect 25053 6273 25087 6307
rect 25605 6273 25639 6307
rect 25789 6273 25823 6307
rect 25881 6273 25915 6307
rect 25973 6273 26007 6307
rect 26985 6273 27019 6307
rect 27169 6273 27203 6307
rect 27261 6273 27295 6307
rect 27399 6273 27433 6307
rect 2145 6205 2179 6239
rect 6653 6205 6687 6239
rect 6929 6205 6963 6239
rect 12633 6205 12667 6239
rect 12725 6205 12759 6239
rect 12817 6205 12851 6239
rect 13645 6205 13679 6239
rect 17877 6205 17911 6239
rect 20637 6205 20671 6239
rect 22753 6205 22787 6239
rect 23949 6205 23983 6239
rect 28181 6273 28215 6307
rect 29193 6273 29227 6307
rect 30665 6273 30699 6307
rect 30941 6273 30975 6307
rect 31125 6273 31159 6307
rect 29469 6205 29503 6239
rect 20913 6137 20947 6171
rect 27721 6137 27755 6171
rect 28365 6137 28399 6171
rect 5457 6069 5491 6103
rect 10701 6069 10735 6103
rect 11713 6069 11747 6103
rect 12817 6069 12851 6103
rect 16129 6069 16163 6103
rect 21097 6069 21131 6103
rect 22293 6069 22327 6103
rect 22661 6069 22695 6103
rect 23489 6069 23523 6103
rect 23857 6069 23891 6103
rect 26157 6069 26191 6103
rect 27537 6069 27571 6103
rect 1593 5865 1627 5899
rect 1961 5865 1995 5899
rect 25973 5865 26007 5899
rect 27721 5865 27755 5899
rect 29929 5865 29963 5899
rect 30481 5865 30515 5899
rect 2329 5797 2363 5831
rect 3157 5797 3191 5831
rect 4721 5797 4755 5831
rect 6469 5797 6503 5831
rect 8401 5797 8435 5831
rect 11529 5797 11563 5831
rect 13001 5797 13035 5831
rect 14657 5797 14691 5831
rect 16589 5797 16623 5831
rect 18245 5797 18279 5831
rect 20637 5797 20671 5831
rect 26433 5797 26467 5831
rect 2789 5729 2823 5763
rect 4353 5729 4387 5763
rect 1409 5661 1443 5695
rect 4169 5661 4203 5695
rect 7481 5729 7515 5763
rect 9505 5729 9539 5763
rect 10149 5729 10183 5763
rect 17877 5729 17911 5763
rect 5089 5661 5123 5695
rect 8217 5661 8251 5695
rect 9413 5661 9447 5695
rect 10416 5661 10450 5695
rect 11989 5661 12023 5695
rect 12173 5661 12207 5695
rect 12817 5661 12851 5695
rect 13093 5661 13127 5695
rect 14841 5661 14875 5695
rect 14933 5661 14967 5695
rect 15117 5661 15151 5695
rect 15209 5661 15243 5695
rect 15301 5661 15335 5695
rect 15669 5661 15703 5695
rect 15853 5661 15887 5695
rect 16773 5661 16807 5695
rect 17049 5661 17083 5695
rect 17233 5661 17267 5695
rect 19257 5661 19291 5695
rect 21833 5661 21867 5695
rect 22100 5661 22134 5695
rect 24593 5661 24627 5695
rect 26617 5661 26651 5695
rect 26709 5661 26743 5695
rect 27084 5661 27118 5695
rect 27225 5661 27259 5695
rect 27542 5661 27576 5695
rect 28549 5661 28583 5695
rect 28825 5661 28859 5695
rect 29009 5661 29043 5695
rect 29745 5661 29779 5695
rect 29929 5661 29963 5695
rect 30665 5661 30699 5695
rect 30941 5661 30975 5695
rect 31125 5661 31159 5695
rect 2145 5593 2179 5627
rect 4721 5593 4755 5627
rect 5356 5593 5390 5627
rect 7297 5593 7331 5627
rect 7389 5593 7423 5627
rect 9321 5593 9355 5627
rect 12081 5593 12115 5627
rect 19524 5593 19558 5627
rect 21189 5593 21223 5627
rect 24838 5593 24872 5627
rect 27353 5593 27387 5627
rect 27445 5593 27479 5627
rect 3249 5525 3283 5559
rect 3801 5525 3835 5559
rect 4261 5525 4295 5559
rect 6929 5525 6963 5559
rect 8953 5525 8987 5559
rect 12633 5525 12667 5559
rect 15301 5525 15335 5559
rect 16037 5525 16071 5559
rect 18337 5525 18371 5559
rect 21281 5525 21315 5559
rect 23213 5525 23247 5559
rect 26709 5525 26743 5559
rect 28365 5525 28399 5559
rect 29561 5525 29595 5559
rect 5365 5321 5399 5355
rect 7757 5321 7791 5355
rect 9045 5321 9079 5355
rect 27169 5321 27203 5355
rect 4721 5253 4755 5287
rect 4905 5253 4939 5287
rect 8125 5253 8159 5287
rect 8493 5253 8527 5287
rect 8861 5253 8895 5287
rect 17049 5253 17083 5287
rect 18420 5253 18454 5287
rect 20913 5253 20947 5287
rect 21113 5253 21147 5287
rect 24194 5253 24228 5287
rect 26157 5253 26191 5287
rect 2053 5185 2087 5219
rect 2237 5185 2271 5219
rect 2789 5185 2823 5219
rect 3056 5185 3090 5219
rect 5549 5185 5583 5219
rect 6377 5185 6411 5219
rect 6561 5185 6595 5219
rect 6837 5185 6871 5219
rect 7021 5185 7055 5219
rect 8033 5185 8067 5219
rect 11989 5185 12023 5219
rect 14013 5185 14047 5219
rect 14197 5185 14231 5219
rect 14473 5185 14507 5219
rect 14657 5185 14691 5219
rect 15485 5185 15519 5219
rect 15577 5185 15611 5219
rect 16681 5185 16715 5219
rect 16773 5185 16807 5219
rect 16957 5185 16991 5219
rect 17141 5185 17175 5219
rect 20177 5185 20211 5219
rect 22273 5185 22307 5219
rect 23949 5185 23983 5219
rect 25789 5185 25823 5219
rect 25882 5185 25916 5219
rect 26065 5185 26099 5219
rect 26295 5185 26329 5219
rect 26985 5185 27019 5219
rect 27988 5185 28022 5219
rect 30196 5185 30230 5219
rect 2329 5117 2363 5151
rect 5825 5117 5859 5151
rect 6193 5117 6227 5151
rect 9597 5117 9631 5151
rect 9873 5117 9907 5151
rect 12265 5117 12299 5151
rect 12725 5117 12759 5151
rect 13001 5117 13035 5151
rect 15117 5117 15151 5151
rect 15301 5117 15335 5151
rect 15393 5117 15427 5151
rect 18153 5117 18187 5151
rect 20453 5117 20487 5151
rect 22017 5117 22051 5151
rect 27721 5117 27755 5151
rect 29929 5117 29963 5151
rect 12173 5049 12207 5083
rect 16681 5049 16715 5083
rect 23397 5049 23431 5083
rect 26433 5049 26467 5083
rect 1869 4981 1903 5015
rect 4169 4981 4203 5015
rect 5733 4981 5767 5015
rect 6193 4981 6227 5015
rect 11805 4981 11839 5015
rect 17325 4981 17359 5015
rect 19533 4981 19567 5015
rect 19993 4981 20027 5015
rect 20361 4981 20395 5015
rect 21097 4981 21131 5015
rect 21281 4981 21315 5015
rect 25329 4981 25363 5015
rect 29101 4981 29135 5015
rect 31309 4981 31343 5015
rect 2789 4777 2823 4811
rect 7941 4777 7975 4811
rect 18153 4777 18187 4811
rect 7757 4709 7791 4743
rect 12909 4709 12943 4743
rect 15945 4709 15979 4743
rect 19533 4777 19567 4811
rect 20821 4777 20855 4811
rect 19257 4709 19291 4743
rect 1409 4641 1443 4675
rect 11529 4641 11563 4675
rect 13461 4641 13495 4675
rect 13645 4641 13679 4675
rect 14381 4641 14415 4675
rect 18153 4641 18187 4675
rect 18245 4641 18279 4675
rect 18613 4641 18647 4675
rect 1676 4573 1710 4607
rect 4353 4573 4387 4607
rect 6193 4573 6227 4607
rect 6469 4573 6503 4607
rect 6653 4573 6687 4607
rect 9505 4573 9539 4607
rect 11796 4573 11830 4607
rect 13369 4573 13403 4607
rect 13553 4573 13587 4607
rect 949 4505 983 4539
rect 3985 4505 4019 4539
rect 4261 4505 4295 4539
rect 4721 4505 4755 4539
rect 7481 4505 7515 4539
rect 9772 4505 9806 4539
rect 20269 4641 20303 4675
rect 20361 4641 20395 4675
rect 21281 4641 21315 4675
rect 23489 4641 23523 4675
rect 24593 4641 24627 4675
rect 24869 4641 24903 4675
rect 26525 4641 26559 4675
rect 28181 4641 28215 4675
rect 29561 4641 29595 4675
rect 14105 4573 14139 4607
rect 15413 4573 15447 4607
rect 15669 4573 15703 4607
rect 15807 4573 15841 4607
rect 16957 4573 16991 4607
rect 17233 4573 17267 4607
rect 18489 4573 18523 4607
rect 18701 4573 18735 4607
rect 18889 4573 18923 4607
rect 19257 4573 19291 4607
rect 19441 4573 19475 4607
rect 19533 4573 19567 4607
rect 20085 4573 20119 4607
rect 21005 4573 21039 4607
rect 21189 4573 21223 4607
rect 21741 4573 21775 4607
rect 26249 4573 26283 4607
rect 27721 4573 27755 4607
rect 28457 4573 28491 4607
rect 15577 4505 15611 4539
rect 5089 4437 5123 4471
rect 5273 4437 5307 4471
rect 6009 4437 6043 4471
rect 10885 4437 10919 4471
rect 13645 4437 13679 4471
rect 29806 4505 29840 4539
rect 18889 4437 18923 4471
rect 19901 4437 19935 4471
rect 27537 4437 27571 4471
rect 30941 4437 30975 4471
rect 1961 4233 1995 4267
rect 3065 4233 3099 4267
rect 6745 4233 6779 4267
rect 10333 4233 10367 4267
rect 15117 4233 15151 4267
rect 17601 4233 17635 4267
rect 18153 4233 18187 4267
rect 21281 4233 21315 4267
rect 29377 4233 29411 4267
rect 11897 4165 11931 4199
rect 17233 4165 17267 4199
rect 27353 4165 27387 4199
rect 2145 4097 2179 4131
rect 2421 4097 2455 4131
rect 2605 4097 2639 4131
rect 3433 4097 3467 4131
rect 3525 4097 3559 4131
rect 4261 4097 4295 4131
rect 4528 4097 4562 4131
rect 6837 4097 6871 4131
rect 8585 4097 8619 4131
rect 9413 4097 9447 4131
rect 9689 4097 9723 4131
rect 9873 4097 9907 4131
rect 10517 4097 10551 4131
rect 10793 4097 10827 4131
rect 14289 4097 14323 4131
rect 14565 4097 14599 4131
rect 14749 4097 14783 4131
rect 15117 4097 15151 4131
rect 15393 4097 15427 4131
rect 15669 4097 15703 4131
rect 15853 4097 15887 4131
rect 16964 4097 16998 4131
rect 17105 4097 17139 4131
rect 17325 4097 17359 4131
rect 17422 4097 17456 4131
rect 18337 4097 18371 4131
rect 18613 4097 18647 4131
rect 18797 4097 18831 4131
rect 19441 4097 19475 4131
rect 19901 4097 19935 4131
rect 20168 4097 20202 4131
rect 22017 4097 22051 4131
rect 22569 4097 22603 4131
rect 23857 4097 23891 4131
rect 25329 4097 25363 4131
rect 25605 4097 25639 4131
rect 25789 4097 25823 4131
rect 26433 4097 26467 4131
rect 26985 4097 27019 4131
rect 27078 4097 27112 4131
rect 27261 4097 27295 4131
rect 27450 4097 27484 4131
rect 28273 4097 28307 4131
rect 28549 4097 28583 4131
rect 28733 4097 28767 4131
rect 29561 4097 29595 4131
rect 29837 4097 29871 4131
rect 30481 4097 30515 4131
rect 30757 4097 30791 4131
rect 30941 4097 30975 4131
rect 3709 4029 3743 4063
rect 7021 4029 7055 4063
rect 7573 4029 7607 4063
rect 8769 4029 8803 4063
rect 22845 4029 22879 4063
rect 24133 4029 24167 4063
rect 30297 4029 30331 4063
rect 5641 3961 5675 3995
rect 7941 3961 7975 3995
rect 15209 3961 15243 3995
rect 26249 3961 26283 3995
rect 29745 3961 29779 3995
rect 6377 3893 6411 3927
rect 8033 3893 8067 3927
rect 9229 3893 9263 3927
rect 10701 3893 10735 3927
rect 13185 3893 13219 3927
rect 14105 3893 14139 3927
rect 19257 3893 19291 3927
rect 21833 3893 21867 3927
rect 25145 3893 25179 3927
rect 27629 3893 27663 3927
rect 28089 3893 28123 3927
rect 2329 3689 2363 3723
rect 5457 3689 5491 3723
rect 5825 3689 5859 3723
rect 7941 3689 7975 3723
rect 12909 3689 12943 3723
rect 17325 3689 17359 3723
rect 19257 3689 19291 3723
rect 19901 3689 19935 3723
rect 21005 3689 21039 3723
rect 23397 3689 23431 3723
rect 23765 3689 23799 3723
rect 26525 3689 26559 3723
rect 30665 3689 30699 3723
rect 3157 3621 3191 3655
rect 3525 3621 3559 3655
rect 13369 3621 13403 3655
rect 31033 3621 31067 3655
rect 1961 3553 1995 3587
rect 4169 3553 4203 3587
rect 5917 3553 5951 3587
rect 11529 3553 11563 3587
rect 15393 3553 15427 3587
rect 31125 3553 31159 3587
rect 2145 3485 2179 3519
rect 2973 3485 3007 3519
rect 3249 3485 3283 3519
rect 3525 3485 3559 3519
rect 4445 3485 4479 3519
rect 5641 3485 5675 3519
rect 6929 3485 6963 3519
rect 9229 3485 9263 3519
rect 9505 3485 9539 3519
rect 9689 3485 9723 3519
rect 10333 3485 10367 3519
rect 10609 3485 10643 3519
rect 10793 3485 10827 3519
rect 11796 3485 11830 3519
rect 13369 3485 13403 3519
rect 13553 3485 13587 3519
rect 14289 3485 14323 3519
rect 14565 3485 14599 3519
rect 14749 3485 14783 3519
rect 15669 3485 15703 3519
rect 16681 3485 16715 3519
rect 16774 3485 16808 3519
rect 16957 3485 16991 3519
rect 17146 3485 17180 3519
rect 18245 3485 18279 3519
rect 18521 3485 18555 3519
rect 18705 3485 18739 3519
rect 19441 3485 19475 3519
rect 20085 3485 20119 3519
rect 20361 3485 20395 3519
rect 20545 3485 20579 3519
rect 21189 3485 21223 3519
rect 21465 3485 21499 3519
rect 21649 3485 21683 3519
rect 22293 3485 22327 3519
rect 22569 3485 22603 3519
rect 22753 3485 22787 3519
rect 23581 3485 23615 3519
rect 23857 3485 23891 3519
rect 24961 3485 24995 3519
rect 25237 3485 25271 3519
rect 25421 3485 25455 3519
rect 25973 3485 26007 3519
rect 26157 3485 26191 3519
rect 26341 3485 26375 3519
rect 26985 3485 27019 3519
rect 29745 3485 29779 3519
rect 30021 3485 30055 3519
rect 30205 3485 30239 3519
rect 30849 3485 30883 3519
rect 6653 3417 6687 3451
rect 7021 3417 7055 3451
rect 7389 3417 7423 3451
rect 17049 3417 17083 3451
rect 26249 3417 26283 3451
rect 28733 3417 28767 3451
rect 2789 3349 2823 3383
rect 7757 3349 7791 3383
rect 9045 3349 9079 3383
rect 10149 3349 10183 3383
rect 14105 3349 14139 3383
rect 18061 3349 18095 3383
rect 22109 3349 22143 3383
rect 24777 3349 24811 3383
rect 29561 3349 29595 3383
rect 14197 3145 14231 3179
rect 15853 3145 15887 3179
rect 18889 3145 18923 3179
rect 20453 3145 20487 3179
rect 28733 3145 28767 3179
rect 30757 3145 30791 3179
rect 6009 3077 6043 3111
rect 6377 3077 6411 3111
rect 9137 3077 9171 3111
rect 11161 3077 11195 3111
rect 2145 3009 2179 3043
rect 2421 3009 2455 3043
rect 2605 3009 2639 3043
rect 3249 3009 3283 3043
rect 3525 3009 3559 3043
rect 3709 3009 3743 3043
rect 4445 3009 4479 3043
rect 4712 3009 4746 3043
rect 5825 2873 5859 2907
rect 6561 3009 6595 3043
rect 6837 3009 6871 3043
rect 7021 3009 7055 3043
rect 7389 3009 7423 3043
rect 7941 3009 7975 3043
rect 8953 3009 8987 3043
rect 9597 3009 9631 3043
rect 9864 3009 9898 3043
rect 8033 2941 8067 2975
rect 8217 2941 8251 2975
rect 8769 2941 8803 2975
rect 7389 2873 7423 2907
rect 7573 2873 7607 2907
rect 10977 2873 11011 2907
rect 1961 2805 1995 2839
rect 3065 2805 3099 2839
rect 6009 2805 6043 2839
rect 11713 3009 11747 3043
rect 12817 3009 12851 3043
rect 13084 3009 13118 3043
rect 14841 3009 14875 3043
rect 15117 3009 15151 3043
rect 15301 3009 15335 3043
rect 15761 3009 15795 3043
rect 15945 3009 15979 3043
rect 16865 3009 16899 3043
rect 17141 3009 17175 3043
rect 17325 3009 17359 3043
rect 18061 3009 18095 3043
rect 18337 3009 18371 3043
rect 18613 3009 18647 3043
rect 18797 3009 18831 3043
rect 18889 3009 18923 3043
rect 19717 3009 19751 3043
rect 20637 3009 20671 3043
rect 20913 3009 20947 3043
rect 21097 3009 21131 3043
rect 21189 3009 21223 3043
rect 22293 3009 22327 3043
rect 22569 3009 22603 3043
rect 22753 3009 22787 3043
rect 23213 3009 23247 3043
rect 23469 3009 23503 3043
rect 25513 3009 25547 3043
rect 25789 3009 25823 3043
rect 25973 3009 26007 3043
rect 27629 3009 27663 3043
rect 27905 3009 27939 3043
rect 28089 3009 28123 3043
rect 28917 3009 28951 3043
rect 29644 3009 29678 3043
rect 11529 2941 11563 2975
rect 11989 2941 12023 2975
rect 19993 2941 20027 2975
rect 18061 2873 18095 2907
rect 19901 2873 19935 2907
rect 29377 2941 29411 2975
rect 24593 2873 24627 2907
rect 11161 2805 11195 2839
rect 11897 2805 11931 2839
rect 14657 2805 14691 2839
rect 16681 2805 16715 2839
rect 18153 2805 18187 2839
rect 19533 2805 19567 2839
rect 21189 2805 21223 2839
rect 22109 2805 22143 2839
rect 25329 2805 25363 2839
rect 27445 2805 27479 2839
rect 2973 2601 3007 2635
rect 5181 2601 5215 2635
rect 6377 2601 6411 2635
rect 10977 2601 11011 2635
rect 12909 2601 12943 2635
rect 13369 2601 13403 2635
rect 20637 2601 20671 2635
rect 22753 2601 22787 2635
rect 24409 2601 24443 2635
rect 1593 2465 1627 2499
rect 3801 2465 3835 2499
rect 949 2397 983 2431
rect 5641 2397 5675 2431
rect 1860 2329 1894 2363
rect 4046 2329 4080 2363
rect 10333 2533 10367 2567
rect 7849 2465 7883 2499
rect 11529 2465 11563 2499
rect 14565 2465 14599 2499
rect 18705 2465 18739 2499
rect 24409 2465 24443 2499
rect 28917 2601 28951 2635
rect 30665 2601 30699 2635
rect 30297 2533 30331 2567
rect 31125 2465 31159 2499
rect 6653 2397 6687 2431
rect 6929 2397 6963 2431
rect 7113 2397 7147 2431
rect 7573 2397 7607 2431
rect 8953 2397 8987 2431
rect 10885 2397 10919 2431
rect 13553 2397 13587 2431
rect 16405 2397 16439 2431
rect 18429 2397 18463 2431
rect 18613 2397 18647 2431
rect 19257 2397 19291 2431
rect 21373 2397 21407 2431
rect 23397 2397 23431 2431
rect 23673 2397 23707 2431
rect 23857 2397 23891 2431
rect 24501 2397 24535 2431
rect 26341 2397 26375 2431
rect 28365 2397 28399 2431
rect 28641 2397 28675 2431
rect 28825 2397 28859 2431
rect 28917 2397 28951 2431
rect 29738 2397 29772 2431
rect 30021 2397 30055 2431
rect 30205 2397 30239 2431
rect 30297 2397 30331 2431
rect 30849 2397 30883 2431
rect 31033 2397 31067 2431
rect 9220 2329 9254 2363
rect 11796 2329 11830 2363
rect 14832 2329 14866 2363
rect 16672 2329 16706 2363
rect 18245 2329 18279 2363
rect 19502 2329 19536 2363
rect 21618 2329 21652 2363
rect 24768 2329 24802 2363
rect 26586 2329 26620 2363
rect 5825 2261 5859 2295
rect 6377 2261 6411 2295
rect 6469 2261 6503 2295
rect 15945 2261 15979 2295
rect 17785 2261 17819 2295
rect 23213 2261 23247 2295
rect 25881 2261 25915 2295
rect 27721 2261 27755 2295
rect 28181 2261 28215 2295
rect 29561 2261 29595 2295
rect 2145 2057 2179 2091
rect 3157 2057 3191 2091
rect 5825 2057 5859 2091
rect 8585 2057 8619 2091
rect 10977 2057 11011 2091
rect 21281 2057 21315 2091
rect 23305 2057 23339 2091
rect 25421 2057 25455 2091
rect 25973 2057 26007 2091
rect 31125 2057 31159 2091
rect 1501 1989 1535 2023
rect 4712 1989 4746 2023
rect 11774 1989 11808 2023
rect 13369 1989 13403 2023
rect 2329 1921 2363 1955
rect 2513 1921 2547 1955
rect 3341 1921 3375 1955
rect 3617 1921 3651 1955
rect 4445 1921 4479 1955
rect 6745 1921 6779 1955
rect 7205 1921 7239 1955
rect 7472 1921 7506 1955
rect 9597 1921 9631 1955
rect 9853 1921 9887 1955
rect 11529 1921 11563 1955
rect 13553 1921 13587 1955
rect 14565 1921 14599 1955
rect 14832 1921 14866 1955
rect 17049 1921 17083 1955
rect 17325 1921 17359 1955
rect 17509 1921 17543 1955
rect 18061 1921 18095 1955
rect 18328 1921 18362 1955
rect 19901 1921 19935 1955
rect 20157 1921 20191 1955
rect 21925 1921 21959 1955
rect 22192 1921 22226 1955
rect 24041 1921 24075 1955
rect 24308 1921 24342 1955
rect 26157 1921 26191 1955
rect 26341 1921 26375 1955
rect 26433 1921 26467 1955
rect 27445 1921 27479 1955
rect 27712 1921 27746 1955
rect 29285 1921 29319 1955
rect 29552 1921 29586 1955
rect 31309 1921 31343 1955
rect 2605 1853 2639 1887
rect 3525 1853 3559 1887
rect 13829 1853 13863 1887
rect 12909 1785 12943 1819
rect 28825 1785 28859 1819
rect 30665 1785 30699 1819
rect 1593 1717 1627 1751
rect 6561 1717 6595 1751
rect 13737 1717 13771 1751
rect 15945 1717 15979 1751
rect 16865 1717 16899 1751
rect 19441 1717 19475 1751
rect 1961 1513 1995 1547
rect 2697 1513 2731 1547
rect 6377 1513 6411 1547
rect 7297 1513 7331 1547
rect 10241 1513 10275 1547
rect 13093 1513 13127 1547
rect 13461 1513 13495 1547
rect 14381 1513 14415 1547
rect 14749 1513 14783 1547
rect 15669 1513 15703 1547
rect 16681 1513 16715 1547
rect 18245 1513 18279 1547
rect 18613 1513 18647 1547
rect 22477 1513 22511 1547
rect 24685 1513 24719 1547
rect 25789 1513 25823 1547
rect 26157 1513 26191 1547
rect 27905 1513 27939 1547
rect 28825 1513 28859 1547
rect 30665 1513 30699 1547
rect 4813 1445 4847 1479
rect 6837 1377 6871 1411
rect 11529 1377 11563 1411
rect 2513 1309 2547 1343
rect 3893 1309 3927 1343
rect 4629 1309 4663 1343
rect 5825 1309 5859 1343
rect 6561 1309 6595 1343
rect 6745 1309 6779 1343
rect 7481 1309 7515 1343
rect 7665 1309 7699 1343
rect 7757 1309 7791 1343
rect 8401 1309 8435 1343
rect 8953 1309 8987 1343
rect 9229 1309 9263 1343
rect 10425 1309 10459 1343
rect 10609 1309 10643 1343
rect 10701 1309 10735 1343
rect 11713 1309 11747 1343
rect 12541 1309 12575 1343
rect 13001 1309 13035 1343
rect 13277 1309 13311 1343
rect 13553 1309 13587 1343
rect 14289 1309 14323 1343
rect 1869 1241 1903 1275
rect 11897 1241 11931 1275
rect 27261 1445 27295 1479
rect 27537 1445 27571 1479
rect 15209 1377 15243 1411
rect 17141 1377 17175 1411
rect 20913 1377 20947 1411
rect 22845 1377 22879 1411
rect 23765 1377 23799 1411
rect 25145 1377 25179 1411
rect 26249 1377 26283 1411
rect 14933 1309 14967 1343
rect 15117 1309 15151 1343
rect 15301 1309 15335 1343
rect 15853 1309 15887 1343
rect 16037 1309 16071 1343
rect 16129 1309 16163 1343
rect 16865 1309 16899 1343
rect 17049 1309 17083 1343
rect 17233 1309 17267 1343
rect 17785 1309 17819 1343
rect 18429 1309 18463 1343
rect 18705 1309 18739 1343
rect 19625 1309 19659 1343
rect 20269 1309 20303 1343
rect 21097 1309 21131 1343
rect 21373 1309 21407 1343
rect 22017 1309 22051 1343
rect 22661 1309 22695 1343
rect 22937 1309 22971 1343
rect 23581 1309 23615 1343
rect 23857 1309 23891 1343
rect 24869 1309 24903 1343
rect 25053 1309 25087 1343
rect 25237 1309 25271 1343
rect 25973 1309 26007 1343
rect 27445 1309 27479 1343
rect 3985 1173 4019 1207
rect 5641 1173 5675 1207
rect 8217 1173 8251 1207
rect 12357 1173 12391 1207
rect 13001 1173 13035 1207
rect 14105 1173 14139 1207
rect 14381 1173 14415 1207
rect 15301 1173 15335 1207
rect 31033 1377 31067 1411
rect 28089 1309 28123 1343
rect 28273 1309 28307 1343
rect 28365 1309 28399 1343
rect 29009 1309 29043 1343
rect 29745 1309 29779 1343
rect 30849 1309 30883 1343
rect 31125 1309 31159 1343
rect 27537 1241 27571 1275
rect 17233 1173 17267 1207
rect 17601 1173 17635 1207
rect 19441 1173 19475 1207
rect 20085 1173 20119 1207
rect 21281 1173 21315 1207
rect 21373 1173 21407 1207
rect 21833 1173 21867 1207
rect 23397 1173 23431 1207
rect 25237 1173 25271 1207
rect 29561 1173 29595 1207
rect 17233 969 17267 1003
rect 17233 629 17267 663
<< metal1 >>
rect 0 42616 800 42630
rect 0 42588 888 42616
rect 0 42574 800 42588
rect 860 42480 888 42588
rect 25774 42576 25780 42628
rect 25832 42616 25838 42628
rect 29730 42616 29736 42628
rect 25832 42588 29736 42616
rect 25832 42576 25838 42588
rect 29730 42576 29736 42588
rect 29788 42576 29794 42628
rect 32320 42616 33120 42630
rect 32232 42588 33120 42616
rect 25590 42508 25596 42560
rect 25648 42548 25654 42560
rect 30098 42548 30104 42560
rect 25648 42520 30104 42548
rect 25648 42508 25654 42520
rect 30098 42508 30104 42520
rect 30156 42508 30162 42560
rect 32232 42480 32260 42588
rect 32320 42574 33120 42588
rect 768 42452 888 42480
rect 1104 42458 32016 42480
rect 768 42276 796 42452
rect 1104 42406 7288 42458
rect 7340 42406 17592 42458
rect 17644 42406 27896 42458
rect 27948 42406 32016 42458
rect 32232 42452 32352 42480
rect 1104 42384 32016 42406
rect 1210 42304 1216 42356
rect 1268 42344 1274 42356
rect 4341 42347 4399 42353
rect 4341 42344 4353 42347
rect 1268 42316 4353 42344
rect 1268 42304 1274 42316
rect 4341 42313 4353 42316
rect 4387 42313 4399 42347
rect 4341 42307 4399 42313
rect 7469 42347 7527 42353
rect 7469 42313 7481 42347
rect 7515 42344 7527 42347
rect 8202 42344 8208 42356
rect 7515 42316 8208 42344
rect 7515 42313 7527 42316
rect 7469 42307 7527 42313
rect 8202 42304 8208 42316
rect 8260 42304 8266 42356
rect 16209 42347 16267 42353
rect 16209 42313 16221 42347
rect 16255 42344 16267 42347
rect 20438 42344 20444 42356
rect 16255 42316 20444 42344
rect 16255 42313 16267 42316
rect 16209 42307 16267 42313
rect 20438 42304 20444 42316
rect 20496 42304 20502 42356
rect 21177 42347 21235 42353
rect 21177 42313 21189 42347
rect 21223 42313 21235 42347
rect 21177 42307 21235 42313
rect 22281 42347 22339 42353
rect 22281 42313 22293 42347
rect 22327 42344 22339 42347
rect 22327 42316 31754 42344
rect 22327 42313 22339 42316
rect 22281 42307 22339 42313
rect 4249 42279 4307 42285
rect 4249 42276 4261 42279
rect 768 42248 4261 42276
rect 4249 42245 4261 42248
rect 4295 42245 4307 42279
rect 21192 42276 21220 42307
rect 23661 42279 23719 42285
rect 23661 42276 23673 42279
rect 4249 42239 4307 42245
rect 15396 42248 21220 42276
rect 22066 42248 23673 42276
rect 1486 42168 1492 42220
rect 1544 42208 1550 42220
rect 1857 42211 1915 42217
rect 1857 42208 1869 42211
rect 1544 42180 1869 42208
rect 1544 42168 1550 42180
rect 1857 42177 1869 42180
rect 1903 42177 1915 42211
rect 2866 42208 2872 42220
rect 2827 42180 2872 42208
rect 1857 42171 1915 42177
rect 2866 42168 2872 42180
rect 2924 42168 2930 42220
rect 7650 42208 7656 42220
rect 7611 42180 7656 42208
rect 7650 42168 7656 42180
rect 7708 42168 7714 42220
rect 8110 42168 8116 42220
rect 8168 42208 8174 42220
rect 8205 42211 8263 42217
rect 8205 42208 8217 42211
rect 8168 42180 8217 42208
rect 8168 42168 8174 42180
rect 8205 42177 8217 42180
rect 8251 42177 8263 42211
rect 9122 42208 9128 42220
rect 9083 42180 9128 42208
rect 8205 42171 8263 42177
rect 9122 42168 9128 42180
rect 9180 42168 9186 42220
rect 10045 42211 10103 42217
rect 10045 42177 10057 42211
rect 10091 42208 10103 42211
rect 10226 42208 10232 42220
rect 10091 42180 10232 42208
rect 10091 42177 10103 42180
rect 10045 42171 10103 42177
rect 10226 42168 10232 42180
rect 10284 42168 10290 42220
rect 12710 42208 12716 42220
rect 12671 42180 12716 42208
rect 12710 42168 12716 42180
rect 12768 42168 12774 42220
rect 15396 42217 15424 42248
rect 15381 42211 15439 42217
rect 15381 42177 15393 42211
rect 15427 42177 15439 42211
rect 15381 42171 15439 42177
rect 15933 42211 15991 42217
rect 15933 42177 15945 42211
rect 15979 42208 15991 42211
rect 16209 42211 16267 42217
rect 16209 42208 16221 42211
rect 15979 42180 16221 42208
rect 15979 42177 15991 42180
rect 15933 42171 15991 42177
rect 16209 42177 16221 42180
rect 16255 42177 16267 42211
rect 16209 42171 16267 42177
rect 16853 42211 16911 42217
rect 16853 42177 16865 42211
rect 16899 42177 16911 42211
rect 18138 42208 18144 42220
rect 18099 42180 18144 42208
rect 16853 42171 16911 42177
rect 3145 42143 3203 42149
rect 3145 42109 3157 42143
rect 3191 42140 3203 42143
rect 3234 42140 3240 42152
rect 3191 42112 3240 42140
rect 3191 42109 3203 42112
rect 3145 42103 3203 42109
rect 3234 42100 3240 42112
rect 3292 42100 3298 42152
rect 8386 42100 8392 42152
rect 8444 42140 8450 42152
rect 9401 42143 9459 42149
rect 9401 42140 9413 42143
rect 8444 42112 9413 42140
rect 8444 42100 8450 42112
rect 9401 42109 9413 42112
rect 9447 42109 9459 42143
rect 12986 42140 12992 42152
rect 12947 42112 12992 42140
rect 9401 42103 9459 42109
rect 12986 42100 12992 42112
rect 13044 42100 13050 42152
rect 16390 42100 16396 42152
rect 16448 42140 16454 42152
rect 16868 42140 16896 42171
rect 18138 42168 18144 42180
rect 18196 42168 18202 42220
rect 19886 42168 19892 42220
rect 19944 42208 19950 42220
rect 20053 42211 20111 42217
rect 20053 42208 20065 42211
rect 19944 42180 20065 42208
rect 19944 42168 19950 42180
rect 20053 42177 20065 42180
rect 20099 42177 20111 42211
rect 20053 42171 20111 42177
rect 20438 42168 20444 42220
rect 20496 42208 20502 42220
rect 22066 42208 22094 42248
rect 23661 42245 23673 42248
rect 23707 42245 23719 42279
rect 28997 42279 29055 42285
rect 28997 42276 29009 42279
rect 23661 42239 23719 42245
rect 24504 42248 29009 42276
rect 20496 42180 22094 42208
rect 22465 42211 22523 42217
rect 20496 42168 20502 42180
rect 22465 42177 22477 42211
rect 22511 42177 22523 42211
rect 22465 42171 22523 42177
rect 23109 42211 23167 42217
rect 23109 42177 23121 42211
rect 23155 42208 23167 42211
rect 24504 42208 24532 42248
rect 28997 42245 29009 42248
rect 29043 42245 29055 42279
rect 28997 42239 29055 42245
rect 23155 42180 24532 42208
rect 24581 42211 24639 42217
rect 23155 42177 23167 42180
rect 23109 42171 23167 42177
rect 24581 42177 24593 42211
rect 24627 42177 24639 42211
rect 24581 42171 24639 42177
rect 16448 42112 16896 42140
rect 17129 42143 17187 42149
rect 16448 42100 16454 42112
rect 17129 42109 17141 42143
rect 17175 42140 17187 42143
rect 17218 42140 17224 42152
rect 17175 42112 17224 42140
rect 17175 42109 17187 42112
rect 17129 42103 17187 42109
rect 17218 42100 17224 42112
rect 17276 42100 17282 42152
rect 18046 42100 18052 42152
rect 18104 42140 18110 42152
rect 18417 42143 18475 42149
rect 18417 42140 18429 42143
rect 18104 42112 18429 42140
rect 18104 42100 18110 42112
rect 18417 42109 18429 42112
rect 18463 42109 18475 42143
rect 18417 42103 18475 42109
rect 19334 42100 19340 42152
rect 19392 42140 19398 42152
rect 19797 42143 19855 42149
rect 19797 42140 19809 42143
rect 19392 42112 19809 42140
rect 19392 42100 19398 42112
rect 19797 42109 19809 42112
rect 19843 42109 19855 42143
rect 22480 42140 22508 42171
rect 24596 42140 24624 42171
rect 25406 42168 25412 42220
rect 25464 42208 25470 42220
rect 25774 42208 25780 42220
rect 25464 42180 25780 42208
rect 25464 42168 25470 42180
rect 25774 42168 25780 42180
rect 25832 42168 25838 42220
rect 26421 42211 26479 42217
rect 26421 42177 26433 42211
rect 26467 42177 26479 42211
rect 27154 42208 27160 42220
rect 27115 42180 27160 42208
rect 26421 42171 26479 42177
rect 26436 42140 26464 42171
rect 27154 42168 27160 42180
rect 27212 42168 27218 42220
rect 28626 42208 28632 42220
rect 27255 42180 27568 42208
rect 28587 42180 28632 42208
rect 26602 42140 26608 42152
rect 22480 42112 24532 42140
rect 24596 42112 26608 42140
rect 19797 42103 19855 42109
rect 2590 42032 2596 42084
rect 2648 42072 2654 42084
rect 3053 42075 3111 42081
rect 3053 42072 3065 42075
rect 2648 42044 3065 42072
rect 2648 42032 2654 42044
rect 3053 42041 3065 42044
rect 3099 42041 3111 42075
rect 3053 42035 3111 42041
rect 9030 42032 9036 42084
rect 9088 42072 9094 42084
rect 9861 42075 9919 42081
rect 9861 42072 9873 42075
rect 9088 42044 9873 42072
rect 9088 42032 9094 42044
rect 9861 42041 9873 42044
rect 9907 42041 9919 42075
rect 9861 42035 9919 42041
rect 16022 42032 16028 42084
rect 16080 42072 16086 42084
rect 16117 42075 16175 42081
rect 16117 42072 16129 42075
rect 16080 42044 16129 42072
rect 16080 42032 16086 42044
rect 16117 42041 16129 42044
rect 16163 42072 16175 42075
rect 17037 42075 17095 42081
rect 17037 42072 17049 42075
rect 16163 42044 17049 42072
rect 16163 42041 16175 42044
rect 16117 42035 16175 42041
rect 17037 42041 17049 42044
rect 17083 42041 17095 42075
rect 17037 42035 17095 42041
rect 17957 42075 18015 42081
rect 17957 42041 17969 42075
rect 18003 42072 18015 42075
rect 18598 42072 18604 42084
rect 18003 42044 18604 42072
rect 18003 42041 18015 42044
rect 17957 42035 18015 42041
rect 18598 42032 18604 42044
rect 18656 42032 18662 42084
rect 23014 42032 23020 42084
rect 23072 42072 23078 42084
rect 24397 42075 24455 42081
rect 24397 42072 24409 42075
rect 23072 42044 24409 42072
rect 23072 42032 23078 42044
rect 24397 42041 24409 42044
rect 24443 42041 24455 42075
rect 24504 42072 24532 42112
rect 26602 42100 26608 42112
rect 26660 42100 26666 42152
rect 27255 42072 27283 42180
rect 27338 42100 27344 42152
rect 27396 42140 27402 42152
rect 27433 42143 27491 42149
rect 27433 42140 27445 42143
rect 27396 42112 27445 42140
rect 27396 42100 27402 42112
rect 27433 42109 27445 42112
rect 27479 42109 27491 42143
rect 27540 42140 27568 42180
rect 28626 42168 28632 42180
rect 28684 42168 28690 42220
rect 29730 42208 29736 42220
rect 28736 42180 29112 42208
rect 29691 42180 29736 42208
rect 28736 42140 28764 42180
rect 27540 42112 28764 42140
rect 27433 42103 27491 42109
rect 28810 42100 28816 42152
rect 28868 42140 28874 42152
rect 28905 42143 28963 42149
rect 28905 42140 28917 42143
rect 28868 42112 28917 42140
rect 28868 42100 28874 42112
rect 28905 42109 28917 42112
rect 28951 42109 28963 42143
rect 29084 42140 29112 42180
rect 29730 42168 29736 42180
rect 29788 42168 29794 42220
rect 30377 42211 30435 42217
rect 30377 42177 30389 42211
rect 30423 42177 30435 42211
rect 30377 42171 30435 42177
rect 31297 42211 31355 42217
rect 31297 42177 31309 42211
rect 31343 42208 31355 42211
rect 31386 42208 31392 42220
rect 31343 42180 31392 42208
rect 31343 42177 31355 42180
rect 31297 42171 31355 42177
rect 30392 42140 30420 42171
rect 31386 42168 31392 42180
rect 31444 42168 31450 42220
rect 31478 42140 31484 42152
rect 29084 42112 30328 42140
rect 30392 42112 31484 42140
rect 28905 42103 28963 42109
rect 27614 42072 27620 42084
rect 24504 42044 27283 42072
rect 27356 42044 27620 42072
rect 24397 42035 24455 42041
rect 1578 41964 1584 42016
rect 1636 42004 1642 42016
rect 1949 42007 2007 42013
rect 1949 42004 1961 42007
rect 1636 41976 1961 42004
rect 1636 41964 1642 41976
rect 1949 41973 1961 41976
rect 1995 41973 2007 42007
rect 2682 42004 2688 42016
rect 2643 41976 2688 42004
rect 1949 41967 2007 41973
rect 2682 41964 2688 41976
rect 2740 41964 2746 42016
rect 8297 42007 8355 42013
rect 8297 41973 8309 42007
rect 8343 42004 8355 42007
rect 8570 42004 8576 42016
rect 8343 41976 8576 42004
rect 8343 41973 8355 41976
rect 8297 41967 8355 41973
rect 8570 41964 8576 41976
rect 8628 41964 8634 42016
rect 8938 42004 8944 42016
rect 8899 41976 8944 42004
rect 8938 41964 8944 41976
rect 8996 41964 9002 42016
rect 9309 42007 9367 42013
rect 9309 41973 9321 42007
rect 9355 42004 9367 42007
rect 10778 42004 10784 42016
rect 9355 41976 10784 42004
rect 9355 41973 9367 41976
rect 9309 41967 9367 41973
rect 10778 41964 10784 41976
rect 10836 41964 10842 42016
rect 12342 41964 12348 42016
rect 12400 42004 12406 42016
rect 12529 42007 12587 42013
rect 12529 42004 12541 42007
rect 12400 41976 12541 42004
rect 12400 41964 12406 41976
rect 12529 41973 12541 41976
rect 12575 41973 12587 42007
rect 12894 42004 12900 42016
rect 12855 41976 12900 42004
rect 12529 41967 12587 41973
rect 12894 41964 12900 41976
rect 12952 41964 12958 42016
rect 15197 42007 15255 42013
rect 15197 41973 15209 42007
rect 15243 42004 15255 42007
rect 16206 42004 16212 42016
rect 15243 41976 16212 42004
rect 15243 41973 15255 41976
rect 15197 41967 15255 41973
rect 16206 41964 16212 41976
rect 16264 41964 16270 42016
rect 16666 42004 16672 42016
rect 16627 41976 16672 42004
rect 16666 41964 16672 41976
rect 16724 41964 16730 42016
rect 18325 42007 18383 42013
rect 18325 41973 18337 42007
rect 18371 42004 18383 42007
rect 19058 42004 19064 42016
rect 18371 41976 19064 42004
rect 18371 41973 18383 41976
rect 18325 41967 18383 41973
rect 19058 41964 19064 41976
rect 19116 41964 19122 42016
rect 22925 42007 22983 42013
rect 22925 41973 22937 42007
rect 22971 42004 22983 42007
rect 23566 42004 23572 42016
rect 22971 41976 23572 42004
rect 22971 41973 22983 41976
rect 22925 41967 22983 41973
rect 23566 41964 23572 41976
rect 23624 41964 23630 42016
rect 23658 41964 23664 42016
rect 23716 42004 23722 42016
rect 23753 42007 23811 42013
rect 23753 42004 23765 42007
rect 23716 41976 23765 42004
rect 23716 41964 23722 41976
rect 23753 41973 23765 41976
rect 23799 41973 23811 42007
rect 25590 42004 25596 42016
rect 25551 41976 25596 42004
rect 23753 41967 23811 41973
rect 25590 41964 25596 41976
rect 25648 41964 25654 42016
rect 26234 42004 26240 42016
rect 26195 41976 26240 42004
rect 26234 41964 26240 41976
rect 26292 41964 26298 42016
rect 26973 42007 27031 42013
rect 26973 41973 26985 42007
rect 27019 42004 27031 42007
rect 27246 42004 27252 42016
rect 27019 41976 27252 42004
rect 27019 41973 27031 41976
rect 26973 41967 27031 41973
rect 27246 41964 27252 41976
rect 27304 41964 27310 42016
rect 27356 42013 27384 42044
rect 27614 42032 27620 42044
rect 27672 42072 27678 42084
rect 28534 42072 28540 42084
rect 27672 42044 28540 42072
rect 27672 42032 27678 42044
rect 28534 42032 28540 42044
rect 28592 42072 28598 42084
rect 28592 42044 28856 42072
rect 28592 42032 28598 42044
rect 27341 42007 27399 42013
rect 27341 41973 27353 42007
rect 27387 41973 27399 42007
rect 28442 42004 28448 42016
rect 28403 41976 28448 42004
rect 27341 41967 27399 41973
rect 28442 41964 28448 41976
rect 28500 41964 28506 42016
rect 28828 42013 28856 42044
rect 29362 42032 29368 42084
rect 29420 42072 29426 42084
rect 30193 42075 30251 42081
rect 30193 42072 30205 42075
rect 29420 42044 30205 42072
rect 29420 42032 29426 42044
rect 30193 42041 30205 42044
rect 30239 42041 30251 42075
rect 30300 42072 30328 42112
rect 31478 42100 31484 42112
rect 31536 42100 31542 42152
rect 31113 42075 31171 42081
rect 31113 42072 31125 42075
rect 30300 42044 31125 42072
rect 30193 42035 30251 42041
rect 31113 42041 31125 42044
rect 31159 42041 31171 42075
rect 31726 42072 31754 42316
rect 32324 42072 32352 42452
rect 31726 42044 32352 42072
rect 31113 42035 31171 42041
rect 28813 42007 28871 42013
rect 28813 41973 28825 42007
rect 28859 41973 28871 42007
rect 28813 41967 28871 41973
rect 28997 42007 29055 42013
rect 28997 41973 29009 42007
rect 29043 42004 29055 42007
rect 29549 42007 29607 42013
rect 29549 42004 29561 42007
rect 29043 41976 29561 42004
rect 29043 41973 29055 41976
rect 28997 41967 29055 41973
rect 29549 41973 29561 41976
rect 29595 41973 29607 42007
rect 29549 41967 29607 41973
rect 1104 41914 32016 41936
rect 1104 41862 2136 41914
rect 2188 41862 12440 41914
rect 12492 41862 22744 41914
rect 22796 41862 32016 41914
rect 1104 41840 32016 41862
rect 6181 41803 6239 41809
rect 6181 41769 6193 41803
rect 6227 41800 6239 41803
rect 8386 41800 8392 41812
rect 6227 41772 8248 41800
rect 8347 41772 8392 41800
rect 6227 41769 6239 41772
rect 6181 41763 6239 41769
rect 3237 41735 3295 41741
rect 3237 41701 3249 41735
rect 3283 41732 3295 41735
rect 8220 41732 8248 41772
rect 8386 41760 8392 41772
rect 8444 41760 8450 41812
rect 19058 41760 19064 41812
rect 19116 41800 19122 41812
rect 19613 41803 19671 41809
rect 19613 41800 19625 41803
rect 19116 41772 19625 41800
rect 19116 41760 19122 41772
rect 19613 41769 19625 41772
rect 19659 41769 19671 41803
rect 19613 41763 19671 41769
rect 26605 41803 26663 41809
rect 26605 41769 26617 41803
rect 26651 41800 26663 41803
rect 27614 41800 27620 41812
rect 26651 41772 27620 41800
rect 26651 41769 26663 41772
rect 26605 41763 26663 41769
rect 27614 41760 27620 41772
rect 27672 41760 27678 41812
rect 8570 41732 8576 41744
rect 3283 41704 4292 41732
rect 8220 41704 8576 41732
rect 3283 41701 3295 41704
rect 3237 41695 3295 41701
rect 1394 41556 1400 41608
rect 1452 41596 1458 41608
rect 1857 41599 1915 41605
rect 1857 41596 1869 41599
rect 1452 41568 1869 41596
rect 1452 41556 1458 41568
rect 1857 41565 1869 41568
rect 1903 41565 1915 41599
rect 1857 41559 1915 41565
rect 2124 41599 2182 41605
rect 2124 41565 2136 41599
rect 2170 41596 2182 41599
rect 2682 41596 2688 41608
rect 2170 41568 2688 41596
rect 2170 41565 2182 41568
rect 2124 41559 2182 41565
rect 2682 41556 2688 41568
rect 2740 41556 2746 41608
rect 3970 41596 3976 41608
rect 3931 41568 3976 41596
rect 3970 41556 3976 41568
rect 4028 41556 4034 41608
rect 4264 41605 4292 41704
rect 8570 41692 8576 41704
rect 8628 41732 8634 41744
rect 9309 41735 9367 41741
rect 9309 41732 9321 41735
rect 8628 41704 9321 41732
rect 8628 41692 8634 41704
rect 9309 41701 9321 41704
rect 9355 41701 9367 41735
rect 9309 41695 9367 41701
rect 18785 41735 18843 41741
rect 18785 41701 18797 41735
rect 18831 41732 18843 41735
rect 19426 41732 19432 41744
rect 18831 41704 19432 41732
rect 18831 41701 18843 41704
rect 18785 41695 18843 41701
rect 19426 41692 19432 41704
rect 19484 41692 19490 41744
rect 25777 41735 25835 41741
rect 25777 41701 25789 41735
rect 25823 41701 25835 41735
rect 25777 41695 25835 41701
rect 28997 41735 29055 41741
rect 28997 41701 29009 41735
rect 29043 41732 29055 41735
rect 29043 41704 29868 41732
rect 29043 41701 29055 41704
rect 28997 41695 29055 41701
rect 5258 41624 5264 41676
rect 5316 41664 5322 41676
rect 6273 41667 6331 41673
rect 6273 41664 6285 41667
rect 5316 41636 6285 41664
rect 5316 41624 5322 41636
rect 6273 41633 6285 41636
rect 6319 41633 6331 41667
rect 6273 41627 6331 41633
rect 8754 41624 8760 41676
rect 8812 41664 8818 41676
rect 9401 41667 9459 41673
rect 9401 41664 9413 41667
rect 8812 41636 9413 41664
rect 8812 41624 8818 41636
rect 9401 41633 9413 41636
rect 9447 41633 9459 41667
rect 9401 41627 9459 41633
rect 18049 41667 18107 41673
rect 18049 41633 18061 41667
rect 18095 41664 18107 41667
rect 18095 41636 19472 41664
rect 18095 41633 18107 41636
rect 18049 41627 18107 41633
rect 4157 41599 4215 41605
rect 4157 41565 4169 41599
rect 4203 41565 4215 41599
rect 4157 41559 4215 41565
rect 4249 41599 4307 41605
rect 4249 41565 4261 41599
rect 4295 41596 4307 41599
rect 4338 41596 4344 41608
rect 4295 41568 4344 41596
rect 4295 41565 4307 41568
rect 4249 41559 4307 41565
rect 4172 41528 4200 41559
rect 4338 41556 4344 41568
rect 4396 41556 4402 41608
rect 4893 41599 4951 41605
rect 4893 41596 4905 41599
rect 4448 41568 4905 41596
rect 2700 41500 4200 41528
rect 2700 41472 2728 41500
rect 2682 41420 2688 41472
rect 2740 41420 2746 41472
rect 3789 41463 3847 41469
rect 3789 41429 3801 41463
rect 3835 41460 3847 41463
rect 3878 41460 3884 41472
rect 3835 41432 3884 41460
rect 3835 41429 3847 41432
rect 3789 41423 3847 41429
rect 3878 41420 3884 41432
rect 3936 41420 3942 41472
rect 4062 41420 4068 41472
rect 4120 41460 4126 41472
rect 4448 41460 4476 41568
rect 4893 41565 4905 41568
rect 4939 41565 4951 41599
rect 4893 41559 4951 41565
rect 4982 41556 4988 41608
rect 5040 41596 5046 41608
rect 5169 41599 5227 41605
rect 5169 41596 5181 41599
rect 5040 41568 5181 41596
rect 5040 41556 5046 41568
rect 5169 41565 5181 41568
rect 5215 41565 5227 41599
rect 5350 41596 5356 41608
rect 5311 41568 5356 41596
rect 5169 41559 5227 41565
rect 5350 41556 5356 41568
rect 5408 41556 5414 41608
rect 5997 41599 6055 41605
rect 5997 41565 6009 41599
rect 6043 41565 6055 41599
rect 7006 41596 7012 41608
rect 6967 41568 7012 41596
rect 5997 41559 6055 41565
rect 4709 41531 4767 41537
rect 4709 41497 4721 41531
rect 4755 41528 4767 41531
rect 6012 41528 6040 41559
rect 7006 41556 7012 41568
rect 7064 41556 7070 41608
rect 8386 41556 8392 41608
rect 8444 41596 8450 41608
rect 9125 41599 9183 41605
rect 9125 41596 9137 41599
rect 8444 41568 9137 41596
rect 8444 41556 8450 41568
rect 9125 41565 9137 41568
rect 9171 41565 9183 41599
rect 9125 41559 9183 41565
rect 10045 41599 10103 41605
rect 10045 41565 10057 41599
rect 10091 41596 10103 41599
rect 11882 41596 11888 41608
rect 10091 41568 11888 41596
rect 10091 41565 10103 41568
rect 10045 41559 10103 41565
rect 11882 41556 11888 41568
rect 11940 41596 11946 41608
rect 12342 41605 12348 41608
rect 12069 41599 12127 41605
rect 12069 41596 12081 41599
rect 11940 41568 12081 41596
rect 11940 41556 11946 41568
rect 12069 41565 12081 41568
rect 12115 41565 12127 41599
rect 12336 41596 12348 41605
rect 12303 41568 12348 41596
rect 12069 41559 12127 41565
rect 12336 41559 12348 41568
rect 12342 41556 12348 41559
rect 12400 41556 12406 41608
rect 13998 41556 14004 41608
rect 14056 41596 14062 41608
rect 14093 41599 14151 41605
rect 14093 41596 14105 41599
rect 14056 41568 14105 41596
rect 14056 41556 14062 41568
rect 14093 41565 14105 41568
rect 14139 41596 14151 41599
rect 15933 41599 15991 41605
rect 15933 41596 15945 41599
rect 14139 41568 15945 41596
rect 14139 41565 14151 41568
rect 14093 41559 14151 41565
rect 15933 41565 15945 41568
rect 15979 41565 15991 41599
rect 15933 41559 15991 41565
rect 16200 41599 16258 41605
rect 16200 41565 16212 41599
rect 16246 41596 16258 41599
rect 16666 41596 16672 41608
rect 16246 41568 16672 41596
rect 16246 41565 16258 41568
rect 16200 41559 16258 41565
rect 16666 41556 16672 41568
rect 16724 41556 16730 41608
rect 18230 41596 18236 41608
rect 18191 41568 18236 41596
rect 18230 41556 18236 41568
rect 18288 41556 18294 41608
rect 18506 41596 18512 41608
rect 18467 41568 18512 41596
rect 18506 41556 18512 41568
rect 18564 41556 18570 41608
rect 19444 41605 19472 41636
rect 19518 41624 19524 41676
rect 19576 41664 19582 41676
rect 19705 41667 19763 41673
rect 19705 41664 19717 41667
rect 19576 41636 19717 41664
rect 19576 41624 19582 41636
rect 19705 41633 19717 41636
rect 19751 41633 19763 41667
rect 19705 41627 19763 41633
rect 23566 41624 23572 41676
rect 23624 41664 23630 41676
rect 23624 41636 24532 41664
rect 23624 41624 23630 41636
rect 18693 41599 18751 41605
rect 18693 41565 18705 41599
rect 18739 41596 18751 41599
rect 18785 41599 18843 41605
rect 18785 41596 18797 41599
rect 18739 41568 18797 41596
rect 18739 41565 18751 41568
rect 18693 41559 18751 41565
rect 18785 41565 18797 41568
rect 18831 41565 18843 41599
rect 18785 41559 18843 41565
rect 19429 41599 19487 41605
rect 19429 41565 19441 41599
rect 19475 41565 19487 41599
rect 19429 41559 19487 41565
rect 20625 41599 20683 41605
rect 20625 41565 20637 41599
rect 20671 41596 20683 41599
rect 21634 41596 21640 41608
rect 20671 41568 21640 41596
rect 20671 41565 20683 41568
rect 20625 41559 20683 41565
rect 10318 41537 10324 41540
rect 4755 41500 6040 41528
rect 7276 41531 7334 41537
rect 4755 41497 4767 41500
rect 4709 41491 4767 41497
rect 7276 41497 7288 41531
rect 7322 41528 7334 41531
rect 8941 41531 8999 41537
rect 8941 41528 8953 41531
rect 7322 41500 8953 41528
rect 7322 41497 7334 41500
rect 7276 41491 7334 41497
rect 8941 41497 8953 41500
rect 8987 41497 8999 41531
rect 8941 41491 8999 41497
rect 10312 41491 10324 41537
rect 10376 41528 10382 41540
rect 14360 41531 14418 41537
rect 10376 41500 10412 41528
rect 10318 41488 10324 41491
rect 10376 41488 10382 41500
rect 14360 41497 14372 41531
rect 14406 41528 14418 41531
rect 15102 41528 15108 41540
rect 14406 41500 15108 41528
rect 14406 41497 14418 41500
rect 14360 41491 14418 41497
rect 15102 41488 15108 41500
rect 15160 41488 15166 41540
rect 19334 41488 19340 41540
rect 19392 41528 19398 41540
rect 20640 41528 20668 41559
rect 21634 41556 21640 41568
rect 21692 41596 21698 41608
rect 22465 41599 22523 41605
rect 22465 41596 22477 41599
rect 21692 41568 22477 41596
rect 21692 41556 21698 41568
rect 22465 41565 22477 41568
rect 22511 41565 22523 41599
rect 24394 41596 24400 41608
rect 24355 41568 24400 41596
rect 22465 41559 22523 41565
rect 24394 41556 24400 41568
rect 24452 41556 24458 41608
rect 24504 41596 24532 41636
rect 25590 41624 25596 41676
rect 25648 41664 25654 41676
rect 25792 41664 25820 41695
rect 26697 41667 26755 41673
rect 26697 41664 26709 41667
rect 25648 41636 26709 41664
rect 25648 41624 25654 41636
rect 26697 41633 26709 41636
rect 26743 41633 26755 41667
rect 26697 41627 26755 41633
rect 29840 41608 29868 41704
rect 29917 41667 29975 41673
rect 29917 41633 29929 41667
rect 29963 41664 29975 41667
rect 31018 41664 31024 41676
rect 29963 41636 31024 41664
rect 29963 41633 29975 41636
rect 29917 41627 29975 41633
rect 31018 41624 31024 41636
rect 31076 41624 31082 41676
rect 26418 41596 26424 41608
rect 24504 41568 26280 41596
rect 26379 41568 26424 41596
rect 19392 41500 20668 41528
rect 20892 41531 20950 41537
rect 19392 41488 19398 41500
rect 20892 41497 20904 41531
rect 20938 41528 20950 41531
rect 21818 41528 21824 41540
rect 20938 41500 21824 41528
rect 20938 41497 20950 41500
rect 20892 41491 20950 41497
rect 21818 41488 21824 41500
rect 21876 41488 21882 41540
rect 22732 41531 22790 41537
rect 22732 41497 22744 41531
rect 22778 41528 22790 41531
rect 23290 41528 23296 41540
rect 22778 41500 23296 41528
rect 22778 41497 22790 41500
rect 22732 41491 22790 41497
rect 23290 41488 23296 41500
rect 23348 41488 23354 41540
rect 24664 41531 24722 41537
rect 24664 41497 24676 41531
rect 24710 41528 24722 41531
rect 24762 41528 24768 41540
rect 24710 41500 24768 41528
rect 24710 41497 24722 41500
rect 24664 41491 24722 41497
rect 24762 41488 24768 41500
rect 24820 41488 24826 41540
rect 26252 41528 26280 41568
rect 26418 41556 26424 41568
rect 26476 41556 26482 41608
rect 27614 41596 27620 41608
rect 27575 41568 27620 41596
rect 27614 41556 27620 41568
rect 27672 41556 27678 41608
rect 27884 41599 27942 41605
rect 27884 41565 27896 41599
rect 27930 41596 27942 41599
rect 28442 41596 28448 41608
rect 27930 41568 28448 41596
rect 27930 41565 27942 41568
rect 27884 41559 27942 41565
rect 28442 41556 28448 41568
rect 28500 41556 28506 41608
rect 29730 41596 29736 41608
rect 29691 41568 29736 41596
rect 29730 41556 29736 41568
rect 29788 41556 29794 41608
rect 29822 41556 29828 41608
rect 29880 41596 29886 41608
rect 30009 41599 30067 41605
rect 30009 41596 30021 41599
rect 29880 41568 30021 41596
rect 29880 41556 29886 41568
rect 30009 41565 30021 41568
rect 30055 41565 30067 41599
rect 30009 41559 30067 41565
rect 30653 41599 30711 41605
rect 30653 41565 30665 41599
rect 30699 41565 30711 41599
rect 31294 41596 31300 41608
rect 31255 41568 31300 41596
rect 30653 41559 30711 41565
rect 28350 41528 28356 41540
rect 26252 41500 28356 41528
rect 28350 41488 28356 41500
rect 28408 41488 28414 41540
rect 30668 41528 30696 41559
rect 31294 41556 31300 41568
rect 31352 41556 31358 41608
rect 31386 41528 31392 41540
rect 30668 41500 31392 41528
rect 31386 41488 31392 41500
rect 31444 41488 31450 41540
rect 5810 41460 5816 41472
rect 4120 41432 4476 41460
rect 5771 41432 5816 41460
rect 4120 41420 4126 41432
rect 5810 41420 5816 41432
rect 5868 41420 5874 41472
rect 11425 41463 11483 41469
rect 11425 41429 11437 41463
rect 11471 41460 11483 41463
rect 12250 41460 12256 41472
rect 11471 41432 12256 41460
rect 11471 41429 11483 41432
rect 11425 41423 11483 41429
rect 12250 41420 12256 41432
rect 12308 41420 12314 41472
rect 13449 41463 13507 41469
rect 13449 41429 13461 41463
rect 13495 41460 13507 41463
rect 14274 41460 14280 41472
rect 13495 41432 14280 41460
rect 13495 41429 13507 41432
rect 13449 41423 13507 41429
rect 14274 41420 14280 41432
rect 14332 41420 14338 41472
rect 15473 41463 15531 41469
rect 15473 41429 15485 41463
rect 15519 41460 15531 41463
rect 15746 41460 15752 41472
rect 15519 41432 15752 41460
rect 15519 41429 15531 41432
rect 15473 41423 15531 41429
rect 15746 41420 15752 41432
rect 15804 41420 15810 41472
rect 17310 41460 17316 41472
rect 17271 41432 17316 41460
rect 17310 41420 17316 41432
rect 17368 41420 17374 41472
rect 19150 41420 19156 41472
rect 19208 41460 19214 41472
rect 19245 41463 19303 41469
rect 19245 41460 19257 41463
rect 19208 41432 19257 41460
rect 19208 41420 19214 41432
rect 19245 41429 19257 41432
rect 19291 41429 19303 41463
rect 19245 41423 19303 41429
rect 22005 41463 22063 41469
rect 22005 41429 22017 41463
rect 22051 41460 22063 41463
rect 23566 41460 23572 41472
rect 22051 41432 23572 41460
rect 22051 41429 22063 41432
rect 22005 41423 22063 41429
rect 23566 41420 23572 41432
rect 23624 41420 23630 41472
rect 23842 41460 23848 41472
rect 23803 41432 23848 41460
rect 23842 41420 23848 41432
rect 23900 41420 23906 41472
rect 26050 41420 26056 41472
rect 26108 41460 26114 41472
rect 26237 41463 26295 41469
rect 26237 41460 26249 41463
rect 26108 41432 26249 41460
rect 26108 41420 26114 41432
rect 26237 41429 26249 41432
rect 26283 41429 26295 41463
rect 26237 41423 26295 41429
rect 29549 41463 29607 41469
rect 29549 41429 29561 41463
rect 29595 41460 29607 41463
rect 29638 41460 29644 41472
rect 29595 41432 29644 41460
rect 29595 41429 29607 41432
rect 29549 41423 29607 41429
rect 29638 41420 29644 41432
rect 29696 41420 29702 41472
rect 30282 41420 30288 41472
rect 30340 41460 30346 41472
rect 30469 41463 30527 41469
rect 30469 41460 30481 41463
rect 30340 41432 30481 41460
rect 30340 41420 30346 41432
rect 30469 41429 30481 41432
rect 30515 41429 30527 41463
rect 31110 41460 31116 41472
rect 31071 41432 31116 41460
rect 30469 41423 30527 41429
rect 31110 41420 31116 41432
rect 31168 41420 31174 41472
rect 1104 41370 32016 41392
rect 1104 41318 7288 41370
rect 7340 41318 17592 41370
rect 17644 41318 27896 41370
rect 27948 41318 32016 41370
rect 1104 41296 32016 41318
rect 10318 41256 10324 41268
rect 10279 41228 10324 41256
rect 10318 41216 10324 41228
rect 10376 41216 10382 41268
rect 11882 41216 11888 41268
rect 11940 41216 11946 41268
rect 12710 41216 12716 41268
rect 12768 41256 12774 41268
rect 13449 41259 13507 41265
rect 13449 41256 13461 41259
rect 12768 41228 13461 41256
rect 12768 41216 12774 41228
rect 13449 41225 13461 41228
rect 13495 41225 13507 41259
rect 13449 41219 13507 41225
rect 15102 41216 15108 41268
rect 15160 41256 15166 41268
rect 15657 41259 15715 41265
rect 15657 41256 15669 41259
rect 15160 41228 15669 41256
rect 15160 41216 15166 41228
rect 15657 41225 15669 41228
rect 15703 41225 15715 41259
rect 15657 41219 15715 41225
rect 22278 41216 22284 41268
rect 22336 41256 22342 41268
rect 22336 41228 27384 41256
rect 22336 41216 22342 41228
rect 4430 41188 4436 41200
rect 1412 41160 4436 41188
rect 1412 41132 1440 41160
rect 1394 41120 1400 41132
rect 1355 41092 1400 41120
rect 1394 41080 1400 41092
rect 1452 41080 1458 41132
rect 1670 41129 1676 41132
rect 1664 41083 1676 41129
rect 1728 41120 1734 41132
rect 3804 41129 3832 41160
rect 4430 41148 4436 41160
rect 4488 41148 4494 41200
rect 7006 41188 7012 41200
rect 6380 41160 7012 41188
rect 3789 41123 3847 41129
rect 1728 41092 1764 41120
rect 1670 41080 1676 41083
rect 1728 41080 1734 41092
rect 3789 41089 3801 41123
rect 3835 41089 3847 41123
rect 3789 41083 3847 41089
rect 3878 41080 3884 41132
rect 3936 41120 3942 41132
rect 4045 41123 4103 41129
rect 4045 41120 4057 41123
rect 3936 41092 4057 41120
rect 3936 41080 3942 41092
rect 4045 41089 4057 41092
rect 4091 41089 4103 41123
rect 4448 41120 4476 41148
rect 6380 41129 6408 41160
rect 7006 41148 7012 41160
rect 7064 41148 7070 41200
rect 8656 41191 8714 41197
rect 8656 41157 8668 41191
rect 8702 41188 8714 41191
rect 8938 41188 8944 41200
rect 8702 41160 8944 41188
rect 8702 41157 8714 41160
rect 8656 41151 8714 41157
rect 8938 41148 8944 41160
rect 8996 41148 9002 41200
rect 11900 41188 11928 41216
rect 14553 41191 14611 41197
rect 11624 41160 11928 41188
rect 13648 41160 14504 41188
rect 6365 41123 6423 41129
rect 6365 41120 6377 41123
rect 4448 41092 6377 41120
rect 4045 41083 4103 41089
rect 6365 41089 6377 41092
rect 6411 41089 6423 41123
rect 6365 41083 6423 41089
rect 6632 41123 6690 41129
rect 6632 41089 6644 41123
rect 6678 41120 6690 41123
rect 6914 41120 6920 41132
rect 6678 41092 6920 41120
rect 6678 41089 6690 41092
rect 6632 41083 6690 41089
rect 6914 41080 6920 41092
rect 6972 41080 6978 41132
rect 7024 41120 7052 41148
rect 8389 41123 8447 41129
rect 8389 41120 8401 41123
rect 7024 41092 8401 41120
rect 8389 41089 8401 41092
rect 8435 41089 8447 41123
rect 8389 41083 8447 41089
rect 10505 41123 10563 41129
rect 10505 41089 10517 41123
rect 10551 41120 10563 41123
rect 11514 41120 11520 41132
rect 10551 41092 11520 41120
rect 10551 41089 10563 41092
rect 10505 41083 10563 41089
rect 11514 41080 11520 41092
rect 11572 41080 11578 41132
rect 11624 41129 11652 41160
rect 11609 41123 11667 41129
rect 11609 41089 11621 41123
rect 11655 41089 11667 41123
rect 11609 41083 11667 41089
rect 11876 41123 11934 41129
rect 11876 41089 11888 41123
rect 11922 41120 11934 41123
rect 12618 41120 12624 41132
rect 11922 41092 12624 41120
rect 11922 41089 11934 41092
rect 11876 41083 11934 41089
rect 12618 41080 12624 41092
rect 12676 41080 12682 41132
rect 13078 41080 13084 41132
rect 13136 41120 13142 41132
rect 13648 41129 13676 41160
rect 13633 41123 13691 41129
rect 13633 41120 13645 41123
rect 13136 41092 13645 41120
rect 13136 41080 13142 41092
rect 13633 41089 13645 41092
rect 13679 41089 13691 41123
rect 13633 41083 13691 41089
rect 13909 41123 13967 41129
rect 13909 41089 13921 41123
rect 13955 41089 13967 41123
rect 14090 41120 14096 41132
rect 14051 41092 14096 41120
rect 13909 41083 13967 41089
rect 10781 41055 10839 41061
rect 10781 41021 10793 41055
rect 10827 41052 10839 41055
rect 11054 41052 11060 41064
rect 10827 41024 11060 41052
rect 10827 41021 10839 41024
rect 10781 41015 10839 41021
rect 11054 41012 11060 41024
rect 11112 41012 11118 41064
rect 13924 41052 13952 41083
rect 14090 41080 14096 41092
rect 14148 41080 14154 41132
rect 14476 41120 14504 41160
rect 14553 41157 14565 41191
rect 14599 41188 14611 41191
rect 18322 41188 18328 41200
rect 14599 41160 15884 41188
rect 14599 41157 14611 41160
rect 14553 41151 14611 41157
rect 14734 41120 14740 41132
rect 14476 41092 14740 41120
rect 14734 41080 14740 41092
rect 14792 41080 14798 41132
rect 15013 41123 15071 41129
rect 15013 41089 15025 41123
rect 15059 41089 15071 41123
rect 15013 41083 15071 41089
rect 15197 41123 15255 41129
rect 15197 41089 15209 41123
rect 15243 41120 15255 41123
rect 15746 41120 15752 41132
rect 15243 41092 15752 41120
rect 15243 41089 15255 41092
rect 15197 41083 15255 41089
rect 14642 41052 14648 41064
rect 13924 41024 14648 41052
rect 14642 41012 14648 41024
rect 14700 41052 14706 41064
rect 15028 41052 15056 41083
rect 15746 41080 15752 41092
rect 15804 41080 15810 41132
rect 15856 41129 15884 41160
rect 16684 41160 18328 41188
rect 16684 41129 16712 41160
rect 18322 41148 18328 41160
rect 18380 41188 18386 41200
rect 18380 41160 18552 41188
rect 18380 41148 18386 41160
rect 15841 41123 15899 41129
rect 15841 41089 15853 41123
rect 15887 41089 15899 41123
rect 15841 41083 15899 41089
rect 16669 41123 16727 41129
rect 16669 41089 16681 41123
rect 16715 41089 16727 41123
rect 16669 41083 16727 41089
rect 16758 41080 16764 41132
rect 16816 41120 16822 41132
rect 18524 41129 18552 41160
rect 18598 41148 18604 41200
rect 18656 41188 18662 41200
rect 18754 41191 18812 41197
rect 18754 41188 18766 41191
rect 18656 41160 18766 41188
rect 18656 41148 18662 41160
rect 18754 41157 18766 41160
rect 18800 41157 18812 41191
rect 18754 41151 18812 41157
rect 25308 41191 25366 41197
rect 25308 41157 25320 41191
rect 25354 41188 25366 41191
rect 26050 41188 26056 41200
rect 25354 41160 26056 41188
rect 25354 41157 25366 41160
rect 25308 41151 25366 41157
rect 26050 41148 26056 41160
rect 26108 41148 26114 41200
rect 27246 41197 27252 41200
rect 27240 41188 27252 41197
rect 27207 41160 27252 41188
rect 27240 41151 27252 41160
rect 27246 41148 27252 41151
rect 27304 41148 27310 41200
rect 27356 41188 27384 41228
rect 28736 41228 29316 41256
rect 28736 41188 28764 41228
rect 27356 41160 28764 41188
rect 29288 41188 29316 41228
rect 31294 41188 31300 41200
rect 29288 41160 31300 41188
rect 31294 41148 31300 41160
rect 31352 41148 31358 41200
rect 16925 41123 16983 41129
rect 16925 41120 16937 41123
rect 16816 41092 16937 41120
rect 16816 41080 16822 41092
rect 16925 41089 16937 41092
rect 16971 41089 16983 41123
rect 16925 41083 16983 41089
rect 18509 41123 18567 41129
rect 18509 41089 18521 41123
rect 18555 41120 18567 41123
rect 19242 41120 19248 41132
rect 18555 41092 19248 41120
rect 18555 41089 18567 41092
rect 18509 41083 18567 41089
rect 19242 41080 19248 41092
rect 19300 41080 19306 41132
rect 20254 41080 20260 41132
rect 20312 41120 20318 41132
rect 20625 41123 20683 41129
rect 20625 41120 20637 41123
rect 20312 41092 20637 41120
rect 20312 41080 20318 41092
rect 20625 41089 20637 41092
rect 20671 41089 20683 41123
rect 21266 41120 21272 41132
rect 21227 41092 21272 41120
rect 20625 41083 20683 41089
rect 21266 41080 21272 41092
rect 21324 41080 21330 41132
rect 22088 41123 22146 41129
rect 22088 41089 22100 41123
rect 22134 41120 22146 41123
rect 23661 41123 23719 41129
rect 23661 41120 23673 41123
rect 22134 41092 23673 41120
rect 22134 41089 22146 41092
rect 22088 41083 22146 41089
rect 23661 41089 23673 41092
rect 23707 41089 23719 41123
rect 23661 41083 23719 41089
rect 23845 41123 23903 41129
rect 23845 41089 23857 41123
rect 23891 41089 23903 41123
rect 23845 41083 23903 41089
rect 14700 41024 15056 41052
rect 16117 41055 16175 41061
rect 14700 41012 14706 41024
rect 16117 41021 16129 41055
rect 16163 41021 16175 41055
rect 16117 41015 16175 41021
rect 14090 40944 14096 40996
rect 14148 40984 14154 40996
rect 16132 40984 16160 41015
rect 21634 41012 21640 41064
rect 21692 41052 21698 41064
rect 21821 41055 21879 41061
rect 21821 41052 21833 41055
rect 21692 41024 21833 41052
rect 21692 41012 21698 41024
rect 21821 41021 21833 41024
rect 21867 41021 21879 41055
rect 21821 41015 21879 41021
rect 22830 41012 22836 41064
rect 22888 41052 22894 41064
rect 23860 41052 23888 41083
rect 25774 41080 25780 41132
rect 25832 41120 25838 41132
rect 26973 41123 27031 41129
rect 26973 41120 26985 41123
rect 25832 41092 26985 41120
rect 25832 41080 25838 41092
rect 26973 41089 26985 41092
rect 27019 41089 27031 41123
rect 26973 41083 27031 41089
rect 27614 41080 27620 41132
rect 27672 41120 27678 41132
rect 28718 41120 28724 41132
rect 27672 41092 28724 41120
rect 27672 41080 27678 41092
rect 28718 41080 28724 41092
rect 28776 41120 28782 41132
rect 28813 41123 28871 41129
rect 28813 41120 28825 41123
rect 28776 41092 28825 41120
rect 28776 41080 28782 41092
rect 28813 41089 28825 41092
rect 28859 41089 28871 41123
rect 28813 41083 28871 41089
rect 28902 41080 28908 41132
rect 28960 41120 28966 41132
rect 29069 41123 29127 41129
rect 29069 41120 29081 41123
rect 28960 41092 29081 41120
rect 28960 41080 28966 41092
rect 29069 41089 29081 41092
rect 29115 41089 29127 41123
rect 29069 41083 29127 41089
rect 30837 41123 30895 41129
rect 30837 41089 30849 41123
rect 30883 41089 30895 41123
rect 30837 41083 30895 41089
rect 22888 41024 23888 41052
rect 24121 41055 24179 41061
rect 22888 41012 22894 41024
rect 24121 41021 24133 41055
rect 24167 41052 24179 41055
rect 24302 41052 24308 41064
rect 24167 41024 24308 41052
rect 24167 41021 24179 41024
rect 24121 41015 24179 41021
rect 14148 40956 16160 40984
rect 14148 40944 14154 40956
rect 19794 40944 19800 40996
rect 19852 40984 19858 40996
rect 20441 40987 20499 40993
rect 20441 40984 20453 40987
rect 19852 40956 20453 40984
rect 19852 40944 19858 40956
rect 20441 40953 20453 40956
rect 20487 40953 20499 40987
rect 20441 40947 20499 40953
rect 23566 40944 23572 40996
rect 23624 40984 23630 40996
rect 24136 40984 24164 41015
rect 24302 41012 24308 41024
rect 24360 41012 24366 41064
rect 25038 41052 25044 41064
rect 24999 41024 25044 41052
rect 25038 41012 25044 41024
rect 25096 41012 25102 41064
rect 29914 41012 29920 41064
rect 29972 41052 29978 41064
rect 30852 41052 30880 41083
rect 29972 41024 30880 41052
rect 29972 41012 29978 41024
rect 23624 40956 24164 40984
rect 30193 40987 30251 40993
rect 23624 40944 23630 40956
rect 30193 40953 30205 40987
rect 30239 40953 30251 40987
rect 30193 40947 30251 40953
rect 2777 40919 2835 40925
rect 2777 40885 2789 40919
rect 2823 40916 2835 40919
rect 3234 40916 3240 40928
rect 2823 40888 3240 40916
rect 2823 40885 2835 40888
rect 2777 40879 2835 40885
rect 3234 40876 3240 40888
rect 3292 40876 3298 40928
rect 5169 40919 5227 40925
rect 5169 40885 5181 40919
rect 5215 40916 5227 40919
rect 5258 40916 5264 40928
rect 5215 40888 5264 40916
rect 5215 40885 5227 40888
rect 5169 40879 5227 40885
rect 5258 40876 5264 40888
rect 5316 40876 5322 40928
rect 7745 40919 7803 40925
rect 7745 40885 7757 40919
rect 7791 40916 7803 40919
rect 8202 40916 8208 40928
rect 7791 40888 8208 40916
rect 7791 40885 7803 40888
rect 7745 40879 7803 40885
rect 8202 40876 8208 40888
rect 8260 40876 8266 40928
rect 9674 40876 9680 40928
rect 9732 40916 9738 40928
rect 9769 40919 9827 40925
rect 9769 40916 9781 40919
rect 9732 40888 9781 40916
rect 9732 40876 9738 40888
rect 9769 40885 9781 40888
rect 9815 40885 9827 40919
rect 9769 40879 9827 40885
rect 10689 40919 10747 40925
rect 10689 40885 10701 40919
rect 10735 40916 10747 40919
rect 10778 40916 10784 40928
rect 10735 40888 10784 40916
rect 10735 40885 10747 40888
rect 10689 40879 10747 40885
rect 10778 40876 10784 40888
rect 10836 40876 10842 40928
rect 12986 40916 12992 40928
rect 12899 40888 12992 40916
rect 12986 40876 12992 40888
rect 13044 40916 13050 40928
rect 13446 40916 13452 40928
rect 13044 40888 13452 40916
rect 13044 40876 13050 40888
rect 13446 40876 13452 40888
rect 13504 40876 13510 40928
rect 15654 40876 15660 40928
rect 15712 40916 15718 40928
rect 16022 40916 16028 40928
rect 15712 40888 16028 40916
rect 15712 40876 15718 40888
rect 16022 40876 16028 40888
rect 16080 40876 16086 40928
rect 18046 40916 18052 40928
rect 18007 40888 18052 40916
rect 18046 40876 18052 40888
rect 18104 40876 18110 40928
rect 19518 40876 19524 40928
rect 19576 40916 19582 40928
rect 19889 40919 19947 40925
rect 19889 40916 19901 40919
rect 19576 40888 19901 40916
rect 19576 40876 19582 40888
rect 19889 40885 19901 40888
rect 19935 40885 19947 40919
rect 21082 40916 21088 40928
rect 21043 40888 21088 40916
rect 19889 40879 19947 40885
rect 21082 40876 21088 40888
rect 21140 40876 21146 40928
rect 23201 40919 23259 40925
rect 23201 40885 23213 40919
rect 23247 40916 23259 40919
rect 23750 40916 23756 40928
rect 23247 40888 23756 40916
rect 23247 40885 23259 40888
rect 23201 40879 23259 40885
rect 23750 40876 23756 40888
rect 23808 40876 23814 40928
rect 24026 40916 24032 40928
rect 23987 40888 24032 40916
rect 24026 40876 24032 40888
rect 24084 40876 24090 40928
rect 26326 40876 26332 40928
rect 26384 40916 26390 40928
rect 26421 40919 26479 40925
rect 26421 40916 26433 40919
rect 26384 40888 26433 40916
rect 26384 40876 26390 40888
rect 26421 40885 26433 40888
rect 26467 40916 26479 40919
rect 27338 40916 27344 40928
rect 26467 40888 27344 40916
rect 26467 40885 26479 40888
rect 26421 40879 26479 40885
rect 27338 40876 27344 40888
rect 27396 40876 27402 40928
rect 27706 40876 27712 40928
rect 27764 40916 27770 40928
rect 28353 40919 28411 40925
rect 28353 40916 28365 40919
rect 27764 40888 28365 40916
rect 27764 40876 27770 40888
rect 28353 40885 28365 40888
rect 28399 40916 28411 40919
rect 28810 40916 28816 40928
rect 28399 40888 28816 40916
rect 28399 40885 28411 40888
rect 28353 40879 28411 40885
rect 28810 40876 28816 40888
rect 28868 40876 28874 40928
rect 28994 40876 29000 40928
rect 29052 40916 29058 40928
rect 30208 40916 30236 40947
rect 29052 40888 30236 40916
rect 29052 40876 29058 40888
rect 30466 40876 30472 40928
rect 30524 40916 30530 40928
rect 30653 40919 30711 40925
rect 30653 40916 30665 40919
rect 30524 40888 30665 40916
rect 30524 40876 30530 40888
rect 30653 40885 30665 40888
rect 30699 40885 30711 40919
rect 30653 40879 30711 40885
rect 1104 40826 32016 40848
rect 0 40780 800 40794
rect 0 40752 980 40780
rect 1104 40774 2136 40826
rect 2188 40774 12440 40826
rect 12492 40774 22744 40826
rect 22796 40774 32016 40826
rect 32320 40780 33120 40794
rect 1104 40752 32016 40774
rect 32048 40752 33120 40780
rect 0 40738 800 40752
rect 952 40712 980 40752
rect 1486 40712 1492 40724
rect 952 40684 1492 40712
rect 1486 40672 1492 40684
rect 1544 40672 1550 40724
rect 1670 40712 1676 40724
rect 1631 40684 1676 40712
rect 1670 40672 1676 40684
rect 1728 40672 1734 40724
rect 2866 40672 2872 40724
rect 2924 40712 2930 40724
rect 3789 40715 3847 40721
rect 3789 40712 3801 40715
rect 2924 40684 3801 40712
rect 2924 40672 2930 40684
rect 3789 40681 3801 40684
rect 3835 40681 3847 40715
rect 7006 40712 7012 40724
rect 6967 40684 7012 40712
rect 3789 40675 3847 40681
rect 7006 40672 7012 40684
rect 7064 40672 7070 40724
rect 11882 40712 11888 40724
rect 9416 40684 11888 40712
rect 6914 40604 6920 40656
rect 6972 40644 6978 40656
rect 7929 40647 7987 40653
rect 7929 40644 7941 40647
rect 6972 40616 7941 40644
rect 6972 40604 6978 40616
rect 7929 40613 7941 40616
rect 7975 40613 7987 40647
rect 7929 40607 7987 40613
rect 2133 40579 2191 40585
rect 2133 40545 2145 40579
rect 2179 40576 2191 40579
rect 2866 40576 2872 40588
rect 2179 40548 2872 40576
rect 2179 40545 2191 40548
rect 2133 40539 2191 40545
rect 2866 40536 2872 40548
rect 2924 40536 2930 40588
rect 4614 40576 4620 40588
rect 3068 40548 4620 40576
rect 1857 40511 1915 40517
rect 1857 40477 1869 40511
rect 1903 40477 1915 40511
rect 1857 40471 1915 40477
rect 2041 40511 2099 40517
rect 2041 40477 2053 40511
rect 2087 40508 2099 40511
rect 2682 40508 2688 40520
rect 2087 40480 2688 40508
rect 2087 40477 2099 40480
rect 2041 40471 2099 40477
rect 1872 40440 1900 40471
rect 2682 40468 2688 40480
rect 2740 40468 2746 40520
rect 3068 40517 3096 40548
rect 2777 40511 2835 40517
rect 2777 40477 2789 40511
rect 2823 40477 2835 40511
rect 2777 40471 2835 40477
rect 3053 40511 3111 40517
rect 3053 40477 3065 40511
rect 3099 40477 3111 40511
rect 3234 40508 3240 40520
rect 3195 40480 3240 40508
rect 3053 40471 3111 40477
rect 2593 40443 2651 40449
rect 2593 40440 2605 40443
rect 1872 40412 2605 40440
rect 2593 40409 2605 40412
rect 2639 40409 2651 40443
rect 2792 40440 2820 40471
rect 3234 40468 3240 40480
rect 3292 40468 3298 40520
rect 3510 40468 3516 40520
rect 3568 40508 3574 40520
rect 3973 40511 4031 40517
rect 3973 40508 3985 40511
rect 3568 40480 3985 40508
rect 3568 40468 3574 40480
rect 3973 40477 3985 40480
rect 4019 40508 4031 40511
rect 4062 40508 4068 40520
rect 4019 40480 4068 40508
rect 4019 40477 4031 40480
rect 3973 40471 4031 40477
rect 4062 40468 4068 40480
rect 4120 40468 4126 40520
rect 4264 40517 4292 40548
rect 4614 40536 4620 40548
rect 4672 40576 4678 40588
rect 4982 40576 4988 40588
rect 4672 40548 4988 40576
rect 4672 40536 4678 40548
rect 4982 40536 4988 40548
rect 5040 40536 5046 40588
rect 5350 40536 5356 40588
rect 5408 40576 5414 40588
rect 9416 40585 9444 40684
rect 11882 40672 11888 40684
rect 11940 40672 11946 40724
rect 16390 40712 16396 40724
rect 16351 40684 16396 40712
rect 16390 40672 16396 40684
rect 16448 40672 16454 40724
rect 22189 40715 22247 40721
rect 22189 40681 22201 40715
rect 22235 40712 22247 40715
rect 22830 40712 22836 40724
rect 22235 40684 22836 40712
rect 22235 40681 22247 40684
rect 22189 40675 22247 40681
rect 22830 40672 22836 40684
rect 22888 40672 22894 40724
rect 23290 40712 23296 40724
rect 23251 40684 23296 40712
rect 23290 40672 23296 40684
rect 23348 40672 23354 40724
rect 26418 40672 26424 40724
rect 26476 40712 26482 40724
rect 27341 40715 27399 40721
rect 27341 40712 27353 40715
rect 26476 40684 27353 40712
rect 26476 40672 26482 40684
rect 27341 40681 27353 40684
rect 27387 40681 27399 40715
rect 27341 40675 27399 40681
rect 28445 40715 28503 40721
rect 28445 40681 28457 40715
rect 28491 40712 28503 40715
rect 28902 40712 28908 40724
rect 28491 40684 28908 40712
rect 28491 40681 28503 40684
rect 28445 40675 28503 40681
rect 28902 40672 28908 40684
rect 28960 40672 28966 40724
rect 29914 40712 29920 40724
rect 29012 40684 29920 40712
rect 17218 40644 17224 40656
rect 15948 40616 17224 40644
rect 8389 40579 8447 40585
rect 8389 40576 8401 40579
rect 5408 40548 8401 40576
rect 5408 40536 5414 40548
rect 8389 40545 8401 40548
rect 8435 40545 8447 40579
rect 8389 40539 8447 40545
rect 9401 40579 9459 40585
rect 9401 40545 9413 40579
rect 9447 40545 9459 40579
rect 9401 40539 9459 40545
rect 4249 40511 4307 40517
rect 4249 40477 4261 40511
rect 4295 40477 4307 40511
rect 4249 40471 4307 40477
rect 4338 40468 4344 40520
rect 4396 40508 4402 40520
rect 4433 40511 4491 40517
rect 4433 40508 4445 40511
rect 4396 40480 4445 40508
rect 4396 40468 4402 40480
rect 4433 40477 4445 40480
rect 4479 40508 4491 40511
rect 5166 40508 5172 40520
rect 4479 40480 5172 40508
rect 4479 40477 4491 40480
rect 4433 40471 4491 40477
rect 5166 40468 5172 40480
rect 5224 40468 5230 40520
rect 7558 40468 7564 40520
rect 7616 40508 7622 40520
rect 8113 40511 8171 40517
rect 8113 40508 8125 40511
rect 7616 40480 8125 40508
rect 7616 40468 7622 40480
rect 8113 40477 8125 40480
rect 8159 40477 8171 40511
rect 8113 40471 8171 40477
rect 8297 40511 8355 40517
rect 8297 40477 8309 40511
rect 8343 40508 8355 40511
rect 8570 40508 8576 40520
rect 8343 40480 8576 40508
rect 8343 40477 8355 40480
rect 8297 40471 8355 40477
rect 8570 40468 8576 40480
rect 8628 40508 8634 40520
rect 8938 40508 8944 40520
rect 8628 40480 8944 40508
rect 8628 40468 8634 40480
rect 8938 40468 8944 40480
rect 8996 40468 9002 40520
rect 11422 40508 11428 40520
rect 11383 40480 11428 40508
rect 11422 40468 11428 40480
rect 11480 40468 11486 40520
rect 11701 40511 11759 40517
rect 11701 40477 11713 40511
rect 11747 40508 11759 40511
rect 11790 40508 11796 40520
rect 11747 40480 11796 40508
rect 11747 40477 11759 40480
rect 11701 40471 11759 40477
rect 11790 40468 11796 40480
rect 11848 40468 11854 40520
rect 11885 40511 11943 40517
rect 11885 40477 11897 40511
rect 11931 40477 11943 40511
rect 11885 40471 11943 40477
rect 12989 40511 13047 40517
rect 12989 40477 13001 40511
rect 13035 40508 13047 40511
rect 13078 40508 13084 40520
rect 13035 40480 13084 40508
rect 13035 40477 13047 40480
rect 12989 40471 13047 40477
rect 3528 40440 3556 40468
rect 2792 40412 3556 40440
rect 5721 40443 5779 40449
rect 2593 40403 2651 40409
rect 5721 40409 5733 40443
rect 5767 40440 5779 40443
rect 9668 40443 9726 40449
rect 5767 40412 8616 40440
rect 5767 40409 5779 40412
rect 5721 40403 5779 40409
rect 8588 40372 8616 40412
rect 9668 40409 9680 40443
rect 9714 40440 9726 40443
rect 9950 40440 9956 40452
rect 9714 40412 9956 40440
rect 9714 40409 9726 40412
rect 9668 40403 9726 40409
rect 9950 40400 9956 40412
rect 10008 40400 10014 40452
rect 11054 40440 11060 40452
rect 10796 40412 11060 40440
rect 10594 40372 10600 40384
rect 8588 40344 10600 40372
rect 10594 40332 10600 40344
rect 10652 40332 10658 40384
rect 10796 40381 10824 40412
rect 11054 40400 11060 40412
rect 11112 40440 11118 40452
rect 11606 40440 11612 40452
rect 11112 40412 11612 40440
rect 11112 40400 11118 40412
rect 11606 40400 11612 40412
rect 11664 40440 11670 40452
rect 11900 40440 11928 40471
rect 13078 40468 13084 40480
rect 13136 40468 13142 40520
rect 13265 40511 13323 40517
rect 13265 40477 13277 40511
rect 13311 40477 13323 40511
rect 13446 40508 13452 40520
rect 13407 40480 13452 40508
rect 13265 40471 13323 40477
rect 11664 40412 11928 40440
rect 13280 40440 13308 40471
rect 13446 40468 13452 40480
rect 13504 40468 13510 40520
rect 13998 40468 14004 40520
rect 14056 40508 14062 40520
rect 14553 40511 14611 40517
rect 14553 40508 14565 40511
rect 14056 40480 14565 40508
rect 14056 40468 14062 40480
rect 14553 40477 14565 40480
rect 14599 40477 14611 40511
rect 14553 40471 14611 40477
rect 14642 40440 14648 40452
rect 13280 40412 14648 40440
rect 11664 40400 11670 40412
rect 14642 40400 14648 40412
rect 14700 40400 14706 40452
rect 14820 40443 14878 40449
rect 14820 40409 14832 40443
rect 14866 40440 14878 40443
rect 15286 40440 15292 40452
rect 14866 40412 15292 40440
rect 14866 40409 14878 40412
rect 14820 40403 14878 40409
rect 15286 40400 15292 40412
rect 15344 40400 15350 40452
rect 10781 40375 10839 40381
rect 10781 40341 10793 40375
rect 10827 40341 10839 40375
rect 10781 40335 10839 40341
rect 10870 40332 10876 40384
rect 10928 40372 10934 40384
rect 11241 40375 11299 40381
rect 11241 40372 11253 40375
rect 10928 40344 11253 40372
rect 10928 40332 10934 40344
rect 11241 40341 11253 40344
rect 11287 40341 11299 40375
rect 12802 40372 12808 40384
rect 12763 40344 12808 40372
rect 11241 40335 11299 40341
rect 12802 40332 12808 40344
rect 12860 40332 12866 40384
rect 15470 40332 15476 40384
rect 15528 40372 15534 40384
rect 15948 40381 15976 40616
rect 17218 40604 17224 40616
rect 17276 40604 17282 40656
rect 25590 40604 25596 40656
rect 25648 40644 25654 40656
rect 26050 40644 26056 40656
rect 25648 40616 26056 40644
rect 25648 40604 25654 40616
rect 26050 40604 26056 40616
rect 26108 40644 26114 40656
rect 26108 40616 26924 40644
rect 26108 40604 26114 40616
rect 18230 40576 18236 40588
rect 16592 40548 18236 40576
rect 16592 40520 16620 40548
rect 16574 40508 16580 40520
rect 16487 40480 16580 40508
rect 16574 40468 16580 40480
rect 16632 40468 16638 40520
rect 16853 40511 16911 40517
rect 16853 40477 16865 40511
rect 16899 40477 16911 40511
rect 16853 40471 16911 40477
rect 17037 40511 17095 40517
rect 17037 40477 17049 40511
rect 17083 40508 17095 40511
rect 17310 40508 17316 40520
rect 17083 40480 17316 40508
rect 17083 40477 17095 40480
rect 17037 40471 17095 40477
rect 16868 40440 16896 40471
rect 17310 40468 17316 40480
rect 17368 40468 17374 40520
rect 17696 40517 17724 40548
rect 18230 40536 18236 40548
rect 18288 40536 18294 40588
rect 19242 40576 19248 40588
rect 19203 40548 19248 40576
rect 19242 40536 19248 40548
rect 19300 40536 19306 40588
rect 23014 40576 23020 40588
rect 22388 40548 23020 40576
rect 17681 40511 17739 40517
rect 17681 40477 17693 40511
rect 17727 40477 17739 40511
rect 17681 40471 17739 40477
rect 17957 40511 18015 40517
rect 17957 40477 17969 40511
rect 18003 40477 18015 40511
rect 17957 40471 18015 40477
rect 17126 40440 17132 40452
rect 16868 40412 17132 40440
rect 17126 40400 17132 40412
rect 17184 40440 17190 40452
rect 17972 40440 18000 40471
rect 18046 40468 18052 40520
rect 18104 40508 18110 40520
rect 18141 40511 18199 40517
rect 18141 40508 18153 40511
rect 18104 40480 18153 40508
rect 18104 40468 18110 40480
rect 18141 40477 18153 40480
rect 18187 40477 18199 40511
rect 18141 40471 18199 40477
rect 19150 40468 19156 40520
rect 19208 40508 19214 40520
rect 19501 40511 19559 40517
rect 19501 40508 19513 40511
rect 19208 40480 19513 40508
rect 19208 40468 19214 40480
rect 19501 40477 19513 40480
rect 19547 40477 19559 40511
rect 19501 40471 19559 40477
rect 20714 40468 20720 40520
rect 20772 40508 20778 40520
rect 21729 40511 21787 40517
rect 21729 40508 21741 40511
rect 20772 40480 21741 40508
rect 20772 40468 20778 40480
rect 21729 40477 21741 40480
rect 21775 40508 21787 40511
rect 22278 40508 22284 40520
rect 21775 40480 22284 40508
rect 21775 40477 21787 40480
rect 21729 40471 21787 40477
rect 22278 40468 22284 40480
rect 22336 40468 22342 40520
rect 22388 40517 22416 40548
rect 23014 40536 23020 40548
rect 23072 40536 23078 40588
rect 24026 40576 24032 40588
rect 23676 40548 24032 40576
rect 22373 40511 22431 40517
rect 22373 40477 22385 40511
rect 22419 40477 22431 40511
rect 22373 40471 22431 40477
rect 22649 40511 22707 40517
rect 22649 40477 22661 40511
rect 22695 40477 22707 40511
rect 22649 40471 22707 40477
rect 22833 40511 22891 40517
rect 22833 40477 22845 40511
rect 22879 40477 22891 40511
rect 23474 40508 23480 40520
rect 23435 40480 23480 40508
rect 22833 40471 22891 40477
rect 18506 40440 18512 40452
rect 17184 40412 18512 40440
rect 17184 40400 17190 40412
rect 18506 40400 18512 40412
rect 18564 40400 18570 40452
rect 22186 40400 22192 40452
rect 22244 40440 22250 40452
rect 22664 40440 22692 40471
rect 22244 40412 22692 40440
rect 22848 40440 22876 40471
rect 23474 40468 23480 40480
rect 23532 40468 23538 40520
rect 23566 40468 23572 40520
rect 23624 40508 23630 40520
rect 23676 40517 23704 40548
rect 24026 40536 24032 40548
rect 24084 40536 24090 40588
rect 23661 40511 23719 40517
rect 23661 40508 23673 40511
rect 23624 40480 23673 40508
rect 23624 40468 23630 40480
rect 23661 40477 23673 40480
rect 23707 40477 23719 40511
rect 23661 40471 23719 40477
rect 23750 40468 23756 40520
rect 23808 40508 23814 40520
rect 24394 40508 24400 40520
rect 23808 40480 23853 40508
rect 24307 40480 24400 40508
rect 23808 40468 23814 40480
rect 24394 40468 24400 40480
rect 24452 40508 24458 40520
rect 25038 40508 25044 40520
rect 24452 40480 25044 40508
rect 24452 40468 24458 40480
rect 25038 40468 25044 40480
rect 25096 40508 25102 40520
rect 25774 40508 25780 40520
rect 25096 40480 25780 40508
rect 25096 40468 25102 40480
rect 25774 40468 25780 40480
rect 25832 40468 25838 40520
rect 26234 40468 26240 40520
rect 26292 40508 26298 40520
rect 26421 40511 26479 40517
rect 26421 40508 26433 40511
rect 26292 40480 26433 40508
rect 26292 40468 26298 40480
rect 26421 40477 26433 40480
rect 26467 40477 26479 40511
rect 26694 40508 26700 40520
rect 26655 40480 26700 40508
rect 26421 40471 26479 40477
rect 26694 40468 26700 40480
rect 26752 40468 26758 40520
rect 26896 40517 26924 40616
rect 26970 40604 26976 40656
rect 27028 40644 27034 40656
rect 29012 40644 29040 40684
rect 29914 40672 29920 40684
rect 29972 40672 29978 40724
rect 30282 40672 30288 40724
rect 30340 40712 30346 40724
rect 32048 40712 32076 40752
rect 32320 40738 33120 40752
rect 30340 40684 32076 40712
rect 30340 40672 30346 40684
rect 27028 40616 29040 40644
rect 27028 40604 27034 40616
rect 27338 40536 27344 40588
rect 27396 40576 27402 40588
rect 27396 40548 28028 40576
rect 27396 40536 27402 40548
rect 26881 40511 26939 40517
rect 26881 40477 26893 40511
rect 26927 40477 26939 40511
rect 26881 40471 26939 40477
rect 26970 40468 26976 40520
rect 27028 40508 27034 40520
rect 27525 40511 27583 40517
rect 27525 40508 27537 40511
rect 27028 40480 27537 40508
rect 27028 40468 27034 40480
rect 27525 40477 27537 40480
rect 27571 40477 27583 40511
rect 27798 40508 27804 40520
rect 27759 40480 27804 40508
rect 27525 40471 27583 40477
rect 27798 40468 27804 40480
rect 27856 40468 27862 40520
rect 28000 40517 28028 40548
rect 28718 40536 28724 40588
rect 28776 40576 28782 40588
rect 29546 40576 29552 40588
rect 28776 40548 29552 40576
rect 28776 40536 28782 40548
rect 29546 40536 29552 40548
rect 29604 40536 29610 40588
rect 27985 40511 28043 40517
rect 27985 40477 27997 40511
rect 28031 40477 28043 40511
rect 27985 40471 28043 40477
rect 28258 40468 28264 40520
rect 28316 40508 28322 40520
rect 28442 40508 28448 40520
rect 28316 40480 28448 40508
rect 28316 40468 28322 40480
rect 28442 40468 28448 40480
rect 28500 40468 28506 40520
rect 28629 40511 28687 40517
rect 28629 40508 28641 40511
rect 28552 40480 28641 40508
rect 23768 40440 23796 40468
rect 22848 40412 23796 40440
rect 22244 40400 22250 40412
rect 24486 40400 24492 40452
rect 24544 40440 24550 40452
rect 24642 40443 24700 40449
rect 24642 40440 24654 40443
rect 24544 40412 24654 40440
rect 24544 40400 24550 40412
rect 24642 40409 24654 40412
rect 24688 40409 24700 40443
rect 24642 40403 24700 40409
rect 28074 40400 28080 40452
rect 28132 40440 28138 40452
rect 28552 40440 28580 40480
rect 28629 40477 28641 40480
rect 28675 40477 28687 40511
rect 28810 40508 28816 40520
rect 28771 40480 28816 40508
rect 28629 40471 28687 40477
rect 28810 40468 28816 40480
rect 28868 40468 28874 40520
rect 28902 40468 28908 40520
rect 28960 40508 28966 40520
rect 28960 40480 29005 40508
rect 28960 40468 28966 40480
rect 29638 40468 29644 40520
rect 29696 40508 29702 40520
rect 29805 40511 29863 40517
rect 29805 40508 29817 40511
rect 29696 40480 29817 40508
rect 29696 40468 29702 40480
rect 29805 40477 29817 40480
rect 29851 40477 29863 40511
rect 29805 40471 29863 40477
rect 28132 40412 28580 40440
rect 28132 40400 28138 40412
rect 15933 40375 15991 40381
rect 15933 40372 15945 40375
rect 15528 40344 15945 40372
rect 15528 40332 15534 40344
rect 15933 40341 15945 40344
rect 15979 40341 15991 40375
rect 15933 40335 15991 40341
rect 16942 40332 16948 40384
rect 17000 40372 17006 40384
rect 17497 40375 17555 40381
rect 17497 40372 17509 40375
rect 17000 40344 17509 40372
rect 17000 40332 17006 40344
rect 17497 40341 17509 40344
rect 17543 40341 17555 40375
rect 17497 40335 17555 40341
rect 19426 40332 19432 40384
rect 19484 40372 19490 40384
rect 20625 40375 20683 40381
rect 20625 40372 20637 40375
rect 19484 40344 20637 40372
rect 19484 40332 19490 40344
rect 20625 40341 20637 40344
rect 20671 40341 20683 40375
rect 20625 40335 20683 40341
rect 21545 40375 21603 40381
rect 21545 40341 21557 40375
rect 21591 40372 21603 40375
rect 22002 40372 22008 40384
rect 21591 40344 22008 40372
rect 21591 40341 21603 40344
rect 21545 40335 21603 40341
rect 22002 40332 22008 40344
rect 22060 40332 22066 40384
rect 25777 40375 25835 40381
rect 25777 40341 25789 40375
rect 25823 40372 25835 40375
rect 25866 40372 25872 40384
rect 25823 40344 25872 40372
rect 25823 40341 25835 40344
rect 25777 40335 25835 40341
rect 25866 40332 25872 40344
rect 25924 40332 25930 40384
rect 26237 40375 26295 40381
rect 26237 40341 26249 40375
rect 26283 40372 26295 40375
rect 28442 40372 28448 40384
rect 26283 40344 28448 40372
rect 26283 40341 26295 40344
rect 26237 40335 26295 40341
rect 28442 40332 28448 40344
rect 28500 40332 28506 40384
rect 30926 40372 30932 40384
rect 30887 40344 30932 40372
rect 30926 40332 30932 40344
rect 30984 40332 30990 40384
rect 1104 40282 32016 40304
rect 1104 40230 7288 40282
rect 7340 40230 17592 40282
rect 17644 40230 27896 40282
rect 27948 40230 32016 40282
rect 1104 40208 32016 40230
rect 3329 40171 3387 40177
rect 3329 40137 3341 40171
rect 3375 40168 3387 40171
rect 3970 40168 3976 40180
rect 3375 40140 3976 40168
rect 3375 40137 3387 40140
rect 3329 40131 3387 40137
rect 3970 40128 3976 40140
rect 4028 40128 4034 40180
rect 5350 40128 5356 40180
rect 5408 40168 5414 40180
rect 5813 40171 5871 40177
rect 5813 40168 5825 40171
rect 5408 40140 5825 40168
rect 5408 40128 5414 40140
rect 5813 40137 5825 40140
rect 5859 40168 5871 40171
rect 7558 40168 7564 40180
rect 5859 40140 6868 40168
rect 7519 40140 7564 40168
rect 5859 40137 5871 40140
rect 5813 40131 5871 40137
rect 5258 40100 5264 40112
rect 3988 40072 5264 40100
rect 1664 40035 1722 40041
rect 1664 40001 1676 40035
rect 1710 40032 1722 40035
rect 2590 40032 2596 40044
rect 1710 40004 2596 40032
rect 1710 40001 1722 40004
rect 1664 39995 1722 40001
rect 2590 39992 2596 40004
rect 2648 39992 2654 40044
rect 3510 40032 3516 40044
rect 3471 40004 3516 40032
rect 3510 39992 3516 40004
rect 3568 39992 3574 40044
rect 3988 40041 4016 40072
rect 5258 40060 5264 40072
rect 5316 40060 5322 40112
rect 6840 40109 6868 40140
rect 7558 40128 7564 40140
rect 7616 40128 7622 40180
rect 8849 40171 8907 40177
rect 8849 40137 8861 40171
rect 8895 40168 8907 40171
rect 9122 40168 9128 40180
rect 8895 40140 9128 40168
rect 8895 40137 8907 40140
rect 8849 40131 8907 40137
rect 9122 40128 9128 40140
rect 9180 40128 9186 40180
rect 9950 40168 9956 40180
rect 9911 40140 9956 40168
rect 9950 40128 9956 40140
rect 10008 40128 10014 40180
rect 11514 40168 11520 40180
rect 11475 40140 11520 40168
rect 11514 40128 11520 40140
rect 11572 40128 11578 40180
rect 13740 40140 18000 40168
rect 6825 40103 6883 40109
rect 6825 40069 6837 40103
rect 6871 40069 6883 40103
rect 7926 40100 7932 40112
rect 6825 40063 6883 40069
rect 7760 40072 7932 40100
rect 3789 40035 3847 40041
rect 3789 40001 3801 40035
rect 3835 40001 3847 40035
rect 3789 39995 3847 40001
rect 3973 40035 4031 40041
rect 3973 40001 3985 40035
rect 4019 40001 4031 40035
rect 4430 40032 4436 40044
rect 4391 40004 4436 40032
rect 3973 39995 4031 40001
rect 1394 39964 1400 39976
rect 1355 39936 1400 39964
rect 1394 39924 1400 39936
rect 1452 39924 1458 39976
rect 3804 39964 3832 39995
rect 4430 39992 4436 40004
rect 4488 39992 4494 40044
rect 4522 39992 4528 40044
rect 4580 39992 4586 40044
rect 4700 40035 4758 40041
rect 4700 40001 4712 40035
rect 4746 40032 4758 40035
rect 5810 40032 5816 40044
rect 4746 40004 5816 40032
rect 4746 40001 4758 40004
rect 4700 39995 4758 40001
rect 5810 39992 5816 40004
rect 5868 39992 5874 40044
rect 6549 40035 6607 40041
rect 6549 40001 6561 40035
rect 6595 40001 6607 40035
rect 6730 40032 6736 40044
rect 6691 40004 6736 40032
rect 6549 39995 6607 40001
rect 4540 39964 4568 39992
rect 3804 39936 4568 39964
rect 6564 39964 6592 39995
rect 6730 39992 6736 40004
rect 6788 39992 6794 40044
rect 6917 40035 6975 40041
rect 6917 40001 6929 40035
rect 6963 40032 6975 40035
rect 7098 40032 7104 40044
rect 6963 40004 7104 40032
rect 6963 40001 6975 40004
rect 6917 39995 6975 40001
rect 7098 39992 7104 40004
rect 7156 39992 7162 40044
rect 7760 40041 7788 40072
rect 7926 40060 7932 40072
rect 7984 40100 7990 40112
rect 7984 40072 9076 40100
rect 7984 40060 7990 40072
rect 9048 40044 9076 40072
rect 10226 40060 10232 40112
rect 10284 40100 10290 40112
rect 10410 40100 10416 40112
rect 10284 40072 10416 40100
rect 10284 40060 10290 40072
rect 10410 40060 10416 40072
rect 10468 40100 10474 40112
rect 13740 40100 13768 40140
rect 10468 40072 13768 40100
rect 10468 40060 10474 40072
rect 7745 40035 7803 40041
rect 7745 40001 7757 40035
rect 7791 40001 7803 40035
rect 7745 39995 7803 40001
rect 8021 40035 8079 40041
rect 8021 40001 8033 40035
rect 8067 40001 8079 40035
rect 8202 40032 8208 40044
rect 8163 40004 8208 40032
rect 8021 39995 8079 40001
rect 8036 39964 8064 39995
rect 8202 39992 8208 40004
rect 8260 39992 8266 40044
rect 9030 40032 9036 40044
rect 8991 40004 9036 40032
rect 9030 39992 9036 40004
rect 9088 39992 9094 40044
rect 9309 40035 9367 40041
rect 9309 40001 9321 40035
rect 9355 40001 9367 40035
rect 9309 39995 9367 40001
rect 9493 40035 9551 40041
rect 9493 40001 9505 40035
rect 9539 40032 9551 40035
rect 9674 40032 9680 40044
rect 9539 40004 9680 40032
rect 9539 40001 9551 40004
rect 9493 39995 9551 40001
rect 8294 39964 8300 39976
rect 6564 39936 6960 39964
rect 8036 39936 8300 39964
rect 6932 39896 6960 39936
rect 8294 39924 8300 39936
rect 8352 39964 8358 39976
rect 9324 39964 9352 39995
rect 9674 39992 9680 40004
rect 9732 39992 9738 40044
rect 10137 40035 10195 40041
rect 10137 40001 10149 40035
rect 10183 40032 10195 40035
rect 10870 40032 10876 40044
rect 10183 40004 10876 40032
rect 10183 40001 10195 40004
rect 10137 39995 10195 40001
rect 10870 39992 10876 40004
rect 10928 39992 10934 40044
rect 11422 39992 11428 40044
rect 11480 40032 11486 40044
rect 11701 40035 11759 40041
rect 11701 40032 11713 40035
rect 11480 40004 11713 40032
rect 11480 39992 11486 40004
rect 11701 40001 11713 40004
rect 11747 40001 11759 40035
rect 11701 39995 11759 40001
rect 8352 39936 9352 39964
rect 9692 39964 9720 39992
rect 10413 39967 10471 39973
rect 10413 39964 10425 39967
rect 9692 39936 10425 39964
rect 8352 39924 8358 39936
rect 10413 39933 10425 39936
rect 10459 39933 10471 39967
rect 10413 39927 10471 39933
rect 8202 39896 8208 39908
rect 6932 39868 8208 39896
rect 8202 39856 8208 39868
rect 8260 39856 8266 39908
rect 11716 39896 11744 39995
rect 11790 39992 11796 40044
rect 11848 40032 11854 40044
rect 11977 40035 12035 40041
rect 11977 40032 11989 40035
rect 11848 40004 11989 40032
rect 11848 39992 11854 40004
rect 11977 40001 11989 40004
rect 12023 40001 12035 40035
rect 11977 39995 12035 40001
rect 12161 40035 12219 40041
rect 12161 40001 12173 40035
rect 12207 40032 12219 40035
rect 12250 40032 12256 40044
rect 12207 40004 12256 40032
rect 12207 40001 12219 40004
rect 12161 39995 12219 40001
rect 11992 39964 12020 39995
rect 12250 39992 12256 40004
rect 12308 39992 12314 40044
rect 12618 40032 12624 40044
rect 12579 40004 12624 40032
rect 12618 39992 12624 40004
rect 12676 39992 12682 40044
rect 12802 40032 12808 40044
rect 12763 40004 12808 40032
rect 12802 39992 12808 40004
rect 12860 39992 12866 40044
rect 13740 40041 13768 40072
rect 14185 40103 14243 40109
rect 14185 40069 14197 40103
rect 14231 40100 14243 40103
rect 15378 40100 15384 40112
rect 14231 40072 15384 40100
rect 14231 40069 14243 40072
rect 14185 40063 14243 40069
rect 15378 40060 15384 40072
rect 15436 40060 15442 40112
rect 16669 40103 16727 40109
rect 16669 40100 16681 40103
rect 15488 40072 16681 40100
rect 13725 40035 13783 40041
rect 13725 40001 13737 40035
rect 13771 40001 13783 40035
rect 13725 39995 13783 40001
rect 14369 40035 14427 40041
rect 14369 40001 14381 40035
rect 14415 40001 14427 40035
rect 14642 40032 14648 40044
rect 14603 40004 14648 40032
rect 14369 39995 14427 40001
rect 12342 39964 12348 39976
rect 11992 39936 12348 39964
rect 12342 39924 12348 39936
rect 12400 39924 12406 39976
rect 13081 39967 13139 39973
rect 13081 39933 13093 39967
rect 13127 39964 13139 39967
rect 13814 39964 13820 39976
rect 13127 39936 13820 39964
rect 13127 39933 13139 39936
rect 13081 39927 13139 39933
rect 13814 39924 13820 39936
rect 13872 39924 13878 39976
rect 12526 39896 12532 39908
rect 11716 39868 12532 39896
rect 12526 39856 12532 39868
rect 12584 39896 12590 39908
rect 13541 39899 13599 39905
rect 13541 39896 13553 39899
rect 12584 39868 13553 39896
rect 12584 39856 12590 39868
rect 13541 39865 13553 39868
rect 13587 39865 13599 39899
rect 14384 39896 14412 39995
rect 14642 39992 14648 40004
rect 14700 39992 14706 40044
rect 14829 40035 14887 40041
rect 14829 40001 14841 40035
rect 14875 40001 14887 40035
rect 15286 40032 15292 40044
rect 15247 40004 15292 40032
rect 14829 39995 14887 40001
rect 14844 39964 14872 39995
rect 15286 39992 15292 40004
rect 15344 39992 15350 40044
rect 15488 40041 15516 40072
rect 16669 40069 16681 40072
rect 16715 40069 16727 40103
rect 16669 40063 16727 40069
rect 17218 40060 17224 40112
rect 17276 40100 17282 40112
rect 17972 40100 18000 40140
rect 18230 40128 18236 40180
rect 18288 40168 18294 40180
rect 19705 40171 19763 40177
rect 19705 40168 19717 40171
rect 18288 40140 19717 40168
rect 18288 40128 18294 40140
rect 19705 40137 19717 40140
rect 19751 40137 19763 40171
rect 19705 40131 19763 40137
rect 22833 40171 22891 40177
rect 22833 40137 22845 40171
rect 22879 40168 22891 40171
rect 23474 40168 23480 40180
rect 22879 40140 23480 40168
rect 22879 40137 22891 40140
rect 22833 40131 22891 40137
rect 23474 40128 23480 40140
rect 23532 40128 23538 40180
rect 26234 40168 26240 40180
rect 25700 40140 26240 40168
rect 17276 40072 17356 40100
rect 17276 40060 17282 40072
rect 15473 40035 15531 40041
rect 15473 40001 15485 40035
rect 15519 40001 15531 40035
rect 15473 39995 15531 40001
rect 16574 39992 16580 40044
rect 16632 40032 16638 40044
rect 16853 40035 16911 40041
rect 16853 40032 16865 40035
rect 16632 40004 16865 40032
rect 16632 39992 16638 40004
rect 16853 40001 16865 40004
rect 16899 40001 16911 40035
rect 17126 40032 17132 40044
rect 17087 40004 17132 40032
rect 16853 39995 16911 40001
rect 17126 39992 17132 40004
rect 17184 39992 17190 40044
rect 17328 40041 17356 40072
rect 17972 40072 19932 40100
rect 17972 40041 18000 40072
rect 17313 40035 17371 40041
rect 17313 40001 17325 40035
rect 17359 40001 17371 40035
rect 17313 39995 17371 40001
rect 17957 40035 18015 40041
rect 17957 40001 17969 40035
rect 18003 40001 18015 40035
rect 17957 39995 18015 40001
rect 18506 39992 18512 40044
rect 18564 40032 18570 40044
rect 19904 40041 19932 40072
rect 22186 40060 22192 40112
rect 22244 40100 22250 40112
rect 22244 40072 23336 40100
rect 22244 40060 22250 40072
rect 23308 40044 23336 40072
rect 24578 40060 24584 40112
rect 24636 40100 24642 40112
rect 25409 40103 25467 40109
rect 25409 40100 25421 40103
rect 24636 40072 25421 40100
rect 24636 40060 24642 40072
rect 25409 40069 25421 40072
rect 25455 40069 25467 40103
rect 25700 40100 25728 40140
rect 26234 40128 26240 40140
rect 26292 40168 26298 40180
rect 26789 40171 26847 40177
rect 26789 40168 26801 40171
rect 26292 40140 26801 40168
rect 26292 40128 26298 40140
rect 26789 40137 26801 40140
rect 26835 40168 26847 40171
rect 26878 40168 26884 40180
rect 26835 40140 26884 40168
rect 26835 40137 26847 40140
rect 26789 40131 26847 40137
rect 26878 40128 26884 40140
rect 26936 40128 26942 40180
rect 26973 40171 27031 40177
rect 26973 40137 26985 40171
rect 27019 40168 27031 40171
rect 27154 40168 27160 40180
rect 27019 40140 27160 40168
rect 27019 40137 27031 40140
rect 26973 40131 27031 40137
rect 27154 40128 27160 40140
rect 27212 40128 27218 40180
rect 28074 40168 28080 40180
rect 28035 40140 28080 40168
rect 28074 40128 28080 40140
rect 28132 40128 28138 40180
rect 28626 40128 28632 40180
rect 28684 40168 28690 40180
rect 29181 40171 29239 40177
rect 29181 40168 29193 40171
rect 28684 40140 29193 40168
rect 28684 40128 28690 40140
rect 29181 40137 29193 40140
rect 29227 40137 29239 40171
rect 29181 40131 29239 40137
rect 26694 40100 26700 40112
rect 25409 40063 25467 40069
rect 25608 40072 25728 40100
rect 25884 40072 26700 40100
rect 18693 40035 18751 40041
rect 18693 40032 18705 40035
rect 18564 40004 18705 40032
rect 18564 39992 18570 40004
rect 18693 40001 18705 40004
rect 18739 40001 18751 40035
rect 18693 39995 18751 40001
rect 19889 40035 19947 40041
rect 19889 40001 19901 40035
rect 19935 40001 19947 40035
rect 21818 40032 21824 40044
rect 21779 40004 21824 40032
rect 19889 39995 19947 40001
rect 21818 39992 21824 40004
rect 21876 39992 21882 40044
rect 22005 40035 22063 40041
rect 22005 40001 22017 40035
rect 22051 40032 22063 40035
rect 22830 40032 22836 40044
rect 22051 40004 22836 40032
rect 22051 40001 22063 40004
rect 22005 39995 22063 40001
rect 22830 39992 22836 40004
rect 22888 39992 22894 40044
rect 23014 40032 23020 40044
rect 22975 40004 23020 40032
rect 23014 39992 23020 40004
rect 23072 39992 23078 40044
rect 23290 40032 23296 40044
rect 23203 40004 23296 40032
rect 23290 39992 23296 40004
rect 23348 39992 23354 40044
rect 23477 40035 23535 40041
rect 23477 40001 23489 40035
rect 23523 40032 23535 40035
rect 23842 40032 23848 40044
rect 23523 40004 23848 40032
rect 23523 40001 23535 40004
rect 23477 39995 23535 40001
rect 23842 39992 23848 40004
rect 23900 39992 23906 40044
rect 25608 40041 25636 40072
rect 25884 40041 25912 40072
rect 26694 40060 26700 40072
rect 26752 40100 26758 40112
rect 27798 40100 27804 40112
rect 26752 40072 27804 40100
rect 26752 40060 26758 40072
rect 25593 40035 25651 40041
rect 25593 40001 25605 40035
rect 25639 40001 25651 40035
rect 25593 39995 25651 40001
rect 25869 40035 25927 40041
rect 25869 40001 25881 40035
rect 25915 40001 25927 40035
rect 25869 39995 25927 40001
rect 25958 39992 25964 40044
rect 26016 40032 26022 40044
rect 27448 40041 27476 40072
rect 27798 40060 27804 40072
rect 27856 40100 27862 40112
rect 30285 40103 30343 40109
rect 27856 40072 28580 40100
rect 27856 40060 27862 40072
rect 26053 40035 26111 40041
rect 26053 40032 26065 40035
rect 26016 40004 26065 40032
rect 26016 39992 26022 40004
rect 26053 40001 26065 40004
rect 26099 40001 26111 40035
rect 26053 39995 26111 40001
rect 26789 40035 26847 40041
rect 26789 40001 26801 40035
rect 26835 40032 26847 40035
rect 27157 40035 27215 40041
rect 27157 40032 27169 40035
rect 26835 40004 27169 40032
rect 26835 40001 26847 40004
rect 26789 39995 26847 40001
rect 27157 40001 27169 40004
rect 27203 40001 27215 40035
rect 27157 39995 27215 40001
rect 27433 40035 27491 40041
rect 27433 40001 27445 40035
rect 27479 40001 27491 40035
rect 27433 39995 27491 40001
rect 27617 40035 27675 40041
rect 27617 40001 27629 40035
rect 27663 40032 27675 40035
rect 27706 40032 27712 40044
rect 27663 40004 27712 40032
rect 27663 40001 27675 40004
rect 27617 39995 27675 40001
rect 15194 39964 15200 39976
rect 14844 39936 15200 39964
rect 15194 39924 15200 39936
rect 15252 39964 15258 39976
rect 15749 39967 15807 39973
rect 15749 39964 15761 39967
rect 15252 39936 15761 39964
rect 15252 39924 15258 39936
rect 15749 39933 15761 39936
rect 15795 39933 15807 39967
rect 15749 39927 15807 39933
rect 16206 39924 16212 39976
rect 16264 39964 16270 39976
rect 18414 39964 18420 39976
rect 16264 39936 17908 39964
rect 18375 39936 18420 39964
rect 16264 39924 16270 39936
rect 14734 39896 14740 39908
rect 14384 39868 14740 39896
rect 13541 39859 13599 39865
rect 14734 39856 14740 39868
rect 14792 39896 14798 39908
rect 17773 39899 17831 39905
rect 17773 39896 17785 39899
rect 14792 39868 17785 39896
rect 14792 39856 14798 39868
rect 17773 39865 17785 39868
rect 17819 39865 17831 39899
rect 17880 39896 17908 39936
rect 18414 39924 18420 39936
rect 18472 39964 18478 39976
rect 19702 39964 19708 39976
rect 18472 39936 19708 39964
rect 18472 39924 18478 39936
rect 19702 39924 19708 39936
rect 19760 39964 19766 39976
rect 20349 39967 20407 39973
rect 20349 39964 20361 39967
rect 19760 39936 20361 39964
rect 19760 39924 19766 39936
rect 20349 39933 20361 39936
rect 20395 39933 20407 39967
rect 20349 39927 20407 39933
rect 20625 39967 20683 39973
rect 20625 39933 20637 39967
rect 20671 39964 20683 39967
rect 22186 39964 22192 39976
rect 20671 39936 22192 39964
rect 20671 39933 20683 39936
rect 20625 39927 20683 39933
rect 22186 39924 22192 39936
rect 22244 39924 22250 39976
rect 22281 39967 22339 39973
rect 22281 39933 22293 39967
rect 22327 39964 22339 39967
rect 22922 39964 22928 39976
rect 22327 39936 22928 39964
rect 22327 39933 22339 39936
rect 22281 39927 22339 39933
rect 22922 39924 22928 39936
rect 22980 39924 22986 39976
rect 23658 39924 23664 39976
rect 23716 39964 23722 39976
rect 24121 39967 24179 39973
rect 24121 39964 24133 39967
rect 23716 39936 24133 39964
rect 23716 39924 23722 39936
rect 24121 39933 24133 39936
rect 24167 39933 24179 39967
rect 24121 39927 24179 39933
rect 24397 39967 24455 39973
rect 24397 39933 24409 39967
rect 24443 39964 24455 39967
rect 27172 39964 27200 39995
rect 27706 39992 27712 40004
rect 27764 39992 27770 40044
rect 28552 40041 28580 40072
rect 30285 40069 30297 40103
rect 30331 40100 30343 40103
rect 30650 40100 30656 40112
rect 30331 40072 30656 40100
rect 30331 40069 30343 40072
rect 30285 40063 30343 40069
rect 30650 40060 30656 40072
rect 30708 40060 30714 40112
rect 28261 40035 28319 40041
rect 28261 40001 28273 40035
rect 28307 40001 28319 40035
rect 28261 39995 28319 40001
rect 28537 40035 28595 40041
rect 28537 40001 28549 40035
rect 28583 40001 28595 40035
rect 28718 40032 28724 40044
rect 28679 40004 28724 40032
rect 28537 39995 28595 40001
rect 28276 39964 28304 39995
rect 28718 39992 28724 40004
rect 28776 40032 28782 40044
rect 28902 40032 28908 40044
rect 28776 40004 28908 40032
rect 28776 39992 28782 40004
rect 28902 39992 28908 40004
rect 28960 39992 28966 40044
rect 29365 40035 29423 40041
rect 29365 40001 29377 40035
rect 29411 40001 29423 40035
rect 29638 40032 29644 40044
rect 29599 40004 29644 40032
rect 29365 39995 29423 40001
rect 29380 39964 29408 39995
rect 29638 39992 29644 40004
rect 29696 39992 29702 40044
rect 29822 40032 29828 40044
rect 29783 40004 29828 40032
rect 29822 39992 29828 40004
rect 29880 39992 29886 40044
rect 30466 40032 30472 40044
rect 30427 40004 30472 40032
rect 30466 39992 30472 40004
rect 30524 39992 30530 40044
rect 30745 40035 30803 40041
rect 30745 40032 30757 40035
rect 30576 40004 30757 40032
rect 29454 39964 29460 39976
rect 24443 39936 27108 39964
rect 27172 39936 28304 39964
rect 29367 39936 29460 39964
rect 24443 39933 24455 39936
rect 24397 39927 24455 39933
rect 24854 39896 24860 39908
rect 17880 39868 24860 39896
rect 17773 39859 17831 39865
rect 24854 39856 24860 39868
rect 24912 39856 24918 39908
rect 27080 39896 27108 39936
rect 29454 39924 29460 39936
rect 29512 39964 29518 39976
rect 30484 39964 30512 39992
rect 29512 39936 30512 39964
rect 29512 39924 29518 39936
rect 28258 39896 28264 39908
rect 27080 39868 28264 39896
rect 28258 39856 28264 39868
rect 28316 39896 28322 39908
rect 28810 39896 28816 39908
rect 28316 39868 28816 39896
rect 28316 39856 28322 39868
rect 28810 39856 28816 39868
rect 28868 39856 28874 39908
rect 29638 39856 29644 39908
rect 29696 39896 29702 39908
rect 30576 39896 30604 40004
rect 30745 40001 30757 40004
rect 30791 40001 30803 40035
rect 30745 39995 30803 40001
rect 30929 40035 30987 40041
rect 30929 40001 30941 40035
rect 30975 40032 30987 40035
rect 31294 40032 31300 40044
rect 30975 40004 31300 40032
rect 30975 40001 30987 40004
rect 30929 39995 30987 40001
rect 31294 39992 31300 40004
rect 31352 39992 31358 40044
rect 29696 39868 30604 39896
rect 29696 39856 29702 39868
rect 2777 39831 2835 39837
rect 2777 39797 2789 39831
rect 2823 39828 2835 39831
rect 2866 39828 2872 39840
rect 2823 39800 2872 39828
rect 2823 39797 2835 39800
rect 2777 39791 2835 39797
rect 2866 39788 2872 39800
rect 2924 39828 2930 39840
rect 3786 39828 3792 39840
rect 2924 39800 3792 39828
rect 2924 39788 2930 39800
rect 3786 39788 3792 39800
rect 3844 39788 3850 39840
rect 5902 39788 5908 39840
rect 5960 39828 5966 39840
rect 7101 39831 7159 39837
rect 7101 39828 7113 39831
rect 5960 39800 7113 39828
rect 5960 39788 5966 39800
rect 7101 39797 7113 39800
rect 7147 39797 7159 39831
rect 7101 39791 7159 39797
rect 7190 39788 7196 39840
rect 7248 39828 7254 39840
rect 9030 39828 9036 39840
rect 7248 39800 9036 39828
rect 7248 39788 7254 39800
rect 9030 39788 9036 39800
rect 9088 39788 9094 39840
rect 10321 39831 10379 39837
rect 10321 39797 10333 39831
rect 10367 39828 10379 39831
rect 10778 39828 10784 39840
rect 10367 39800 10784 39828
rect 10367 39797 10379 39800
rect 10321 39791 10379 39797
rect 10778 39788 10784 39800
rect 10836 39788 10842 39840
rect 12618 39788 12624 39840
rect 12676 39828 12682 39840
rect 12894 39828 12900 39840
rect 12676 39800 12900 39828
rect 12676 39788 12682 39800
rect 12894 39788 12900 39800
rect 12952 39828 12958 39840
rect 12989 39831 13047 39837
rect 12989 39828 13001 39831
rect 12952 39800 13001 39828
rect 12952 39788 12958 39800
rect 12989 39797 13001 39800
rect 13035 39797 13047 39831
rect 15654 39828 15660 39840
rect 15615 39800 15660 39828
rect 12989 39791 13047 39797
rect 15654 39788 15660 39800
rect 15712 39788 15718 39840
rect 22189 39831 22247 39837
rect 22189 39797 22201 39831
rect 22235 39828 22247 39831
rect 22462 39828 22468 39840
rect 22235 39800 22468 39828
rect 22235 39797 22247 39800
rect 22189 39791 22247 39797
rect 22462 39788 22468 39800
rect 22520 39828 22526 39840
rect 23566 39828 23572 39840
rect 22520 39800 23572 39828
rect 22520 39788 22526 39800
rect 23566 39788 23572 39800
rect 23624 39788 23630 39840
rect 1104 39738 32016 39760
rect 1104 39686 2136 39738
rect 2188 39686 12440 39738
rect 12492 39686 22744 39738
rect 22796 39686 32016 39738
rect 1104 39664 32016 39686
rect 2590 39624 2596 39636
rect 2551 39596 2596 39624
rect 2590 39584 2596 39596
rect 2648 39584 2654 39636
rect 4249 39627 4307 39633
rect 4249 39593 4261 39627
rect 4295 39624 4307 39627
rect 7190 39624 7196 39636
rect 4295 39596 7196 39624
rect 4295 39593 4307 39596
rect 4249 39587 4307 39593
rect 7190 39584 7196 39596
rect 7248 39584 7254 39636
rect 7745 39627 7803 39633
rect 7745 39593 7757 39627
rect 7791 39624 7803 39627
rect 8386 39624 8392 39636
rect 7791 39596 8392 39624
rect 7791 39593 7803 39596
rect 7745 39587 7803 39593
rect 8386 39584 8392 39596
rect 8444 39584 8450 39636
rect 12253 39627 12311 39633
rect 12253 39593 12265 39627
rect 12299 39624 12311 39627
rect 12618 39624 12624 39636
rect 12299 39596 12624 39624
rect 12299 39593 12311 39596
rect 12253 39587 12311 39593
rect 12618 39584 12624 39596
rect 12676 39584 12682 39636
rect 16758 39624 16764 39636
rect 16719 39596 16764 39624
rect 16758 39584 16764 39596
rect 16816 39584 16822 39636
rect 18049 39627 18107 39633
rect 18049 39593 18061 39627
rect 18095 39624 18107 39627
rect 18138 39624 18144 39636
rect 18095 39596 18144 39624
rect 18095 39593 18107 39596
rect 18049 39587 18107 39593
rect 18138 39584 18144 39596
rect 18196 39584 18202 39636
rect 22830 39624 22836 39636
rect 22791 39596 22836 39624
rect 22830 39584 22836 39596
rect 22888 39584 22894 39636
rect 24397 39627 24455 39633
rect 24397 39593 24409 39627
rect 24443 39624 24455 39627
rect 24486 39624 24492 39636
rect 24443 39596 24492 39624
rect 24443 39593 24455 39596
rect 24397 39587 24455 39593
rect 24486 39584 24492 39596
rect 24544 39584 24550 39636
rect 7285 39559 7343 39565
rect 7285 39525 7297 39559
rect 7331 39556 7343 39559
rect 12066 39556 12072 39568
rect 7331 39528 12072 39556
rect 7331 39525 7343 39528
rect 7285 39519 7343 39525
rect 12066 39516 12072 39528
rect 12124 39516 12130 39568
rect 15654 39516 15660 39568
rect 15712 39556 15718 39568
rect 15749 39559 15807 39565
rect 15749 39556 15761 39559
rect 15712 39528 15761 39556
rect 15712 39516 15718 39528
rect 15749 39525 15761 39528
rect 15795 39556 15807 39559
rect 17129 39559 17187 39565
rect 17129 39556 17141 39559
rect 15795 39528 17141 39556
rect 15795 39525 15807 39528
rect 15749 39519 15807 39525
rect 17129 39525 17141 39528
rect 17175 39525 17187 39559
rect 17129 39519 17187 39525
rect 23566 39516 23572 39568
rect 23624 39556 23630 39568
rect 24765 39559 24823 39565
rect 24765 39556 24777 39559
rect 23624 39528 24777 39556
rect 23624 39516 23630 39528
rect 24765 39525 24777 39528
rect 24811 39525 24823 39559
rect 24765 39519 24823 39525
rect 25958 39516 25964 39568
rect 26016 39556 26022 39568
rect 28721 39559 28779 39565
rect 28721 39556 28733 39559
rect 26016 39528 28733 39556
rect 26016 39516 26022 39528
rect 28721 39525 28733 39528
rect 28767 39525 28779 39559
rect 28721 39519 28779 39525
rect 2682 39448 2688 39500
rect 2740 39488 2746 39500
rect 2961 39491 3019 39497
rect 2961 39488 2973 39491
rect 2740 39460 2973 39488
rect 2740 39448 2746 39460
rect 2961 39457 2973 39460
rect 3007 39457 3019 39491
rect 2961 39451 3019 39457
rect 3234 39448 3240 39500
rect 3292 39488 3298 39500
rect 4614 39488 4620 39500
rect 3292 39460 4476 39488
rect 4575 39460 4620 39488
rect 3292 39448 3298 39460
rect 2774 39380 2780 39432
rect 2832 39420 2838 39432
rect 3050 39420 3056 39432
rect 2832 39392 2877 39420
rect 3011 39392 3056 39420
rect 2832 39380 2838 39392
rect 3050 39380 3056 39392
rect 3108 39380 3114 39432
rect 4246 39420 4252 39432
rect 4159 39392 4252 39420
rect 4246 39380 4252 39392
rect 4304 39420 4310 39432
rect 4341 39423 4399 39429
rect 4341 39420 4353 39423
rect 4304 39392 4353 39420
rect 4304 39380 4310 39392
rect 4341 39389 4353 39392
rect 4387 39389 4399 39423
rect 4448 39420 4476 39460
rect 4614 39448 4620 39460
rect 4672 39448 4678 39500
rect 9217 39491 9275 39497
rect 9217 39488 9229 39491
rect 6012 39460 7144 39488
rect 6012 39429 6040 39460
rect 7116 39432 7144 39460
rect 8312 39460 9229 39488
rect 8312 39432 8340 39460
rect 9217 39457 9229 39460
rect 9263 39457 9275 39491
rect 12805 39491 12863 39497
rect 12805 39488 12817 39491
rect 9217 39451 9275 39457
rect 12084 39460 12817 39488
rect 5629 39423 5687 39429
rect 5629 39420 5641 39423
rect 4448 39392 5641 39420
rect 4341 39383 4399 39389
rect 5629 39389 5641 39392
rect 5675 39389 5687 39423
rect 5905 39423 5963 39429
rect 5905 39420 5917 39423
rect 5629 39383 5687 39389
rect 5736 39392 5917 39420
rect 1765 39355 1823 39361
rect 1765 39352 1777 39355
rect 768 39324 1777 39352
rect 768 39148 796 39324
rect 1765 39321 1777 39324
rect 1811 39321 1823 39355
rect 1765 39315 1823 39321
rect 3786 39312 3792 39364
rect 3844 39352 3850 39364
rect 5736 39352 5764 39392
rect 5905 39389 5917 39392
rect 5951 39389 5963 39423
rect 5905 39383 5963 39389
rect 5997 39423 6055 39429
rect 5997 39389 6009 39423
rect 6043 39389 6055 39423
rect 5997 39383 6055 39389
rect 6733 39423 6791 39429
rect 6733 39389 6745 39423
rect 6779 39389 6791 39423
rect 7098 39420 7104 39432
rect 7059 39392 7104 39420
rect 6733 39383 6791 39389
rect 3844 39324 5764 39352
rect 5813 39355 5871 39361
rect 3844 39312 3850 39324
rect 5813 39321 5825 39355
rect 5859 39352 5871 39355
rect 6638 39352 6644 39364
rect 5859 39324 6644 39352
rect 5859 39321 5871 39324
rect 5813 39315 5871 39321
rect 6638 39312 6644 39324
rect 6696 39312 6702 39364
rect 1854 39284 1860 39296
rect 1815 39256 1860 39284
rect 1854 39244 1860 39256
rect 1912 39244 1918 39296
rect 5442 39244 5448 39296
rect 5500 39284 5506 39296
rect 6181 39287 6239 39293
rect 6181 39284 6193 39287
rect 5500 39256 6193 39284
rect 5500 39244 5506 39256
rect 6181 39253 6193 39256
rect 6227 39253 6239 39287
rect 6748 39284 6776 39383
rect 7098 39380 7104 39392
rect 7156 39380 7162 39432
rect 7926 39420 7932 39432
rect 7887 39392 7932 39420
rect 7926 39380 7932 39392
rect 7984 39380 7990 39432
rect 8205 39423 8263 39429
rect 8205 39389 8217 39423
rect 8251 39420 8263 39423
rect 8294 39420 8300 39432
rect 8251 39392 8300 39420
rect 8251 39389 8263 39392
rect 8205 39383 8263 39389
rect 8294 39380 8300 39392
rect 8352 39380 8358 39432
rect 8389 39423 8447 39429
rect 8389 39389 8401 39423
rect 8435 39420 8447 39423
rect 8478 39420 8484 39432
rect 8435 39392 8484 39420
rect 8435 39389 8447 39392
rect 8389 39383 8447 39389
rect 6822 39312 6828 39364
rect 6880 39352 6886 39364
rect 6917 39355 6975 39361
rect 6917 39352 6929 39355
rect 6880 39324 6929 39352
rect 6880 39312 6886 39324
rect 6917 39321 6929 39324
rect 6963 39321 6975 39355
rect 6917 39315 6975 39321
rect 7009 39355 7067 39361
rect 7009 39321 7021 39355
rect 7055 39352 7067 39355
rect 8404 39352 8432 39383
rect 8478 39380 8484 39392
rect 8536 39380 8542 39432
rect 8941 39423 8999 39429
rect 8941 39389 8953 39423
rect 8987 39420 8999 39423
rect 9030 39420 9036 39432
rect 8987 39392 9036 39420
rect 8987 39389 8999 39392
rect 8941 39383 8999 39389
rect 9030 39380 9036 39392
rect 9088 39380 9094 39432
rect 10318 39380 10324 39432
rect 10376 39420 10382 39432
rect 10597 39423 10655 39429
rect 10597 39420 10609 39423
rect 10376 39392 10609 39420
rect 10376 39380 10382 39392
rect 10597 39389 10609 39392
rect 10643 39389 10655 39423
rect 10778 39420 10784 39432
rect 10739 39392 10784 39420
rect 10597 39383 10655 39389
rect 10778 39380 10784 39392
rect 10836 39380 10842 39432
rect 12084 39429 12112 39460
rect 12805 39457 12817 39460
rect 12851 39457 12863 39491
rect 14369 39491 14427 39497
rect 14369 39488 14381 39491
rect 12805 39451 12863 39457
rect 13280 39460 14381 39488
rect 10873 39423 10931 39429
rect 10873 39389 10885 39423
rect 10919 39389 10931 39423
rect 10873 39383 10931 39389
rect 12069 39423 12127 39429
rect 12069 39389 12081 39423
rect 12115 39389 12127 39423
rect 12069 39383 12127 39389
rect 12345 39423 12403 39429
rect 12345 39389 12357 39423
rect 12391 39389 12403 39423
rect 12345 39383 12403 39389
rect 12989 39423 13047 39429
rect 12989 39389 13001 39423
rect 13035 39420 13047 39423
rect 13078 39420 13084 39432
rect 13035 39392 13084 39420
rect 13035 39389 13047 39392
rect 12989 39383 13047 39389
rect 7055 39324 8432 39352
rect 10888 39352 10916 39383
rect 12250 39352 12256 39364
rect 10888 39324 12256 39352
rect 7055 39321 7067 39324
rect 7009 39315 7067 39321
rect 12250 39312 12256 39324
rect 12308 39312 12314 39364
rect 9674 39284 9680 39296
rect 6748 39256 9680 39284
rect 6181 39247 6239 39253
rect 9674 39244 9680 39256
rect 9732 39244 9738 39296
rect 9766 39244 9772 39296
rect 9824 39284 9830 39296
rect 10413 39287 10471 39293
rect 10413 39284 10425 39287
rect 9824 39256 10425 39284
rect 9824 39244 9830 39256
rect 10413 39253 10425 39256
rect 10459 39253 10471 39287
rect 10413 39247 10471 39253
rect 11885 39287 11943 39293
rect 11885 39253 11897 39287
rect 11931 39284 11943 39287
rect 11974 39284 11980 39296
rect 11931 39256 11980 39284
rect 11931 39253 11943 39256
rect 11885 39247 11943 39253
rect 11974 39244 11980 39256
rect 12032 39244 12038 39296
rect 12360 39284 12388 39383
rect 13078 39380 13084 39392
rect 13136 39380 13142 39432
rect 13280 39429 13308 39460
rect 14369 39457 14381 39460
rect 14415 39488 14427 39491
rect 14642 39488 14648 39500
rect 14415 39460 14648 39488
rect 14415 39457 14427 39460
rect 14369 39451 14427 39457
rect 14642 39448 14648 39460
rect 14700 39448 14706 39500
rect 17221 39491 17279 39497
rect 17221 39457 17233 39491
rect 17267 39488 17279 39491
rect 17310 39488 17316 39500
rect 17267 39460 17316 39488
rect 17267 39457 17279 39460
rect 17221 39451 17279 39457
rect 17310 39448 17316 39460
rect 17368 39488 17374 39500
rect 17494 39488 17500 39500
rect 17368 39460 17500 39488
rect 17368 39448 17374 39460
rect 17494 39448 17500 39460
rect 17552 39448 17558 39500
rect 18414 39488 18420 39500
rect 18064 39460 18420 39488
rect 13265 39423 13323 39429
rect 13265 39389 13277 39423
rect 13311 39389 13323 39423
rect 13265 39383 13323 39389
rect 13449 39423 13507 39429
rect 13449 39389 13461 39423
rect 13495 39420 13507 39423
rect 13814 39420 13820 39432
rect 13495 39392 13820 39420
rect 13495 39389 13507 39392
rect 13449 39383 13507 39389
rect 13814 39380 13820 39392
rect 13872 39380 13878 39432
rect 14093 39423 14151 39429
rect 14093 39389 14105 39423
rect 14139 39389 14151 39423
rect 14093 39383 14151 39389
rect 14108 39352 14136 39383
rect 15378 39380 15384 39432
rect 15436 39420 15442 39432
rect 15565 39423 15623 39429
rect 15565 39420 15577 39423
rect 15436 39392 15577 39420
rect 15436 39380 15442 39392
rect 15565 39389 15577 39392
rect 15611 39389 15623 39423
rect 15565 39383 15623 39389
rect 15838 39380 15844 39432
rect 15896 39420 15902 39432
rect 16942 39420 16948 39432
rect 15896 39392 15941 39420
rect 16903 39392 16948 39420
rect 15896 39380 15902 39392
rect 16942 39380 16948 39392
rect 17000 39380 17006 39432
rect 18064 39420 18092 39460
rect 18414 39448 18420 39460
rect 18472 39448 18478 39500
rect 19613 39491 19671 39497
rect 19613 39457 19625 39491
rect 19659 39488 19671 39491
rect 20990 39488 20996 39500
rect 19659 39460 20996 39488
rect 19659 39457 19671 39460
rect 19613 39451 19671 39457
rect 20990 39448 20996 39460
rect 21048 39448 21054 39500
rect 23842 39448 23848 39500
rect 23900 39488 23906 39500
rect 24670 39488 24676 39500
rect 23900 39460 24676 39488
rect 23900 39448 23906 39460
rect 24670 39448 24676 39460
rect 24728 39488 24734 39500
rect 24857 39491 24915 39497
rect 24857 39488 24869 39491
rect 24728 39460 24869 39488
rect 24728 39448 24734 39460
rect 24857 39457 24869 39460
rect 24903 39457 24915 39491
rect 24857 39451 24915 39457
rect 27617 39491 27675 39497
rect 27617 39457 27629 39491
rect 27663 39488 27675 39491
rect 27798 39488 27804 39500
rect 27663 39460 27804 39488
rect 27663 39457 27675 39460
rect 27617 39451 27675 39457
rect 27798 39448 27804 39460
rect 27856 39448 27862 39500
rect 29546 39448 29552 39500
rect 29604 39488 29610 39500
rect 29917 39491 29975 39497
rect 29917 39488 29929 39491
rect 29604 39460 29929 39488
rect 29604 39448 29610 39460
rect 29917 39457 29929 39460
rect 29963 39457 29975 39491
rect 29917 39451 29975 39457
rect 18230 39420 18236 39432
rect 17328 39392 18092 39420
rect 18191 39392 18236 39420
rect 17328 39352 17356 39392
rect 18230 39380 18236 39392
rect 18288 39380 18294 39432
rect 18506 39420 18512 39432
rect 18467 39392 18512 39420
rect 18506 39380 18512 39392
rect 18564 39380 18570 39432
rect 18693 39423 18751 39429
rect 18693 39389 18705 39423
rect 18739 39389 18751 39423
rect 19426 39420 19432 39432
rect 19387 39392 19432 39420
rect 18693 39383 18751 39389
rect 14108 39324 17356 39352
rect 17402 39312 17408 39364
rect 17460 39352 17466 39364
rect 18708 39352 18736 39383
rect 19426 39380 19432 39392
rect 19484 39380 19490 39432
rect 19705 39423 19763 39429
rect 19705 39389 19717 39423
rect 19751 39420 19763 39423
rect 21174 39420 21180 39432
rect 19751 39392 21180 39420
rect 19751 39389 19763 39392
rect 19705 39383 19763 39389
rect 21174 39380 21180 39392
rect 21232 39380 21238 39432
rect 23014 39420 23020 39432
rect 22975 39392 23020 39420
rect 23014 39380 23020 39392
rect 23072 39380 23078 39432
rect 23290 39420 23296 39432
rect 23251 39392 23296 39420
rect 23290 39380 23296 39392
rect 23348 39380 23354 39432
rect 23477 39423 23535 39429
rect 23477 39389 23489 39423
rect 23523 39420 23535 39423
rect 24302 39420 24308 39432
rect 23523 39392 24308 39420
rect 23523 39389 23535 39392
rect 23477 39383 23535 39389
rect 24302 39380 24308 39392
rect 24360 39380 24366 39432
rect 24578 39420 24584 39432
rect 24539 39392 24584 39420
rect 24578 39380 24584 39392
rect 24636 39380 24642 39432
rect 25866 39420 25872 39432
rect 25827 39392 25872 39420
rect 25866 39380 25872 39392
rect 25924 39380 25930 39432
rect 26234 39420 26240 39432
rect 26195 39392 26240 39420
rect 26234 39380 26240 39392
rect 26292 39380 26298 39432
rect 27341 39423 27399 39429
rect 27341 39389 27353 39423
rect 27387 39389 27399 39423
rect 28626 39420 28632 39432
rect 28587 39392 28632 39420
rect 27341 39383 27399 39389
rect 19518 39352 19524 39364
rect 17460 39324 19524 39352
rect 17460 39312 17466 39324
rect 19518 39312 19524 39324
rect 19576 39312 19582 39364
rect 20622 39352 20628 39364
rect 20583 39324 20628 39352
rect 20622 39312 20628 39324
rect 20680 39312 20686 39364
rect 25590 39312 25596 39364
rect 25648 39352 25654 39364
rect 26053 39355 26111 39361
rect 26053 39352 26065 39355
rect 25648 39324 26065 39352
rect 25648 39312 25654 39324
rect 26053 39321 26065 39324
rect 26099 39321 26111 39355
rect 26053 39315 26111 39321
rect 26145 39355 26203 39361
rect 26145 39321 26157 39355
rect 26191 39352 26203 39355
rect 26326 39352 26332 39364
rect 26191 39324 26332 39352
rect 26191 39321 26203 39324
rect 26145 39315 26203 39321
rect 26326 39312 26332 39324
rect 26384 39312 26390 39364
rect 27356 39352 27384 39383
rect 28626 39380 28632 39392
rect 28684 39380 28690 39432
rect 29178 39352 29184 39364
rect 27356 39324 29184 39352
rect 29178 39312 29184 39324
rect 29236 39312 29242 39364
rect 30184 39355 30242 39361
rect 30184 39321 30196 39355
rect 30230 39352 30242 39355
rect 30466 39352 30472 39364
rect 30230 39324 30472 39352
rect 30230 39321 30242 39324
rect 30184 39315 30242 39321
rect 30466 39312 30472 39324
rect 30524 39312 30530 39364
rect 13354 39284 13360 39296
rect 12360 39256 13360 39284
rect 13354 39244 13360 39256
rect 13412 39244 13418 39296
rect 15378 39284 15384 39296
rect 15339 39256 15384 39284
rect 15378 39244 15384 39256
rect 15436 39244 15442 39296
rect 19245 39287 19303 39293
rect 19245 39253 19257 39287
rect 19291 39284 19303 39287
rect 20070 39284 20076 39296
rect 19291 39256 20076 39284
rect 19291 39253 19303 39256
rect 19245 39247 19303 39253
rect 20070 39244 20076 39256
rect 20128 39244 20134 39296
rect 21634 39244 21640 39296
rect 21692 39284 21698 39296
rect 21913 39287 21971 39293
rect 21913 39284 21925 39287
rect 21692 39256 21925 39284
rect 21692 39244 21698 39256
rect 21913 39253 21925 39256
rect 21959 39253 21971 39287
rect 21913 39247 21971 39253
rect 26421 39287 26479 39293
rect 26421 39253 26433 39287
rect 26467 39284 26479 39287
rect 27154 39284 27160 39296
rect 26467 39256 27160 39284
rect 26467 39253 26479 39256
rect 26421 39247 26479 39253
rect 27154 39244 27160 39256
rect 27212 39244 27218 39296
rect 31294 39284 31300 39296
rect 31255 39256 31300 39284
rect 31294 39244 31300 39256
rect 31352 39244 31358 39296
rect 1104 39194 32016 39216
rect 768 39120 888 39148
rect 1104 39142 7288 39194
rect 7340 39142 17592 39194
rect 17644 39142 27896 39194
rect 27948 39142 32016 39194
rect 1104 39120 32016 39142
rect 0 39012 800 39026
rect 860 39012 888 39120
rect 2774 39040 2780 39092
rect 2832 39080 2838 39092
rect 3145 39083 3203 39089
rect 3145 39080 3157 39083
rect 2832 39052 3157 39080
rect 2832 39040 2838 39052
rect 3145 39049 3157 39052
rect 3191 39049 3203 39083
rect 3510 39080 3516 39092
rect 3145 39043 3203 39049
rect 3344 39052 3516 39080
rect 0 38984 888 39012
rect 0 38970 800 38984
rect 2406 38944 2412 38956
rect 2367 38916 2412 38944
rect 2406 38904 2412 38916
rect 2464 38904 2470 38956
rect 3344 38953 3372 39052
rect 3510 39040 3516 39052
rect 3568 39080 3574 39092
rect 6365 39083 6423 39089
rect 6365 39080 6377 39083
rect 3568 39052 6377 39080
rect 3568 39040 3574 39052
rect 6365 39049 6377 39052
rect 6411 39049 6423 39083
rect 8110 39080 8116 39092
rect 6365 39043 6423 39049
rect 6932 39052 8116 39080
rect 4614 39012 4620 39024
rect 3620 38984 4620 39012
rect 3620 38953 3648 38984
rect 4614 38972 4620 38984
rect 4672 38972 4678 39024
rect 5902 39012 5908 39024
rect 5092 38984 5908 39012
rect 3329 38947 3387 38953
rect 3329 38913 3341 38947
rect 3375 38913 3387 38947
rect 3329 38907 3387 38913
rect 3605 38947 3663 38953
rect 3605 38913 3617 38947
rect 3651 38913 3663 38947
rect 3786 38944 3792 38956
rect 3747 38916 3792 38944
rect 3605 38907 3663 38913
rect 3786 38904 3792 38916
rect 3844 38904 3850 38956
rect 5092 38953 5120 38984
rect 5902 38972 5908 38984
rect 5960 38972 5966 39024
rect 4433 38947 4491 38953
rect 4433 38913 4445 38947
rect 4479 38913 4491 38947
rect 4433 38907 4491 38913
rect 5077 38947 5135 38953
rect 5077 38913 5089 38947
rect 5123 38913 5135 38947
rect 5077 38907 5135 38913
rect 2685 38879 2743 38885
rect 2685 38845 2697 38879
rect 2731 38876 2743 38879
rect 2774 38876 2780 38888
rect 2731 38848 2780 38876
rect 2731 38845 2743 38848
rect 2685 38839 2743 38845
rect 2774 38836 2780 38848
rect 2832 38836 2838 38888
rect 4448 38876 4476 38907
rect 5166 38904 5172 38956
rect 5224 38944 5230 38956
rect 5350 38944 5356 38956
rect 5224 38916 5269 38944
rect 5311 38916 5356 38944
rect 5224 38904 5230 38916
rect 5350 38904 5356 38916
rect 5408 38904 5414 38956
rect 5626 38953 5632 38956
rect 5445 38947 5503 38953
rect 5445 38913 5457 38947
rect 5491 38913 5503 38947
rect 5445 38907 5503 38913
rect 5583 38947 5632 38953
rect 5583 38913 5595 38947
rect 5629 38913 5632 38947
rect 5583 38907 5632 38913
rect 4448 38848 5212 38876
rect 4617 38811 4675 38817
rect 4617 38808 4629 38811
rect 3068 38780 4629 38808
rect 2222 38740 2228 38752
rect 2183 38712 2228 38740
rect 2222 38700 2228 38712
rect 2280 38700 2286 38752
rect 2593 38743 2651 38749
rect 2593 38709 2605 38743
rect 2639 38740 2651 38743
rect 2682 38740 2688 38752
rect 2639 38712 2688 38740
rect 2639 38709 2651 38712
rect 2593 38703 2651 38709
rect 2682 38700 2688 38712
rect 2740 38740 2746 38752
rect 3068 38740 3096 38780
rect 4617 38777 4629 38780
rect 4663 38777 4675 38811
rect 5184 38808 5212 38848
rect 5258 38836 5264 38888
rect 5316 38876 5322 38888
rect 5460 38876 5488 38907
rect 5626 38904 5632 38907
rect 5684 38904 5690 38956
rect 6546 38944 6552 38956
rect 6507 38916 6552 38944
rect 6546 38904 6552 38916
rect 6604 38904 6610 38956
rect 5316 38848 5488 38876
rect 5316 38836 5322 38848
rect 6932 38808 6960 39052
rect 8110 39040 8116 39052
rect 8168 39040 8174 39092
rect 8202 39040 8208 39092
rect 8260 39080 8266 39092
rect 10318 39080 10324 39092
rect 8260 39052 9720 39080
rect 10279 39052 10324 39080
rect 8260 39040 8266 39052
rect 7009 39015 7067 39021
rect 7009 38981 7021 39015
rect 7055 39012 7067 39015
rect 7055 38984 9444 39012
rect 7055 38981 7067 38984
rect 7009 38975 7067 38981
rect 7193 38947 7251 38953
rect 7193 38913 7205 38947
rect 7239 38913 7251 38947
rect 7193 38907 7251 38913
rect 7469 38947 7527 38953
rect 7469 38913 7481 38947
rect 7515 38913 7527 38947
rect 7650 38944 7656 38956
rect 7611 38916 7656 38944
rect 7469 38907 7527 38913
rect 5184 38780 6960 38808
rect 7208 38808 7236 38907
rect 7484 38876 7512 38907
rect 7650 38904 7656 38916
rect 7708 38904 7714 38956
rect 7926 38904 7932 38956
rect 7984 38944 7990 38956
rect 8297 38947 8355 38953
rect 8297 38944 8309 38947
rect 7984 38916 8309 38944
rect 7984 38904 7990 38916
rect 8297 38913 8309 38916
rect 8343 38913 8355 38947
rect 8297 38907 8355 38913
rect 8573 38947 8631 38953
rect 8573 38913 8585 38947
rect 8619 38913 8631 38947
rect 8754 38944 8760 38956
rect 8715 38916 8760 38944
rect 8573 38907 8631 38913
rect 8386 38876 8392 38888
rect 7484 38848 8392 38876
rect 8386 38836 8392 38848
rect 8444 38876 8450 38888
rect 8588 38876 8616 38907
rect 8754 38904 8760 38916
rect 8812 38904 8818 38956
rect 9416 38953 9444 38984
rect 9692 38953 9720 39052
rect 10318 39040 10324 39052
rect 10376 39040 10382 39092
rect 10778 39040 10784 39092
rect 10836 39080 10842 39092
rect 16025 39083 16083 39089
rect 16025 39080 16037 39083
rect 10836 39052 16037 39080
rect 10836 39040 10842 39052
rect 16025 39049 16037 39052
rect 16071 39049 16083 39083
rect 16025 39043 16083 39049
rect 19426 39040 19432 39092
rect 19484 39080 19490 39092
rect 21821 39083 21879 39089
rect 21821 39080 21833 39083
rect 19484 39052 21833 39080
rect 19484 39040 19490 39052
rect 21821 39049 21833 39052
rect 21867 39049 21879 39083
rect 22833 39083 22891 39089
rect 22833 39080 22845 39083
rect 21821 39043 21879 39049
rect 22066 39052 22845 39080
rect 12526 39012 12532 39024
rect 10520 38984 12532 39012
rect 10520 38953 10548 38984
rect 12526 38972 12532 38984
rect 12584 38972 12590 39024
rect 14268 39015 14326 39021
rect 14268 38981 14280 39015
rect 14314 39012 14326 39015
rect 15378 39012 15384 39024
rect 14314 38984 15384 39012
rect 14314 38981 14326 38984
rect 14268 38975 14326 38981
rect 15378 38972 15384 38984
rect 15436 38972 15442 39024
rect 17497 39015 17555 39021
rect 17497 39012 17509 39015
rect 15488 38984 17509 39012
rect 9401 38947 9459 38953
rect 9401 38913 9413 38947
rect 9447 38913 9459 38947
rect 9401 38907 9459 38913
rect 9677 38947 9735 38953
rect 9677 38913 9689 38947
rect 9723 38913 9735 38947
rect 9677 38907 9735 38913
rect 10505 38947 10563 38953
rect 10505 38913 10517 38947
rect 10551 38913 10563 38947
rect 10505 38907 10563 38913
rect 10781 38947 10839 38953
rect 10781 38913 10793 38947
rect 10827 38913 10839 38947
rect 10962 38944 10968 38956
rect 10923 38916 10968 38944
rect 10781 38907 10839 38913
rect 10796 38876 10824 38907
rect 10962 38904 10968 38916
rect 11020 38904 11026 38956
rect 11882 38944 11888 38956
rect 11843 38916 11888 38944
rect 11882 38904 11888 38916
rect 11940 38904 11946 38956
rect 11974 38904 11980 38956
rect 12032 38944 12038 38956
rect 12141 38947 12199 38953
rect 12141 38944 12153 38947
rect 12032 38916 12153 38944
rect 12032 38904 12038 38916
rect 12141 38913 12153 38916
rect 12187 38913 12199 38947
rect 12141 38907 12199 38913
rect 15286 38904 15292 38956
rect 15344 38944 15350 38956
rect 15488 38944 15516 38984
rect 17497 38981 17509 38984
rect 17543 38981 17555 39015
rect 17497 38975 17555 38981
rect 17589 39015 17647 39021
rect 17589 38981 17601 39015
rect 17635 39012 17647 39015
rect 18046 39012 18052 39024
rect 17635 38984 18052 39012
rect 17635 38981 17647 38984
rect 17589 38975 17647 38981
rect 18046 38972 18052 38984
rect 18104 38972 18110 39024
rect 21542 39012 21548 39024
rect 18156 38984 20208 39012
rect 15930 38944 15936 38956
rect 15344 38916 15516 38944
rect 15891 38916 15936 38944
rect 15344 38904 15350 38916
rect 15930 38904 15936 38916
rect 15988 38904 15994 38956
rect 17218 38944 17224 38956
rect 17179 38916 17224 38944
rect 17218 38904 17224 38916
rect 17276 38904 17282 38956
rect 17313 38947 17371 38953
rect 17313 38913 17325 38947
rect 17359 38944 17371 38947
rect 17402 38944 17408 38956
rect 17359 38916 17408 38944
rect 17359 38913 17371 38916
rect 17313 38907 17371 38913
rect 17402 38904 17408 38916
rect 17460 38904 17466 38956
rect 17681 38947 17739 38953
rect 17681 38913 17693 38947
rect 17727 38913 17739 38947
rect 17681 38907 17739 38913
rect 11790 38876 11796 38888
rect 8444 38848 8616 38876
rect 8864 38848 10732 38876
rect 10796 38848 11796 38876
rect 8444 38836 8450 38848
rect 7926 38808 7932 38820
rect 7208 38780 7932 38808
rect 4617 38771 4675 38777
rect 7926 38768 7932 38780
rect 7984 38768 7990 38820
rect 8202 38768 8208 38820
rect 8260 38808 8266 38820
rect 8864 38808 8892 38848
rect 8260 38780 8892 38808
rect 8260 38768 8266 38780
rect 8938 38768 8944 38820
rect 8996 38808 9002 38820
rect 9585 38811 9643 38817
rect 9585 38808 9597 38811
rect 8996 38780 9597 38808
rect 8996 38768 9002 38780
rect 9585 38777 9597 38780
rect 9631 38777 9643 38811
rect 9585 38771 9643 38777
rect 5718 38740 5724 38752
rect 2740 38712 3096 38740
rect 5679 38712 5724 38740
rect 2740 38700 2746 38712
rect 5718 38700 5724 38712
rect 5776 38700 5782 38752
rect 7742 38700 7748 38752
rect 7800 38740 7806 38752
rect 8113 38743 8171 38749
rect 8113 38740 8125 38743
rect 7800 38712 8125 38740
rect 7800 38700 7806 38712
rect 8113 38709 8125 38712
rect 8159 38709 8171 38743
rect 8113 38703 8171 38709
rect 8294 38700 8300 38752
rect 8352 38740 8358 38752
rect 9217 38743 9275 38749
rect 9217 38740 9229 38743
rect 8352 38712 9229 38740
rect 8352 38700 8358 38712
rect 9217 38709 9229 38712
rect 9263 38709 9275 38743
rect 10704 38740 10732 38848
rect 11790 38836 11796 38848
rect 11848 38836 11854 38888
rect 13998 38876 14004 38888
rect 13959 38848 14004 38876
rect 13998 38836 14004 38848
rect 14056 38836 14062 38888
rect 15562 38836 15568 38888
rect 15620 38876 15626 38888
rect 17696 38876 17724 38907
rect 15620 38848 17724 38876
rect 15620 38836 15626 38848
rect 15194 38768 15200 38820
rect 15252 38808 15258 38820
rect 15381 38811 15439 38817
rect 15381 38808 15393 38811
rect 15252 38780 15393 38808
rect 15252 38768 15258 38780
rect 15381 38777 15393 38780
rect 15427 38777 15439 38811
rect 15381 38771 15439 38777
rect 17402 38768 17408 38820
rect 17460 38808 17466 38820
rect 18156 38808 18184 38984
rect 18233 38947 18291 38953
rect 18233 38913 18245 38947
rect 18279 38944 18291 38947
rect 18322 38944 18328 38956
rect 18279 38916 18328 38944
rect 18279 38913 18291 38916
rect 18233 38907 18291 38913
rect 18322 38904 18328 38916
rect 18380 38904 18386 38956
rect 18500 38947 18558 38953
rect 18500 38913 18512 38947
rect 18546 38944 18558 38947
rect 18874 38944 18880 38956
rect 18546 38916 18880 38944
rect 18546 38913 18558 38916
rect 18500 38907 18558 38913
rect 18874 38904 18880 38916
rect 18932 38904 18938 38956
rect 20180 38953 20208 38984
rect 20456 38984 21548 39012
rect 20456 38956 20484 38984
rect 21542 38972 21548 38984
rect 21600 39012 21606 39024
rect 22066 39012 22094 39052
rect 22833 39049 22845 39052
rect 22879 39049 22891 39083
rect 22833 39043 22891 39049
rect 23290 39040 23296 39092
rect 23348 39080 23354 39092
rect 27157 39083 27215 39089
rect 23348 39052 24072 39080
rect 23348 39040 23354 39052
rect 21600 38984 22094 39012
rect 22204 38984 22692 39012
rect 21600 38972 21606 38984
rect 20165 38947 20223 38953
rect 20165 38913 20177 38947
rect 20211 38913 20223 38947
rect 20438 38944 20444 38956
rect 20399 38916 20444 38944
rect 20165 38907 20223 38913
rect 20438 38904 20444 38916
rect 20496 38904 20502 38956
rect 22005 38947 22063 38953
rect 22005 38913 22017 38947
rect 22051 38944 22063 38947
rect 22204 38944 22232 38984
rect 22051 38916 22232 38944
rect 22051 38913 22063 38916
rect 22005 38907 22063 38913
rect 22278 38904 22284 38956
rect 22336 38944 22342 38956
rect 22465 38947 22523 38953
rect 22336 38916 22381 38944
rect 22336 38904 22342 38916
rect 22465 38913 22477 38947
rect 22511 38944 22523 38947
rect 22557 38947 22615 38953
rect 22557 38944 22569 38947
rect 22511 38916 22569 38944
rect 22511 38913 22523 38916
rect 22465 38907 22523 38913
rect 22557 38913 22569 38916
rect 22603 38913 22615 38947
rect 22664 38944 22692 38984
rect 22922 38972 22928 39024
rect 22980 39012 22986 39024
rect 22980 38984 23612 39012
rect 22980 38972 22986 38984
rect 23014 38944 23020 38956
rect 22664 38916 23020 38944
rect 22557 38907 22615 38913
rect 23014 38904 23020 38916
rect 23072 38944 23078 38956
rect 23109 38947 23167 38953
rect 23109 38944 23121 38947
rect 23072 38916 23121 38944
rect 23072 38904 23078 38916
rect 23109 38913 23121 38916
rect 23155 38913 23167 38947
rect 23382 38944 23388 38956
rect 23343 38916 23388 38944
rect 23109 38907 23167 38913
rect 23382 38904 23388 38916
rect 23440 38904 23446 38956
rect 23584 38953 23612 38984
rect 24044 38953 24072 39052
rect 27157 39049 27169 39083
rect 27203 39080 27215 39083
rect 28718 39080 28724 39092
rect 27203 39052 28724 39080
rect 27203 39049 27215 39052
rect 27157 39043 27215 39049
rect 28718 39040 28724 39052
rect 28776 39040 28782 39092
rect 30466 39080 30472 39092
rect 30427 39052 30472 39080
rect 30466 39040 30472 39052
rect 30524 39040 30530 39092
rect 25590 38972 25596 39024
rect 25648 39012 25654 39024
rect 27433 39015 27491 39021
rect 27433 39012 27445 39015
rect 25648 38984 27445 39012
rect 25648 38972 25654 38984
rect 27433 38981 27445 38984
rect 27479 38981 27491 39015
rect 27433 38975 27491 38981
rect 27525 39015 27583 39021
rect 27525 38981 27537 39015
rect 27571 39012 27583 39015
rect 31294 39012 31300 39024
rect 27571 38984 31300 39012
rect 27571 38981 27583 38984
rect 27525 38975 27583 38981
rect 31294 38972 31300 38984
rect 31352 38972 31358 39024
rect 32320 39012 33120 39026
rect 31726 38984 33120 39012
rect 23569 38947 23627 38953
rect 23569 38913 23581 38947
rect 23615 38913 23627 38947
rect 23569 38907 23627 38913
rect 24029 38947 24087 38953
rect 24029 38913 24041 38947
rect 24075 38913 24087 38947
rect 24029 38907 24087 38913
rect 24213 38947 24271 38953
rect 24213 38913 24225 38947
rect 24259 38944 24271 38947
rect 24578 38944 24584 38956
rect 24259 38916 24584 38944
rect 24259 38913 24271 38916
rect 24213 38907 24271 38913
rect 24578 38904 24584 38916
rect 24636 38904 24642 38956
rect 24673 38947 24731 38953
rect 24673 38913 24685 38947
rect 24719 38913 24731 38947
rect 24673 38907 24731 38913
rect 27157 38947 27215 38953
rect 27157 38913 27169 38947
rect 27203 38944 27215 38947
rect 27249 38947 27307 38953
rect 27249 38944 27261 38947
rect 27203 38916 27261 38944
rect 27203 38913 27215 38916
rect 27157 38907 27215 38913
rect 27249 38913 27261 38916
rect 27295 38913 27307 38947
rect 27614 38944 27620 38956
rect 27575 38916 27620 38944
rect 27249 38907 27307 38913
rect 20622 38836 20628 38888
rect 20680 38876 20686 38888
rect 24688 38876 24716 38907
rect 27614 38904 27620 38916
rect 27672 38904 27678 38956
rect 28442 38944 28448 38956
rect 28403 38916 28448 38944
rect 28442 38904 28448 38916
rect 28500 38904 28506 38956
rect 28629 38947 28687 38953
rect 28629 38913 28641 38947
rect 28675 38944 28687 38947
rect 28810 38944 28816 38956
rect 28675 38916 28816 38944
rect 28675 38913 28687 38916
rect 28629 38907 28687 38913
rect 28810 38904 28816 38916
rect 28868 38904 28874 38956
rect 30650 38944 30656 38956
rect 30611 38916 30656 38944
rect 30650 38904 30656 38916
rect 30708 38904 30714 38956
rect 30837 38947 30895 38953
rect 30837 38913 30849 38947
rect 30883 38944 30895 38947
rect 31018 38944 31024 38956
rect 30883 38916 31024 38944
rect 30883 38913 30895 38916
rect 30837 38907 30895 38913
rect 31018 38904 31024 38916
rect 31076 38904 31082 38956
rect 20680 38848 24716 38876
rect 20680 38836 20686 38848
rect 25866 38836 25872 38888
rect 25924 38876 25930 38888
rect 28721 38879 28779 38885
rect 28721 38876 28733 38879
rect 25924 38848 28733 38876
rect 25924 38836 25930 38848
rect 28721 38845 28733 38848
rect 28767 38845 28779 38879
rect 29178 38876 29184 38888
rect 29139 38848 29184 38876
rect 28721 38839 28779 38845
rect 29178 38836 29184 38848
rect 29236 38836 29242 38888
rect 29457 38879 29515 38885
rect 29457 38845 29469 38879
rect 29503 38876 29515 38879
rect 29638 38876 29644 38888
rect 29503 38848 29644 38876
rect 29503 38845 29515 38848
rect 29457 38839 29515 38845
rect 29638 38836 29644 38848
rect 29696 38876 29702 38888
rect 30006 38876 30012 38888
rect 29696 38848 30012 38876
rect 29696 38836 29702 38848
rect 30006 38836 30012 38848
rect 30064 38836 30070 38888
rect 30926 38876 30932 38888
rect 30887 38848 30932 38876
rect 30926 38836 30932 38848
rect 30984 38836 30990 38888
rect 17460 38780 18184 38808
rect 17460 38768 17466 38780
rect 20898 38768 20904 38820
rect 20956 38808 20962 38820
rect 21910 38808 21916 38820
rect 20956 38780 21916 38808
rect 20956 38768 20962 38780
rect 21910 38768 21916 38780
rect 21968 38808 21974 38820
rect 22557 38811 22615 38817
rect 22557 38808 22569 38811
rect 21968 38780 22569 38808
rect 21968 38768 21974 38780
rect 22557 38777 22569 38780
rect 22603 38777 22615 38811
rect 22557 38771 22615 38777
rect 22833 38811 22891 38817
rect 22833 38777 22845 38811
rect 22879 38808 22891 38811
rect 23658 38808 23664 38820
rect 22879 38780 23664 38808
rect 22879 38777 22891 38780
rect 22833 38771 22891 38777
rect 23658 38768 23664 38780
rect 23716 38768 23722 38820
rect 24762 38768 24768 38820
rect 24820 38808 24826 38820
rect 28261 38811 28319 38817
rect 28261 38808 28273 38811
rect 24820 38780 28273 38808
rect 24820 38768 24826 38780
rect 28261 38777 28273 38780
rect 28307 38777 28319 38811
rect 28261 38771 28319 38777
rect 28350 38768 28356 38820
rect 28408 38808 28414 38820
rect 31726 38808 31754 38984
rect 32320 38970 33120 38984
rect 28408 38780 31754 38808
rect 28408 38768 28414 38780
rect 11514 38740 11520 38752
rect 10704 38712 11520 38740
rect 9217 38703 9275 38709
rect 11514 38700 11520 38712
rect 11572 38740 11578 38752
rect 12158 38740 12164 38752
rect 11572 38712 12164 38740
rect 11572 38700 11578 38712
rect 12158 38700 12164 38712
rect 12216 38700 12222 38752
rect 13265 38743 13323 38749
rect 13265 38709 13277 38743
rect 13311 38740 13323 38743
rect 13814 38740 13820 38752
rect 13311 38712 13820 38740
rect 13311 38709 13323 38712
rect 13265 38703 13323 38709
rect 13814 38700 13820 38712
rect 13872 38740 13878 38752
rect 14642 38740 14648 38752
rect 13872 38712 14648 38740
rect 13872 38700 13878 38712
rect 14642 38700 14648 38712
rect 14700 38700 14706 38752
rect 16574 38700 16580 38752
rect 16632 38740 16638 38752
rect 17221 38743 17279 38749
rect 17221 38740 17233 38743
rect 16632 38712 17233 38740
rect 16632 38700 16638 38712
rect 17221 38709 17233 38712
rect 17267 38709 17279 38743
rect 17221 38703 17279 38709
rect 18506 38700 18512 38752
rect 18564 38740 18570 38752
rect 19613 38743 19671 38749
rect 19613 38740 19625 38743
rect 18564 38712 19625 38740
rect 18564 38700 18570 38712
rect 19613 38709 19625 38712
rect 19659 38709 19671 38743
rect 19613 38703 19671 38709
rect 22278 38700 22284 38752
rect 22336 38740 22342 38752
rect 22925 38743 22983 38749
rect 22925 38740 22937 38743
rect 22336 38712 22937 38740
rect 22336 38700 22342 38712
rect 22925 38709 22937 38712
rect 22971 38709 22983 38743
rect 22925 38703 22983 38709
rect 24029 38743 24087 38749
rect 24029 38709 24041 38743
rect 24075 38740 24087 38743
rect 24210 38740 24216 38752
rect 24075 38712 24216 38740
rect 24075 38709 24087 38712
rect 24029 38703 24087 38709
rect 24210 38700 24216 38712
rect 24268 38700 24274 38752
rect 25774 38700 25780 38752
rect 25832 38740 25838 38752
rect 25961 38743 26019 38749
rect 25961 38740 25973 38743
rect 25832 38712 25973 38740
rect 25832 38700 25838 38712
rect 25961 38709 25973 38712
rect 26007 38709 26019 38743
rect 27798 38740 27804 38752
rect 27759 38712 27804 38740
rect 25961 38703 26019 38709
rect 27798 38700 27804 38712
rect 27856 38700 27862 38752
rect 1104 38650 32016 38672
rect 1104 38598 2136 38650
rect 2188 38598 12440 38650
rect 12492 38598 22744 38650
rect 22796 38598 32016 38650
rect 1104 38576 32016 38598
rect 3050 38496 3056 38548
rect 3108 38536 3114 38548
rect 3237 38539 3295 38545
rect 3237 38536 3249 38539
rect 3108 38508 3249 38536
rect 3108 38496 3114 38508
rect 3237 38505 3249 38508
rect 3283 38505 3295 38539
rect 5442 38536 5448 38548
rect 5403 38508 5448 38536
rect 3237 38499 3295 38505
rect 3252 38400 3280 38499
rect 5442 38496 5448 38508
rect 5500 38496 5506 38548
rect 6546 38496 6552 38548
rect 6604 38536 6610 38548
rect 8297 38539 8355 38545
rect 8297 38536 8309 38539
rect 6604 38508 8309 38536
rect 6604 38496 6610 38508
rect 8297 38505 8309 38508
rect 8343 38505 8355 38539
rect 11882 38536 11888 38548
rect 11843 38508 11888 38536
rect 8297 38499 8355 38505
rect 11882 38496 11888 38508
rect 11940 38496 11946 38548
rect 12066 38496 12072 38548
rect 12124 38536 12130 38548
rect 14093 38539 14151 38545
rect 14093 38536 14105 38539
rect 12124 38508 14105 38536
rect 12124 38496 12130 38508
rect 14093 38505 14105 38508
rect 14139 38505 14151 38539
rect 14093 38499 14151 38505
rect 14274 38496 14280 38548
rect 14332 38536 14338 38548
rect 14332 38508 16988 38536
rect 14332 38496 14338 38508
rect 4430 38428 4436 38480
rect 4488 38428 4494 38480
rect 4522 38428 4528 38480
rect 4580 38468 4586 38480
rect 5350 38468 5356 38480
rect 4580 38440 5356 38468
rect 4580 38428 4586 38440
rect 5350 38428 5356 38440
rect 5408 38428 5414 38480
rect 7650 38468 7656 38480
rect 7611 38440 7656 38468
rect 7650 38428 7656 38440
rect 7708 38428 7714 38480
rect 8754 38428 8760 38480
rect 8812 38468 8818 38480
rect 9493 38471 9551 38477
rect 8812 38440 9260 38468
rect 8812 38428 8818 38440
rect 4448 38400 4476 38428
rect 5442 38400 5448 38412
rect 3252 38372 4384 38400
rect 4448 38372 5448 38400
rect 1394 38292 1400 38344
rect 1452 38332 1458 38344
rect 1857 38335 1915 38341
rect 1857 38332 1869 38335
rect 1452 38304 1869 38332
rect 1452 38292 1458 38304
rect 1857 38301 1869 38304
rect 1903 38301 1915 38335
rect 1857 38295 1915 38301
rect 2866 38292 2872 38344
rect 2924 38332 2930 38344
rect 4356 38341 4384 38372
rect 5442 38360 5448 38372
rect 5500 38400 5506 38412
rect 6273 38403 6331 38409
rect 6273 38400 6285 38403
rect 5500 38372 6285 38400
rect 5500 38360 5506 38372
rect 6273 38369 6285 38372
rect 6319 38369 6331 38403
rect 7668 38400 7696 38428
rect 8018 38400 8024 38412
rect 7668 38372 8024 38400
rect 6273 38363 6331 38369
rect 8018 38360 8024 38372
rect 8076 38400 8082 38412
rect 8076 38372 8984 38400
rect 8076 38360 8082 38372
rect 4065 38335 4123 38341
rect 4065 38332 4077 38335
rect 2924 38304 4077 38332
rect 2924 38292 2930 38304
rect 4065 38301 4077 38304
rect 4111 38301 4123 38335
rect 4065 38295 4123 38301
rect 4341 38335 4399 38341
rect 4341 38301 4353 38335
rect 4387 38301 4399 38335
rect 4341 38295 4399 38301
rect 4430 38292 4436 38344
rect 4488 38332 4494 38344
rect 5353 38335 5411 38341
rect 5353 38332 5365 38335
rect 4488 38304 4533 38332
rect 4632 38304 5365 38332
rect 4488 38292 4494 38304
rect 2124 38267 2182 38273
rect 2124 38233 2136 38267
rect 2170 38264 2182 38267
rect 2222 38264 2228 38276
rect 2170 38236 2228 38264
rect 2170 38233 2182 38236
rect 2124 38227 2182 38233
rect 2222 38224 2228 38236
rect 2280 38224 2286 38276
rect 4249 38267 4307 38273
rect 4249 38233 4261 38267
rect 4295 38264 4307 38267
rect 4522 38264 4528 38276
rect 4295 38236 4528 38264
rect 4295 38233 4307 38236
rect 4249 38227 4307 38233
rect 4522 38224 4528 38236
rect 4580 38224 4586 38276
rect 4632 38205 4660 38304
rect 5353 38301 5365 38304
rect 5399 38301 5411 38335
rect 5534 38332 5540 38344
rect 5495 38304 5540 38332
rect 5353 38295 5411 38301
rect 5534 38292 5540 38304
rect 5592 38292 5598 38344
rect 6540 38335 6598 38341
rect 6540 38301 6552 38335
rect 6586 38332 6598 38335
rect 8294 38332 8300 38344
rect 6586 38304 8300 38332
rect 6586 38301 6598 38304
rect 6540 38295 6598 38301
rect 8294 38292 8300 38304
rect 8352 38292 8358 38344
rect 8956 38341 8984 38372
rect 9232 38341 9260 38440
rect 9493 38437 9505 38471
rect 9539 38437 9551 38471
rect 9493 38431 9551 38437
rect 9508 38400 9536 38431
rect 11698 38428 11704 38480
rect 11756 38468 11762 38480
rect 11756 38440 13676 38468
rect 11756 38428 11762 38440
rect 13648 38400 13676 38440
rect 13998 38428 14004 38480
rect 14056 38468 14062 38480
rect 16301 38471 16359 38477
rect 16301 38468 16313 38471
rect 14056 38440 16313 38468
rect 14056 38428 14062 38440
rect 16301 38437 16313 38440
rect 16347 38437 16359 38471
rect 16301 38431 16359 38437
rect 16960 38400 16988 38508
rect 17218 38496 17224 38548
rect 17276 38536 17282 38548
rect 17773 38539 17831 38545
rect 17773 38536 17785 38539
rect 17276 38508 17785 38536
rect 17276 38496 17282 38508
rect 17773 38505 17785 38508
rect 17819 38505 17831 38539
rect 17773 38499 17831 38505
rect 18601 38539 18659 38545
rect 18601 38505 18613 38539
rect 18647 38536 18659 38539
rect 19058 38536 19064 38548
rect 18647 38508 19064 38536
rect 18647 38505 18659 38508
rect 18601 38499 18659 38505
rect 19058 38496 19064 38508
rect 19116 38496 19122 38548
rect 22922 38496 22928 38548
rect 22980 38536 22986 38548
rect 23017 38539 23075 38545
rect 23017 38536 23029 38539
rect 22980 38508 23029 38536
rect 22980 38496 22986 38508
rect 23017 38505 23029 38508
rect 23063 38505 23075 38539
rect 27614 38536 27620 38548
rect 23017 38499 23075 38505
rect 25148 38508 27620 38536
rect 17129 38471 17187 38477
rect 17129 38437 17141 38471
rect 17175 38468 17187 38471
rect 19334 38468 19340 38480
rect 17175 38440 19340 38468
rect 17175 38437 17187 38440
rect 17129 38431 17187 38437
rect 19334 38428 19340 38440
rect 19392 38428 19398 38480
rect 17034 38400 17040 38412
rect 9508 38372 13584 38400
rect 13648 38372 15148 38400
rect 16947 38372 17040 38400
rect 8941 38335 8999 38341
rect 8941 38301 8953 38335
rect 8987 38301 8999 38335
rect 8941 38295 8999 38301
rect 9217 38335 9275 38341
rect 9217 38301 9229 38335
rect 9263 38301 9275 38335
rect 9217 38295 9275 38301
rect 9306 38292 9312 38344
rect 9364 38342 9370 38344
rect 9364 38332 9444 38342
rect 10137 38335 10195 38341
rect 9364 38304 9457 38332
rect 9364 38292 9370 38304
rect 8202 38264 8208 38276
rect 8163 38236 8208 38264
rect 8202 38224 8208 38236
rect 8260 38224 8266 38276
rect 8386 38224 8392 38276
rect 8444 38264 8450 38276
rect 9125 38267 9183 38273
rect 9125 38264 9137 38267
rect 8444 38236 9137 38264
rect 8444 38224 8450 38236
rect 9125 38233 9137 38236
rect 9171 38233 9183 38267
rect 9416 38264 9444 38304
rect 10137 38301 10149 38335
rect 10183 38332 10195 38335
rect 12066 38332 12072 38344
rect 10183 38304 12072 38332
rect 10183 38301 10195 38304
rect 10137 38295 10195 38301
rect 12066 38292 12072 38304
rect 12124 38292 12130 38344
rect 12526 38292 12532 38344
rect 12584 38332 12590 38344
rect 12989 38335 13047 38341
rect 12989 38332 13001 38335
rect 12584 38304 13001 38332
rect 12584 38292 12590 38304
rect 12989 38301 13001 38304
rect 13035 38301 13047 38335
rect 12989 38295 13047 38301
rect 13078 38292 13084 38344
rect 13136 38332 13142 38344
rect 13265 38335 13323 38341
rect 13265 38332 13277 38335
rect 13136 38304 13277 38332
rect 13136 38292 13142 38304
rect 13265 38301 13277 38304
rect 13311 38301 13323 38335
rect 13265 38295 13323 38301
rect 13354 38292 13360 38344
rect 13412 38332 13418 38344
rect 13449 38335 13507 38341
rect 13449 38332 13461 38335
rect 13412 38304 13461 38332
rect 13412 38292 13418 38304
rect 13449 38301 13461 38304
rect 13495 38301 13507 38335
rect 13556 38332 13584 38372
rect 14093 38335 14151 38341
rect 14093 38332 14105 38335
rect 13556 38304 14105 38332
rect 13449 38295 13507 38301
rect 14093 38301 14105 38304
rect 14139 38301 14151 38335
rect 14093 38295 14151 38301
rect 14182 38292 14188 38344
rect 14240 38332 14246 38344
rect 14240 38304 14285 38332
rect 14240 38292 14246 38304
rect 10226 38264 10232 38276
rect 9416 38236 10232 38264
rect 9125 38227 9183 38233
rect 10226 38224 10232 38236
rect 10284 38224 10290 38276
rect 10594 38264 10600 38276
rect 10555 38236 10600 38264
rect 10594 38224 10600 38236
rect 10652 38264 10658 38276
rect 15013 38267 15071 38273
rect 15013 38264 15025 38267
rect 10652 38236 15025 38264
rect 10652 38224 10658 38236
rect 15013 38233 15025 38236
rect 15059 38233 15071 38267
rect 15120 38264 15148 38372
rect 17034 38360 17040 38372
rect 17092 38400 17098 38412
rect 17092 38372 17448 38400
rect 17092 38360 17098 38372
rect 17420 38341 17448 38372
rect 18506 38360 18512 38412
rect 18564 38400 18570 38412
rect 18693 38403 18751 38409
rect 18693 38400 18705 38403
rect 18564 38372 18705 38400
rect 18564 38360 18570 38372
rect 18693 38369 18705 38372
rect 18739 38369 18751 38403
rect 18693 38363 18751 38369
rect 23750 38360 23756 38412
rect 23808 38400 23814 38412
rect 23808 38372 24532 38400
rect 23808 38360 23814 38372
rect 17129 38335 17187 38341
rect 17129 38301 17141 38335
rect 17175 38332 17187 38335
rect 17221 38335 17279 38341
rect 17221 38332 17233 38335
rect 17175 38304 17233 38332
rect 17175 38301 17187 38304
rect 17129 38295 17187 38301
rect 17221 38301 17233 38304
rect 17267 38301 17279 38335
rect 17221 38295 17279 38301
rect 17405 38335 17463 38341
rect 17405 38301 17417 38335
rect 17451 38301 17463 38335
rect 17405 38295 17463 38301
rect 17494 38292 17500 38344
rect 17552 38332 17558 38344
rect 17678 38341 17684 38344
rect 17635 38335 17684 38341
rect 17552 38304 17597 38332
rect 17552 38292 17558 38304
rect 17635 38301 17647 38335
rect 17681 38301 17684 38335
rect 17635 38295 17684 38301
rect 17678 38292 17684 38295
rect 17736 38292 17742 38344
rect 17770 38292 17776 38344
rect 17828 38332 17834 38344
rect 18417 38335 18475 38341
rect 18417 38332 18429 38335
rect 17828 38304 18429 38332
rect 17828 38292 17834 38304
rect 18417 38301 18429 38304
rect 18463 38301 18475 38335
rect 18417 38295 18475 38301
rect 19610 38292 19616 38344
rect 19668 38332 19674 38344
rect 19797 38335 19855 38341
rect 19797 38332 19809 38335
rect 19668 38304 19809 38332
rect 19668 38292 19674 38304
rect 19797 38301 19809 38304
rect 19843 38332 19855 38335
rect 21634 38332 21640 38344
rect 19843 38304 21640 38332
rect 19843 38301 19855 38304
rect 19797 38295 19855 38301
rect 21634 38292 21640 38304
rect 21692 38292 21698 38344
rect 23658 38332 23664 38344
rect 23619 38304 23664 38332
rect 23658 38292 23664 38304
rect 23716 38292 23722 38344
rect 24394 38332 24400 38344
rect 24355 38304 24400 38332
rect 24394 38292 24400 38304
rect 24452 38292 24458 38344
rect 24504 38341 24532 38372
rect 24670 38360 24676 38412
rect 24728 38360 24734 38412
rect 24490 38335 24548 38341
rect 24490 38301 24502 38335
rect 24536 38301 24548 38335
rect 24688 38332 24716 38360
rect 24765 38335 24823 38341
rect 24765 38332 24777 38335
rect 24688 38304 24777 38332
rect 24490 38295 24548 38301
rect 24765 38301 24777 38304
rect 24811 38301 24823 38335
rect 24765 38295 24823 38301
rect 24854 38292 24860 38344
rect 24912 38341 24918 38344
rect 24912 38332 24920 38341
rect 25148 38332 25176 38508
rect 26234 38468 26240 38480
rect 24912 38304 25176 38332
rect 25240 38440 26240 38468
rect 24912 38295 24920 38304
rect 24912 38292 24918 38295
rect 20070 38273 20076 38276
rect 20064 38264 20076 38273
rect 15120 38236 19748 38264
rect 20031 38236 20076 38264
rect 15013 38227 15071 38233
rect 4617 38199 4675 38205
rect 4617 38165 4629 38199
rect 4663 38165 4675 38199
rect 4617 38159 4675 38165
rect 5721 38199 5779 38205
rect 5721 38165 5733 38199
rect 5767 38196 5779 38199
rect 8110 38196 8116 38208
rect 5767 38168 8116 38196
rect 5767 38165 5779 38168
rect 5721 38159 5779 38165
rect 8110 38156 8116 38168
rect 8168 38156 8174 38208
rect 9950 38196 9956 38208
rect 9911 38168 9956 38196
rect 9950 38156 9956 38168
rect 10008 38156 10014 38208
rect 11790 38156 11796 38208
rect 11848 38196 11854 38208
rect 12805 38199 12863 38205
rect 12805 38196 12817 38199
rect 11848 38168 12817 38196
rect 11848 38156 11854 38168
rect 12805 38165 12817 38168
rect 12851 38165 12863 38199
rect 12805 38159 12863 38165
rect 13814 38156 13820 38208
rect 13872 38196 13878 38208
rect 14461 38199 14519 38205
rect 14461 38196 14473 38199
rect 13872 38168 14473 38196
rect 13872 38156 13878 38168
rect 14461 38165 14473 38168
rect 14507 38165 14519 38199
rect 18230 38196 18236 38208
rect 18191 38168 18236 38196
rect 14461 38159 14519 38165
rect 18230 38156 18236 38168
rect 18288 38156 18294 38208
rect 19720 38196 19748 38236
rect 20064 38227 20076 38236
rect 20070 38224 20076 38227
rect 20128 38224 20134 38276
rect 20990 38224 20996 38276
rect 21048 38264 21054 38276
rect 21904 38267 21962 38273
rect 21048 38236 21312 38264
rect 21048 38224 21054 38236
rect 20898 38196 20904 38208
rect 19720 38168 20904 38196
rect 20898 38156 20904 38168
rect 20956 38196 20962 38208
rect 21177 38199 21235 38205
rect 21177 38196 21189 38199
rect 20956 38168 21189 38196
rect 20956 38156 20962 38168
rect 21177 38165 21189 38168
rect 21223 38165 21235 38199
rect 21284 38196 21312 38236
rect 21904 38233 21916 38267
rect 21950 38264 21962 38267
rect 22094 38264 22100 38276
rect 21950 38236 22100 38264
rect 21950 38233 21962 38236
rect 21904 38227 21962 38233
rect 22094 38224 22100 38236
rect 22152 38224 22158 38276
rect 24673 38267 24731 38273
rect 22940 38236 23152 38264
rect 22940 38196 22968 38236
rect 21284 38168 22968 38196
rect 23124 38196 23152 38236
rect 24673 38233 24685 38267
rect 24719 38264 24731 38267
rect 25240 38264 25268 38440
rect 26234 38428 26240 38440
rect 26292 38428 26298 38480
rect 26605 38403 26663 38409
rect 26605 38400 26617 38403
rect 25700 38372 26617 38400
rect 25700 38341 25728 38372
rect 26605 38369 26617 38372
rect 26651 38369 26663 38403
rect 26605 38363 26663 38369
rect 25685 38335 25743 38341
rect 25685 38301 25697 38335
rect 25731 38301 25743 38335
rect 26142 38332 26148 38344
rect 26103 38304 26148 38332
rect 25685 38295 25743 38301
rect 26142 38292 26148 38304
rect 26200 38292 26206 38344
rect 26804 38341 26832 38508
rect 27614 38496 27620 38508
rect 27672 38496 27678 38548
rect 27798 38496 27804 38548
rect 27856 38536 27862 38548
rect 28629 38539 28687 38545
rect 28629 38536 28641 38539
rect 27856 38508 28641 38536
rect 27856 38496 27862 38508
rect 28629 38505 28641 38508
rect 28675 38505 28687 38539
rect 28629 38499 28687 38505
rect 29549 38539 29607 38545
rect 29549 38505 29561 38539
rect 29595 38536 29607 38539
rect 29730 38536 29736 38548
rect 29595 38508 29736 38536
rect 29595 38505 29607 38508
rect 29549 38499 29607 38505
rect 29730 38496 29736 38508
rect 29788 38496 29794 38548
rect 31018 38536 31024 38548
rect 30979 38508 31024 38536
rect 31018 38496 31024 38508
rect 31076 38496 31082 38548
rect 27706 38468 27712 38480
rect 26896 38440 27712 38468
rect 26896 38341 26924 38440
rect 27706 38428 27712 38440
rect 27764 38428 27770 38480
rect 28169 38471 28227 38477
rect 28169 38437 28181 38471
rect 28215 38468 28227 38471
rect 28537 38471 28595 38477
rect 28537 38468 28549 38471
rect 28215 38440 28549 38468
rect 28215 38437 28227 38440
rect 28169 38431 28227 38437
rect 28537 38437 28549 38440
rect 28583 38437 28595 38471
rect 28537 38431 28595 38437
rect 28997 38471 29055 38477
rect 28997 38437 29009 38471
rect 29043 38437 29055 38471
rect 28997 38431 29055 38437
rect 29012 38400 29040 38431
rect 30926 38400 30932 38412
rect 27540 38372 29040 38400
rect 30208 38372 30932 38400
rect 26789 38335 26847 38341
rect 26789 38301 26801 38335
rect 26835 38301 26847 38335
rect 26789 38295 26847 38301
rect 26881 38335 26939 38341
rect 26881 38301 26893 38335
rect 26927 38301 26939 38335
rect 27062 38332 27068 38344
rect 27023 38304 27068 38332
rect 26881 38295 26939 38301
rect 27062 38292 27068 38304
rect 27120 38292 27126 38344
rect 27154 38292 27160 38344
rect 27212 38332 27218 38344
rect 27212 38304 27257 38332
rect 27212 38292 27218 38304
rect 24719 38236 25268 38264
rect 24719 38233 24731 38236
rect 24673 38227 24731 38233
rect 25314 38224 25320 38276
rect 25372 38264 25378 38276
rect 25777 38267 25835 38273
rect 25777 38264 25789 38267
rect 25372 38236 25789 38264
rect 25372 38224 25378 38236
rect 25777 38233 25789 38236
rect 25823 38233 25835 38267
rect 25777 38227 25835 38233
rect 25866 38224 25872 38276
rect 25924 38264 25930 38276
rect 26007 38267 26065 38273
rect 25924 38236 25969 38264
rect 25924 38224 25930 38236
rect 26007 38233 26019 38267
rect 26053 38264 26065 38267
rect 27540 38264 27568 38372
rect 27617 38335 27675 38341
rect 27617 38301 27629 38335
rect 27663 38301 27675 38335
rect 27798 38332 27804 38344
rect 27759 38304 27804 38332
rect 27617 38295 27675 38301
rect 26053 38236 27568 38264
rect 27632 38264 27660 38295
rect 27798 38292 27804 38304
rect 27856 38292 27862 38344
rect 27982 38332 27988 38344
rect 27943 38304 27988 38332
rect 27982 38292 27988 38304
rect 28040 38292 28046 38344
rect 28537 38335 28595 38341
rect 28537 38301 28549 38335
rect 28583 38332 28595 38335
rect 28629 38335 28687 38341
rect 28629 38332 28641 38335
rect 28583 38304 28641 38332
rect 28583 38301 28595 38304
rect 28537 38295 28595 38301
rect 28629 38301 28641 38304
rect 28675 38301 28687 38335
rect 28629 38295 28687 38301
rect 28718 38292 28724 38344
rect 28776 38332 28782 38344
rect 28776 38304 28821 38332
rect 28776 38292 28782 38304
rect 29454 38292 29460 38344
rect 29512 38332 29518 38344
rect 29730 38332 29736 38344
rect 29512 38304 29736 38332
rect 29512 38292 29518 38304
rect 29730 38292 29736 38304
rect 29788 38292 29794 38344
rect 30006 38332 30012 38344
rect 29967 38304 30012 38332
rect 30006 38292 30012 38304
rect 30064 38292 30070 38344
rect 30208 38341 30236 38372
rect 30926 38360 30932 38372
rect 30984 38360 30990 38412
rect 31113 38403 31171 38409
rect 31113 38369 31125 38403
rect 31159 38400 31171 38403
rect 31294 38400 31300 38412
rect 31159 38372 31300 38400
rect 31159 38369 31171 38372
rect 31113 38363 31171 38369
rect 31294 38360 31300 38372
rect 31352 38360 31358 38412
rect 30193 38335 30251 38341
rect 30193 38332 30205 38335
rect 30116 38304 30205 38332
rect 27893 38267 27951 38273
rect 27632 38236 27844 38264
rect 26053 38233 26065 38236
rect 26007 38227 26065 38233
rect 23753 38199 23811 38205
rect 23753 38196 23765 38199
rect 23124 38168 23765 38196
rect 21177 38159 21235 38165
rect 23753 38165 23765 38168
rect 23799 38165 23811 38199
rect 23753 38159 23811 38165
rect 24486 38156 24492 38208
rect 24544 38196 24550 38208
rect 25041 38199 25099 38205
rect 25041 38196 25053 38199
rect 24544 38168 25053 38196
rect 24544 38156 24550 38168
rect 25041 38165 25053 38168
rect 25087 38165 25099 38199
rect 25041 38159 25099 38165
rect 25501 38199 25559 38205
rect 25501 38165 25513 38199
rect 25547 38196 25559 38199
rect 25682 38196 25688 38208
rect 25547 38168 25688 38196
rect 25547 38165 25559 38168
rect 25501 38159 25559 38165
rect 25682 38156 25688 38168
rect 25740 38156 25746 38208
rect 26326 38156 26332 38208
rect 26384 38196 26390 38208
rect 27430 38196 27436 38208
rect 26384 38168 27436 38196
rect 26384 38156 26390 38168
rect 27430 38156 27436 38168
rect 27488 38156 27494 38208
rect 27816 38196 27844 38236
rect 27893 38233 27905 38267
rect 27939 38264 27951 38267
rect 29822 38264 29828 38276
rect 27939 38236 29828 38264
rect 27939 38233 27951 38236
rect 27893 38227 27951 38233
rect 29822 38224 29828 38236
rect 29880 38224 29886 38276
rect 30116 38196 30144 38304
rect 30193 38301 30205 38304
rect 30239 38301 30251 38335
rect 30193 38295 30251 38301
rect 30282 38292 30288 38344
rect 30340 38332 30346 38344
rect 30837 38335 30895 38341
rect 30837 38332 30849 38335
rect 30340 38304 30849 38332
rect 30340 38292 30346 38304
rect 30837 38301 30849 38304
rect 30883 38301 30895 38335
rect 30837 38295 30895 38301
rect 30650 38196 30656 38208
rect 27816 38168 30144 38196
rect 30611 38168 30656 38196
rect 30650 38156 30656 38168
rect 30708 38156 30714 38208
rect 1104 38106 32016 38128
rect 1104 38054 7288 38106
rect 7340 38054 17592 38106
rect 17644 38054 27896 38106
rect 27948 38054 32016 38106
rect 1104 38032 32016 38054
rect 2406 37952 2412 38004
rect 2464 37992 2470 38004
rect 2685 37995 2743 38001
rect 2685 37992 2697 37995
rect 2464 37964 2697 37992
rect 2464 37952 2470 37964
rect 2685 37961 2697 37964
rect 2731 37961 2743 37995
rect 2685 37955 2743 37961
rect 5534 37952 5540 38004
rect 5592 37992 5598 38004
rect 5721 37995 5779 38001
rect 5721 37992 5733 37995
rect 5592 37964 5733 37992
rect 5592 37952 5598 37964
rect 5721 37961 5733 37964
rect 5767 37961 5779 37995
rect 5721 37955 5779 37961
rect 8389 37995 8447 38001
rect 8389 37961 8401 37995
rect 8435 37992 8447 37995
rect 8754 37992 8760 38004
rect 8435 37964 8760 37992
rect 8435 37961 8447 37964
rect 8389 37955 8447 37961
rect 8754 37952 8760 37964
rect 8812 37952 8818 38004
rect 10873 37995 10931 38001
rect 10873 37961 10885 37995
rect 10919 37992 10931 37995
rect 10962 37992 10968 38004
rect 10919 37964 10968 37992
rect 10919 37961 10931 37964
rect 10873 37955 10931 37961
rect 10962 37952 10968 37964
rect 11020 37952 11026 38004
rect 11882 37952 11888 38004
rect 11940 37952 11946 38004
rect 14182 37992 14188 38004
rect 11992 37964 14188 37992
rect 3050 37884 3056 37936
rect 3108 37924 3114 37936
rect 3108 37896 3372 37924
rect 3108 37884 3114 37896
rect 1302 37816 1308 37868
rect 1360 37856 1366 37868
rect 3344 37865 3372 37896
rect 4430 37884 4436 37936
rect 4488 37924 4494 37936
rect 5626 37924 5632 37936
rect 4488 37896 5632 37924
rect 4488 37884 4494 37896
rect 5626 37884 5632 37896
rect 5684 37924 5690 37936
rect 9306 37924 9312 37936
rect 5684 37896 9312 37924
rect 5684 37884 5690 37896
rect 9306 37884 9312 37896
rect 9364 37884 9370 37936
rect 11900 37924 11928 37952
rect 9508 37896 11928 37924
rect 1857 37859 1915 37865
rect 1857 37856 1869 37859
rect 1360 37828 1869 37856
rect 1360 37816 1366 37828
rect 1857 37825 1869 37828
rect 1903 37825 1915 37859
rect 1857 37819 1915 37825
rect 2869 37859 2927 37865
rect 2869 37825 2881 37859
rect 2915 37856 2927 37859
rect 3145 37859 3203 37865
rect 2915 37828 3096 37856
rect 2915 37825 2927 37828
rect 2869 37819 2927 37825
rect 2133 37655 2191 37661
rect 2133 37621 2145 37655
rect 2179 37652 2191 37655
rect 2314 37652 2320 37664
rect 2179 37624 2320 37652
rect 2179 37621 2191 37624
rect 2133 37615 2191 37621
rect 2314 37612 2320 37624
rect 2372 37612 2378 37664
rect 3068 37652 3096 37828
rect 3145 37825 3157 37859
rect 3191 37856 3203 37859
rect 3329 37859 3387 37865
rect 3191 37828 3280 37856
rect 3191 37825 3203 37828
rect 3145 37819 3203 37825
rect 3252 37720 3280 37828
rect 3329 37825 3341 37859
rect 3375 37825 3387 37859
rect 3329 37819 3387 37825
rect 4065 37859 4123 37865
rect 4065 37825 4077 37859
rect 4111 37856 4123 37859
rect 4246 37856 4252 37868
rect 4111 37828 4252 37856
rect 4111 37825 4123 37828
rect 4065 37819 4123 37825
rect 4246 37816 4252 37828
rect 4304 37816 4310 37868
rect 5534 37856 5540 37868
rect 5495 37828 5540 37856
rect 5534 37816 5540 37828
rect 5592 37816 5598 37868
rect 5810 37816 5816 37868
rect 5868 37856 5874 37868
rect 6546 37856 6552 37868
rect 5868 37828 6552 37856
rect 5868 37816 5874 37828
rect 6546 37816 6552 37828
rect 6604 37816 6610 37868
rect 7276 37859 7334 37865
rect 7276 37825 7288 37859
rect 7322 37856 7334 37859
rect 7558 37856 7564 37868
rect 7322 37828 7564 37856
rect 7322 37825 7334 37828
rect 7276 37819 7334 37825
rect 7558 37816 7564 37828
rect 7616 37816 7622 37868
rect 9508 37865 9536 37896
rect 9766 37865 9772 37868
rect 9493 37859 9551 37865
rect 9493 37825 9505 37859
rect 9539 37825 9551 37859
rect 9760 37856 9772 37865
rect 9727 37828 9772 37856
rect 9493 37819 9551 37825
rect 9760 37819 9772 37828
rect 9766 37816 9772 37819
rect 9824 37816 9830 37868
rect 11790 37816 11796 37868
rect 11848 37856 11854 37868
rect 11885 37859 11943 37865
rect 11885 37856 11897 37859
rect 11848 37828 11897 37856
rect 11848 37816 11854 37828
rect 11885 37825 11897 37828
rect 11931 37825 11943 37859
rect 11885 37819 11943 37825
rect 4154 37748 4160 37800
rect 4212 37788 4218 37800
rect 4341 37791 4399 37797
rect 4341 37788 4353 37791
rect 4212 37760 4353 37788
rect 4212 37748 4218 37760
rect 4341 37757 4353 37760
rect 4387 37757 4399 37791
rect 4341 37751 4399 37757
rect 5442 37748 5448 37800
rect 5500 37788 5506 37800
rect 7009 37791 7067 37797
rect 7009 37788 7021 37791
rect 5500 37760 7021 37788
rect 5500 37748 5506 37760
rect 7009 37757 7021 37760
rect 7055 37757 7067 37791
rect 7009 37751 7067 37757
rect 4172 37720 4200 37748
rect 3252 37692 4200 37720
rect 5534 37680 5540 37732
rect 5592 37720 5598 37732
rect 6086 37720 6092 37732
rect 5592 37692 6092 37720
rect 5592 37680 5598 37692
rect 6086 37680 6092 37692
rect 6144 37720 6150 37732
rect 11992 37720 12020 37964
rect 14182 37952 14188 37964
rect 14240 37952 14246 38004
rect 18874 37992 18880 38004
rect 15396 37964 18368 37992
rect 18835 37964 18880 37992
rect 12066 37884 12072 37936
rect 12124 37924 12130 37936
rect 15396 37924 15424 37964
rect 12124 37896 15424 37924
rect 15473 37927 15531 37933
rect 12124 37884 12130 37896
rect 15473 37893 15485 37927
rect 15519 37924 15531 37927
rect 15838 37924 15844 37936
rect 15519 37896 15844 37924
rect 15519 37893 15531 37896
rect 15473 37887 15531 37893
rect 15838 37884 15844 37896
rect 15896 37884 15902 37936
rect 17304 37927 17362 37933
rect 17304 37893 17316 37927
rect 17350 37924 17362 37927
rect 18230 37924 18236 37936
rect 17350 37896 18236 37924
rect 17350 37893 17362 37896
rect 17304 37887 17362 37893
rect 18230 37884 18236 37896
rect 18288 37884 18294 37936
rect 18340 37924 18368 37964
rect 18874 37952 18880 37964
rect 18932 37952 18938 38004
rect 21174 37992 21180 38004
rect 21135 37964 21180 37992
rect 21174 37952 21180 37964
rect 21232 37952 21238 38004
rect 22094 37952 22100 38004
rect 22152 37992 22158 38004
rect 23477 37995 23535 38001
rect 22152 37964 22197 37992
rect 22152 37952 22158 37964
rect 23477 37961 23489 37995
rect 23523 37992 23535 37995
rect 24394 37992 24400 38004
rect 23523 37964 24400 37992
rect 23523 37961 23535 37964
rect 23477 37955 23535 37961
rect 24394 37952 24400 37964
rect 24452 37952 24458 38004
rect 25317 37995 25375 38001
rect 25317 37961 25329 37995
rect 25363 37992 25375 37995
rect 26142 37992 26148 38004
rect 25363 37964 26148 37992
rect 25363 37961 25375 37964
rect 25317 37955 25375 37961
rect 26142 37952 26148 37964
rect 26200 37952 26206 38004
rect 26510 37952 26516 38004
rect 26568 37992 26574 38004
rect 26568 37964 27108 37992
rect 26568 37952 26574 37964
rect 18340 37896 22094 37924
rect 12621 37859 12679 37865
rect 12621 37856 12633 37859
rect 12084 37828 12633 37856
rect 12084 37800 12112 37828
rect 12621 37825 12633 37828
rect 12667 37856 12679 37859
rect 13630 37856 13636 37868
rect 12667 37828 13636 37856
rect 12667 37825 12679 37828
rect 12621 37819 12679 37825
rect 13630 37816 13636 37828
rect 13688 37816 13694 37868
rect 14001 37859 14059 37865
rect 14001 37825 14013 37859
rect 14047 37856 14059 37859
rect 14093 37859 14151 37865
rect 14093 37856 14105 37859
rect 14047 37828 14105 37856
rect 14047 37825 14059 37828
rect 14001 37819 14059 37825
rect 14093 37825 14105 37828
rect 14139 37825 14151 37859
rect 14274 37856 14280 37868
rect 14235 37828 14280 37856
rect 14093 37819 14151 37825
rect 14274 37816 14280 37828
rect 14332 37816 14338 37868
rect 14369 37859 14427 37865
rect 14369 37825 14381 37859
rect 14415 37825 14427 37859
rect 14369 37819 14427 37825
rect 14461 37859 14519 37865
rect 14461 37825 14473 37859
rect 14507 37825 14519 37859
rect 15105 37859 15163 37865
rect 15105 37856 15117 37859
rect 14461 37819 14519 37825
rect 14660 37828 15117 37856
rect 12066 37748 12072 37800
rect 12124 37748 12130 37800
rect 12161 37791 12219 37797
rect 12161 37757 12173 37791
rect 12207 37788 12219 37791
rect 12529 37791 12587 37797
rect 12529 37788 12541 37791
rect 12207 37760 12541 37788
rect 12207 37757 12219 37760
rect 12161 37751 12219 37757
rect 12529 37757 12541 37760
rect 12575 37757 12587 37791
rect 12529 37751 12587 37757
rect 12897 37791 12955 37797
rect 12897 37757 12909 37791
rect 12943 37788 12955 37791
rect 13722 37788 13728 37800
rect 12943 37760 13728 37788
rect 12943 37757 12955 37760
rect 12897 37751 12955 37757
rect 12618 37720 12624 37732
rect 6144 37692 6500 37720
rect 6144 37680 6150 37692
rect 3786 37652 3792 37664
rect 3068 37624 3792 37652
rect 3786 37612 3792 37624
rect 3844 37652 3850 37664
rect 6365 37655 6423 37661
rect 6365 37652 6377 37655
rect 3844 37624 6377 37652
rect 3844 37612 3850 37624
rect 6365 37621 6377 37624
rect 6411 37621 6423 37655
rect 6472 37652 6500 37692
rect 10428 37692 12020 37720
rect 12084 37692 12624 37720
rect 10428 37652 10456 37692
rect 6472 37624 10456 37652
rect 11701 37655 11759 37661
rect 6365 37615 6423 37621
rect 11701 37621 11713 37655
rect 11747 37652 11759 37655
rect 11974 37652 11980 37664
rect 11747 37624 11980 37652
rect 11747 37621 11759 37624
rect 11701 37615 11759 37621
rect 11974 37612 11980 37624
rect 12032 37612 12038 37664
rect 12084 37661 12112 37692
rect 12618 37680 12624 37692
rect 12676 37680 12682 37732
rect 12710 37680 12716 37732
rect 12768 37720 12774 37732
rect 12912 37720 12940 37751
rect 13722 37748 13728 37760
rect 13780 37748 13786 37800
rect 14182 37748 14188 37800
rect 14240 37788 14246 37800
rect 14384 37788 14412 37819
rect 14240 37760 14412 37788
rect 14240 37748 14246 37760
rect 14476 37732 14504 37819
rect 12768 37692 12940 37720
rect 12768 37680 12774 37692
rect 14458 37680 14464 37732
rect 14516 37680 14522 37732
rect 14660 37729 14688 37828
rect 15105 37825 15117 37828
rect 15151 37825 15163 37859
rect 15105 37819 15163 37825
rect 15194 37816 15200 37868
rect 15252 37856 15258 37868
rect 15252 37828 15297 37856
rect 15252 37816 15258 37828
rect 15378 37816 15384 37868
rect 15436 37856 15442 37868
rect 15436 37828 15481 37856
rect 15436 37816 15442 37828
rect 15562 37816 15568 37868
rect 15620 37865 15626 37868
rect 15620 37856 15628 37865
rect 19058 37856 19064 37868
rect 15620 37828 15665 37856
rect 19019 37828 19064 37856
rect 15620 37819 15628 37828
rect 15620 37816 15626 37819
rect 19058 37816 19064 37828
rect 19116 37816 19122 37868
rect 19334 37856 19340 37868
rect 19295 37828 19340 37856
rect 19334 37816 19340 37828
rect 19392 37816 19398 37868
rect 19610 37816 19616 37868
rect 19668 37856 19674 37868
rect 19797 37859 19855 37865
rect 19797 37856 19809 37859
rect 19668 37828 19809 37856
rect 19668 37816 19674 37828
rect 19797 37825 19809 37828
rect 19843 37825 19855 37859
rect 19797 37819 19855 37825
rect 20064 37859 20122 37865
rect 20064 37825 20076 37859
rect 20110 37856 20122 37859
rect 20530 37856 20536 37868
rect 20110 37828 20536 37856
rect 20110 37825 20122 37828
rect 20064 37819 20122 37825
rect 20530 37816 20536 37828
rect 20588 37816 20594 37868
rect 14645 37723 14703 37729
rect 14645 37689 14657 37723
rect 14691 37689 14703 37723
rect 14645 37683 14703 37689
rect 15194 37680 15200 37732
rect 15252 37720 15258 37732
rect 15580 37720 15608 37816
rect 16850 37748 16856 37800
rect 16908 37788 16914 37800
rect 17037 37791 17095 37797
rect 17037 37788 17049 37791
rect 16908 37760 17049 37788
rect 16908 37748 16914 37760
rect 17037 37757 17049 37760
rect 17083 37757 17095 37791
rect 17037 37751 17095 37757
rect 19150 37748 19156 37800
rect 19208 37788 19214 37800
rect 19245 37791 19303 37797
rect 19245 37788 19257 37791
rect 19208 37760 19257 37788
rect 19208 37748 19214 37760
rect 19245 37757 19257 37760
rect 19291 37757 19303 37791
rect 19245 37751 19303 37757
rect 15252 37692 15608 37720
rect 22066 37720 22094 37896
rect 22922 37884 22928 37936
rect 22980 37924 22986 37936
rect 23109 37927 23167 37933
rect 23109 37924 23121 37927
rect 22980 37896 23121 37924
rect 22980 37884 22986 37896
rect 23109 37893 23121 37896
rect 23155 37893 23167 37927
rect 23109 37887 23167 37893
rect 23325 37927 23383 37933
rect 23325 37893 23337 37927
rect 23371 37924 23383 37927
rect 24762 37924 24768 37936
rect 23371 37896 24768 37924
rect 23371 37893 23383 37896
rect 23325 37887 23383 37893
rect 24762 37884 24768 37896
rect 24820 37884 24826 37936
rect 26326 37924 26332 37936
rect 25792 37896 26332 37924
rect 22278 37856 22284 37868
rect 22239 37828 22284 37856
rect 22278 37816 22284 37828
rect 22336 37816 22342 37868
rect 22462 37856 22468 37868
rect 22423 37828 22468 37856
rect 22462 37816 22468 37828
rect 22520 37816 22526 37868
rect 24210 37856 24216 37868
rect 24171 37828 24216 37856
rect 24210 37816 24216 37828
rect 24268 37816 24274 37868
rect 24302 37816 24308 37868
rect 24360 37856 24366 37868
rect 24486 37856 24492 37868
rect 24360 37828 24405 37856
rect 24447 37828 24492 37856
rect 24360 37816 24366 37828
rect 24486 37816 24492 37828
rect 24544 37816 24550 37868
rect 24581 37859 24639 37865
rect 24581 37825 24593 37859
rect 24627 37856 24639 37859
rect 24673 37859 24731 37865
rect 24673 37856 24685 37859
rect 24627 37828 24685 37856
rect 24627 37825 24639 37828
rect 24581 37819 24639 37825
rect 24673 37825 24685 37828
rect 24719 37825 24731 37859
rect 24673 37819 24731 37825
rect 25314 37816 25320 37868
rect 25372 37856 25378 37868
rect 25792 37865 25820 37896
rect 26326 37884 26332 37896
rect 26384 37884 26390 37936
rect 25501 37859 25559 37865
rect 25501 37856 25513 37859
rect 25372 37828 25513 37856
rect 25372 37816 25378 37828
rect 25501 37825 25513 37828
rect 25547 37825 25559 37859
rect 25501 37819 25559 37825
rect 25777 37859 25835 37865
rect 25777 37825 25789 37859
rect 25823 37825 25835 37859
rect 25958 37856 25964 37868
rect 25919 37828 25964 37856
rect 25777 37819 25835 37825
rect 25958 37816 25964 37828
rect 26016 37816 26022 37868
rect 26970 37856 26976 37868
rect 26931 37828 26976 37856
rect 26970 37816 26976 37828
rect 27028 37816 27034 37868
rect 27080 37865 27108 37964
rect 27430 37952 27436 38004
rect 27488 37992 27494 38004
rect 27617 37995 27675 38001
rect 27617 37992 27629 37995
rect 27488 37964 27629 37992
rect 27488 37952 27494 37964
rect 27617 37961 27629 37964
rect 27663 37961 27675 37995
rect 31110 37992 31116 38004
rect 27617 37955 27675 37961
rect 27899 37964 31116 37992
rect 27066 37859 27124 37865
rect 27066 37825 27078 37859
rect 27112 37825 27124 37859
rect 27246 37856 27252 37868
rect 27207 37828 27252 37856
rect 27066 37819 27124 37825
rect 27246 37816 27252 37828
rect 27304 37816 27310 37868
rect 27338 37850 27344 37902
rect 27396 37865 27402 37902
rect 27396 37850 27407 37865
rect 27349 37825 27361 37850
rect 27395 37825 27407 37850
rect 27349 37819 27407 37825
rect 27479 37859 27537 37865
rect 27479 37825 27491 37859
rect 27525 37856 27537 37859
rect 27614 37856 27620 37868
rect 27525 37828 27620 37856
rect 27525 37825 27537 37828
rect 27479 37819 27537 37825
rect 27614 37816 27620 37828
rect 27672 37816 27678 37868
rect 22557 37791 22615 37797
rect 22557 37757 22569 37791
rect 22603 37788 22615 37791
rect 22922 37788 22928 37800
rect 22603 37760 22928 37788
rect 22603 37757 22615 37760
rect 22557 37751 22615 37757
rect 22922 37748 22928 37760
rect 22980 37748 22986 37800
rect 24029 37791 24087 37797
rect 24029 37757 24041 37791
rect 24075 37788 24087 37791
rect 25866 37788 25872 37800
rect 24075 37760 25872 37788
rect 24075 37757 24087 37760
rect 24029 37751 24087 37757
rect 25866 37748 25872 37760
rect 25924 37748 25930 37800
rect 27264 37788 27292 37816
rect 27798 37788 27804 37800
rect 27264 37760 27804 37788
rect 27798 37748 27804 37760
rect 27856 37748 27862 37800
rect 27899 37720 27927 37964
rect 31110 37952 31116 37964
rect 31168 37952 31174 38004
rect 29546 37924 29552 37936
rect 28092 37896 29552 37924
rect 28092 37865 28120 37896
rect 29546 37884 29552 37896
rect 29604 37924 29610 37936
rect 30184 37927 30242 37933
rect 29604 37896 29684 37924
rect 29604 37884 29610 37896
rect 28077 37859 28135 37865
rect 28077 37825 28089 37859
rect 28123 37825 28135 37859
rect 28077 37819 28135 37825
rect 28344 37859 28402 37865
rect 28344 37825 28356 37859
rect 28390 37856 28402 37859
rect 28390 37828 29500 37856
rect 28390 37825 28402 37828
rect 28344 37819 28402 37825
rect 29472 37788 29500 37828
rect 29656 37800 29684 37896
rect 30184 37893 30196 37927
rect 30230 37924 30242 37927
rect 30650 37924 30656 37936
rect 30230 37896 30656 37924
rect 30230 37893 30242 37896
rect 30184 37887 30242 37893
rect 30650 37884 30656 37896
rect 30708 37884 30714 37936
rect 29546 37788 29552 37800
rect 29472 37760 29552 37788
rect 29546 37748 29552 37760
rect 29604 37748 29610 37800
rect 29638 37748 29644 37800
rect 29696 37788 29702 37800
rect 29917 37791 29975 37797
rect 29917 37788 29929 37791
rect 29696 37760 29929 37788
rect 29696 37748 29702 37760
rect 29917 37757 29929 37760
rect 29963 37757 29975 37791
rect 29917 37751 29975 37757
rect 22066 37692 27927 37720
rect 15252 37680 15258 37692
rect 12069 37655 12127 37661
rect 12069 37621 12081 37655
rect 12115 37621 12127 37655
rect 12069 37615 12127 37621
rect 12529 37655 12587 37661
rect 12529 37621 12541 37655
rect 12575 37652 12587 37655
rect 13262 37652 13268 37664
rect 12575 37624 13268 37652
rect 12575 37621 12587 37624
rect 12529 37615 12587 37621
rect 13262 37612 13268 37624
rect 13320 37612 13326 37664
rect 14001 37655 14059 37661
rect 14001 37621 14013 37655
rect 14047 37652 14059 37655
rect 15470 37652 15476 37664
rect 14047 37624 15476 37652
rect 14047 37621 14059 37624
rect 14001 37615 14059 37621
rect 15470 37612 15476 37624
rect 15528 37612 15534 37664
rect 15746 37652 15752 37664
rect 15707 37624 15752 37652
rect 15746 37612 15752 37624
rect 15804 37612 15810 37664
rect 18046 37612 18052 37664
rect 18104 37652 18110 37664
rect 18414 37652 18420 37664
rect 18104 37624 18420 37652
rect 18104 37612 18110 37624
rect 18414 37612 18420 37624
rect 18472 37612 18478 37664
rect 23290 37652 23296 37664
rect 23251 37624 23296 37652
rect 23290 37612 23296 37624
rect 23348 37612 23354 37664
rect 24394 37612 24400 37664
rect 24452 37652 24458 37664
rect 24673 37655 24731 37661
rect 24673 37652 24685 37655
rect 24452 37624 24685 37652
rect 24452 37612 24458 37624
rect 24673 37621 24685 37624
rect 24719 37652 24731 37655
rect 28718 37652 28724 37664
rect 24719 37624 28724 37652
rect 24719 37621 24731 37624
rect 24673 37615 24731 37621
rect 28718 37612 28724 37624
rect 28776 37612 28782 37664
rect 28994 37612 29000 37664
rect 29052 37652 29058 37664
rect 29457 37655 29515 37661
rect 29457 37652 29469 37655
rect 29052 37624 29469 37652
rect 29052 37612 29058 37624
rect 29457 37621 29469 37624
rect 29503 37621 29515 37655
rect 31294 37652 31300 37664
rect 31255 37624 31300 37652
rect 29457 37615 29515 37621
rect 31294 37612 31300 37624
rect 31352 37612 31358 37664
rect 1104 37562 32016 37584
rect 1104 37510 2136 37562
rect 2188 37510 12440 37562
rect 12492 37510 22744 37562
rect 22796 37510 32016 37562
rect 1104 37488 32016 37510
rect 2774 37408 2780 37460
rect 2832 37448 2838 37460
rect 7558 37448 7564 37460
rect 2832 37420 2877 37448
rect 7519 37420 7564 37448
rect 2832 37408 2838 37420
rect 7558 37408 7564 37420
rect 7616 37408 7622 37460
rect 8573 37451 8631 37457
rect 8573 37417 8585 37451
rect 8619 37448 8631 37451
rect 11609 37451 11667 37457
rect 11609 37448 11621 37451
rect 8619 37420 11621 37448
rect 8619 37417 8631 37420
rect 8573 37411 8631 37417
rect 11609 37417 11621 37420
rect 11655 37417 11667 37451
rect 11609 37411 11667 37417
rect 12342 37408 12348 37460
rect 12400 37448 12406 37460
rect 13078 37448 13084 37460
rect 12400 37420 13084 37448
rect 12400 37408 12406 37420
rect 13078 37408 13084 37420
rect 13136 37408 13142 37460
rect 13630 37408 13636 37460
rect 13688 37448 13694 37460
rect 15930 37448 15936 37460
rect 13688 37420 15936 37448
rect 13688 37408 13694 37420
rect 15930 37408 15936 37420
rect 15988 37448 15994 37460
rect 16669 37451 16727 37457
rect 16669 37448 16681 37451
rect 15988 37420 16681 37448
rect 15988 37408 15994 37420
rect 16669 37417 16681 37420
rect 16715 37417 16727 37451
rect 16669 37411 16727 37417
rect 20530 37408 20536 37460
rect 20588 37448 20594 37460
rect 20625 37451 20683 37457
rect 20625 37448 20637 37451
rect 20588 37420 20637 37448
rect 20588 37408 20594 37420
rect 20625 37417 20637 37420
rect 20671 37417 20683 37451
rect 20625 37411 20683 37417
rect 22925 37451 22983 37457
rect 22925 37417 22937 37451
rect 22971 37448 22983 37451
rect 23290 37448 23296 37460
rect 22971 37420 23296 37448
rect 22971 37417 22983 37420
rect 22925 37411 22983 37417
rect 23290 37408 23296 37420
rect 23348 37408 23354 37460
rect 23474 37408 23480 37460
rect 23532 37448 23538 37460
rect 23661 37451 23719 37457
rect 23661 37448 23673 37451
rect 23532 37420 23673 37448
rect 23532 37408 23538 37420
rect 23661 37417 23673 37420
rect 23707 37417 23719 37451
rect 23661 37411 23719 37417
rect 23845 37451 23903 37457
rect 23845 37417 23857 37451
rect 23891 37448 23903 37451
rect 24670 37448 24676 37460
rect 23891 37420 24676 37448
rect 23891 37417 23903 37420
rect 23845 37411 23903 37417
rect 6822 37380 6828 37392
rect 5276 37352 6828 37380
rect 5276 37312 5304 37352
rect 6822 37340 6828 37352
rect 6880 37340 6886 37392
rect 11698 37380 11704 37392
rect 7116 37352 11704 37380
rect 6086 37312 6092 37324
rect 4724 37284 5304 37312
rect 5644 37284 5948 37312
rect 6047 37284 6092 37312
rect 1394 37244 1400 37256
rect 1355 37216 1400 37244
rect 1394 37204 1400 37216
rect 1452 37204 1458 37256
rect 4338 37244 4344 37256
rect 4299 37216 4344 37244
rect 4338 37204 4344 37216
rect 4396 37204 4402 37256
rect 4434 37247 4492 37253
rect 4434 37213 4446 37247
rect 4480 37213 4492 37247
rect 4434 37207 4492 37213
rect 4617 37247 4675 37253
rect 4617 37213 4629 37247
rect 4663 37244 4675 37247
rect 4724 37244 4752 37284
rect 4663 37216 4752 37244
rect 4847 37247 4905 37253
rect 4663 37213 4675 37216
rect 4617 37207 4675 37213
rect 4847 37213 4859 37247
rect 4893 37244 4905 37247
rect 5644 37244 5672 37284
rect 4893 37216 5672 37244
rect 4893 37213 4905 37216
rect 4847 37207 4905 37213
rect 0 37176 800 37190
rect 1302 37176 1308 37188
rect 0 37148 1308 37176
rect 0 37134 800 37148
rect 1302 37136 1308 37148
rect 1360 37136 1366 37188
rect 1486 37136 1492 37188
rect 1544 37176 1550 37188
rect 1642 37179 1700 37185
rect 1642 37176 1654 37179
rect 1544 37148 1654 37176
rect 1544 37136 1550 37148
rect 1642 37145 1654 37148
rect 1688 37145 1700 37179
rect 1642 37139 1700 37145
rect 3234 37136 3240 37188
rect 3292 37176 3298 37188
rect 4448 37176 4476 37207
rect 5718 37204 5724 37256
rect 5776 37244 5782 37256
rect 5813 37247 5871 37253
rect 5813 37244 5825 37247
rect 5776 37216 5825 37244
rect 5776 37204 5782 37216
rect 5813 37213 5825 37216
rect 5859 37213 5871 37247
rect 5920 37244 5948 37284
rect 6086 37272 6092 37284
rect 6144 37272 6150 37324
rect 7116 37321 7144 37352
rect 11698 37340 11704 37352
rect 11756 37340 11762 37392
rect 13354 37340 13360 37392
rect 13412 37380 13418 37392
rect 13541 37383 13599 37389
rect 13541 37380 13553 37383
rect 13412 37352 13553 37380
rect 13412 37340 13418 37352
rect 13541 37349 13553 37352
rect 13587 37380 13599 37383
rect 13587 37352 14872 37380
rect 13587 37349 13599 37352
rect 13541 37343 13599 37349
rect 7101 37315 7159 37321
rect 7101 37281 7113 37315
rect 7147 37281 7159 37315
rect 8018 37312 8024 37324
rect 7979 37284 8024 37312
rect 7101 37275 7159 37281
rect 8018 37272 8024 37284
rect 8076 37272 8082 37324
rect 8110 37272 8116 37324
rect 8168 37312 8174 37324
rect 10873 37315 10931 37321
rect 10873 37312 10885 37315
rect 8168 37284 10885 37312
rect 8168 37272 8174 37284
rect 10873 37281 10885 37284
rect 10919 37281 10931 37315
rect 10873 37275 10931 37281
rect 11882 37272 11888 37324
rect 11940 37312 11946 37324
rect 12161 37315 12219 37321
rect 12161 37312 12173 37315
rect 11940 37284 12173 37312
rect 11940 37272 11946 37284
rect 12161 37281 12173 37284
rect 12207 37281 12219 37315
rect 12161 37275 12219 37281
rect 5920 37216 6408 37244
rect 5813 37207 5871 37213
rect 3292 37148 4476 37176
rect 3292 37136 3298 37148
rect 4706 37136 4712 37188
rect 4764 37176 4770 37188
rect 5905 37179 5963 37185
rect 5905 37176 5917 37179
rect 4764 37148 4809 37176
rect 5000 37148 5917 37176
rect 4764 37136 4770 37148
rect 5000 37117 5028 37148
rect 5905 37145 5917 37148
rect 5951 37145 5963 37179
rect 6380 37176 6408 37216
rect 6454 37204 6460 37256
rect 6512 37244 6518 37256
rect 6825 37247 6883 37253
rect 6825 37244 6837 37247
rect 6512 37216 6837 37244
rect 6512 37204 6518 37216
rect 6825 37213 6837 37216
rect 6871 37213 6883 37247
rect 7006 37244 7012 37256
rect 6967 37216 7012 37244
rect 6825 37207 6883 37213
rect 7006 37204 7012 37216
rect 7064 37244 7070 37256
rect 7742 37244 7748 37256
rect 7064 37216 7236 37244
rect 7703 37216 7748 37244
rect 7064 37204 7070 37216
rect 7208 37176 7236 37216
rect 7742 37204 7748 37216
rect 7800 37204 7806 37256
rect 7929 37247 7987 37253
rect 7929 37213 7941 37247
rect 7975 37244 7987 37247
rect 8938 37244 8944 37256
rect 7975 37216 8944 37244
rect 7975 37213 7987 37216
rect 7929 37207 7987 37213
rect 8938 37204 8944 37216
rect 8996 37204 9002 37256
rect 9033 37247 9091 37253
rect 9033 37213 9045 37247
rect 9079 37213 9091 37247
rect 9214 37244 9220 37256
rect 9175 37216 9220 37244
rect 9033 37207 9091 37213
rect 8573 37179 8631 37185
rect 8573 37176 8585 37179
rect 6380 37148 7144 37176
rect 7208 37148 8585 37176
rect 5905 37139 5963 37145
rect 7116 37120 7144 37148
rect 8573 37145 8585 37148
rect 8619 37145 8631 37179
rect 8573 37139 8631 37145
rect 8662 37136 8668 37188
rect 8720 37176 8726 37188
rect 9048 37176 9076 37207
rect 9214 37204 9220 37216
rect 9272 37204 9278 37256
rect 9398 37204 9404 37256
rect 9456 37244 9462 37256
rect 10505 37247 10563 37253
rect 10505 37244 10517 37247
rect 9456 37216 10517 37244
rect 9456 37204 9462 37216
rect 10505 37213 10517 37216
rect 10551 37213 10563 37247
rect 10505 37207 10563 37213
rect 10597 37247 10655 37253
rect 10597 37213 10609 37247
rect 10643 37244 10655 37247
rect 10686 37244 10692 37256
rect 10643 37216 10692 37244
rect 10643 37213 10655 37216
rect 10597 37207 10655 37213
rect 10042 37176 10048 37188
rect 8720 37148 10048 37176
rect 8720 37136 8726 37148
rect 10042 37136 10048 37148
rect 10100 37136 10106 37188
rect 4985 37111 5043 37117
rect 4985 37077 4997 37111
rect 5031 37077 5043 37111
rect 4985 37071 5043 37077
rect 5445 37111 5503 37117
rect 5445 37077 5457 37111
rect 5491 37108 5503 37111
rect 6270 37108 6276 37120
rect 5491 37080 6276 37108
rect 5491 37077 5503 37080
rect 5445 37071 5503 37077
rect 6270 37068 6276 37080
rect 6328 37068 6334 37120
rect 6638 37108 6644 37120
rect 6599 37080 6644 37108
rect 6638 37068 6644 37080
rect 6696 37068 6702 37120
rect 7098 37068 7104 37120
rect 7156 37108 7162 37120
rect 9125 37111 9183 37117
rect 9125 37108 9137 37111
rect 7156 37080 9137 37108
rect 7156 37068 7162 37080
rect 9125 37077 9137 37080
rect 9171 37077 9183 37111
rect 10318 37108 10324 37120
rect 10279 37080 10324 37108
rect 9125 37071 9183 37077
rect 10318 37068 10324 37080
rect 10376 37068 10382 37120
rect 10520 37108 10548 37207
rect 10686 37204 10692 37216
rect 10744 37204 10750 37256
rect 10965 37247 11023 37253
rect 10965 37213 10977 37247
rect 11011 37244 11023 37247
rect 11011 37216 11744 37244
rect 11011 37213 11023 37216
rect 10965 37207 11023 37213
rect 11514 37176 11520 37188
rect 11475 37148 11520 37176
rect 11514 37136 11520 37148
rect 11572 37136 11578 37188
rect 11238 37108 11244 37120
rect 10520 37080 11244 37108
rect 11238 37068 11244 37080
rect 11296 37068 11302 37120
rect 11716 37108 11744 37216
rect 12066 37204 12072 37256
rect 12124 37244 12130 37256
rect 14550 37244 14556 37256
rect 12124 37216 14228 37244
rect 14511 37216 14556 37244
rect 12124 37204 12130 37216
rect 11974 37136 11980 37188
rect 12032 37176 12038 37188
rect 12406 37179 12464 37185
rect 12406 37176 12418 37179
rect 12032 37148 12418 37176
rect 12032 37136 12038 37148
rect 12406 37145 12418 37148
rect 12452 37145 12464 37179
rect 13814 37176 13820 37188
rect 12406 37139 12464 37145
rect 13464 37148 13820 37176
rect 13464 37108 13492 37148
rect 13814 37136 13820 37148
rect 13872 37136 13878 37188
rect 11716 37080 13492 37108
rect 14200 37108 14228 37216
rect 14550 37204 14556 37216
rect 14608 37204 14614 37256
rect 14642 37204 14648 37256
rect 14700 37244 14706 37256
rect 14844 37244 14872 37352
rect 14918 37340 14924 37392
rect 14976 37380 14982 37392
rect 15286 37380 15292 37392
rect 14976 37352 15292 37380
rect 14976 37340 14982 37352
rect 15286 37340 15292 37352
rect 15344 37380 15350 37392
rect 16482 37380 16488 37392
rect 15344 37352 16488 37380
rect 15344 37340 15350 37352
rect 16482 37340 16488 37352
rect 16540 37340 16546 37392
rect 19150 37340 19156 37392
rect 19208 37380 19214 37392
rect 21821 37383 21879 37389
rect 21821 37380 21833 37383
rect 19208 37352 21833 37380
rect 19208 37340 19214 37352
rect 21821 37349 21833 37352
rect 21867 37349 21879 37383
rect 23676 37380 23704 37411
rect 24670 37408 24676 37420
rect 24728 37408 24734 37460
rect 25777 37451 25835 37457
rect 25777 37417 25789 37451
rect 25823 37448 25835 37451
rect 27062 37448 27068 37460
rect 25823 37420 27068 37448
rect 25823 37417 25835 37420
rect 25777 37411 25835 37417
rect 27062 37408 27068 37420
rect 27120 37408 27126 37460
rect 27154 37408 27160 37460
rect 27212 37448 27218 37460
rect 27893 37451 27951 37457
rect 27893 37448 27905 37451
rect 27212 37420 27905 37448
rect 27212 37408 27218 37420
rect 27893 37417 27905 37420
rect 27939 37417 27951 37451
rect 27893 37411 27951 37417
rect 28828 37420 29040 37448
rect 24578 37380 24584 37392
rect 23676 37352 24584 37380
rect 21821 37343 21879 37349
rect 24578 37340 24584 37352
rect 24636 37380 24642 37392
rect 25041 37383 25099 37389
rect 25041 37380 25053 37383
rect 24636 37352 25053 37380
rect 24636 37340 24642 37352
rect 25041 37349 25053 37352
rect 25087 37349 25099 37383
rect 25041 37343 25099 37349
rect 26234 37340 26240 37392
rect 26292 37380 26298 37392
rect 26697 37383 26755 37389
rect 26697 37380 26709 37383
rect 26292 37352 26709 37380
rect 26292 37340 26298 37352
rect 26697 37349 26709 37352
rect 26743 37380 26755 37383
rect 27246 37380 27252 37392
rect 26743 37352 27252 37380
rect 26743 37349 26755 37352
rect 26697 37343 26755 37349
rect 27246 37340 27252 37352
rect 27304 37340 27310 37392
rect 27614 37340 27620 37392
rect 27672 37380 27678 37392
rect 28718 37380 28724 37392
rect 27672 37352 28724 37380
rect 27672 37340 27678 37352
rect 28718 37340 28724 37352
rect 28776 37340 28782 37392
rect 15654 37312 15660 37324
rect 15615 37284 15660 37312
rect 15654 37272 15660 37284
rect 15712 37272 15718 37324
rect 19337 37315 19395 37321
rect 19337 37281 19349 37315
rect 19383 37312 19395 37315
rect 19702 37312 19708 37324
rect 19383 37284 19708 37312
rect 19383 37281 19395 37284
rect 19337 37275 19395 37281
rect 19702 37272 19708 37284
rect 19760 37272 19766 37324
rect 21085 37315 21143 37321
rect 21085 37281 21097 37315
rect 21131 37312 21143 37315
rect 21726 37312 21732 37324
rect 21131 37284 21732 37312
rect 21131 37281 21143 37284
rect 21085 37275 21143 37281
rect 21726 37272 21732 37284
rect 21784 37272 21790 37324
rect 24210 37272 24216 37324
rect 24268 37312 24274 37324
rect 27982 37312 27988 37324
rect 24268 37284 27988 37312
rect 24268 37272 24274 37284
rect 14921 37247 14979 37253
rect 14921 37244 14933 37247
rect 14700 37216 14745 37244
rect 14844 37216 14933 37244
rect 14700 37204 14706 37216
rect 14921 37213 14933 37216
rect 14967 37213 14979 37247
rect 14921 37207 14979 37213
rect 15059 37247 15117 37253
rect 15059 37213 15071 37247
rect 15105 37244 15117 37247
rect 15194 37244 15200 37256
rect 15105 37216 15200 37244
rect 15105 37213 15117 37216
rect 15059 37207 15117 37213
rect 15194 37204 15200 37216
rect 15252 37204 15258 37256
rect 15286 37204 15292 37256
rect 15344 37244 15350 37256
rect 15841 37247 15899 37253
rect 15841 37244 15853 37247
rect 15344 37216 15853 37244
rect 15344 37204 15350 37216
rect 15841 37213 15853 37216
rect 15887 37213 15899 37247
rect 17770 37244 17776 37256
rect 17731 37216 17776 37244
rect 15841 37207 15899 37213
rect 17770 37204 17776 37216
rect 17828 37204 17834 37256
rect 17862 37204 17868 37256
rect 17920 37244 17926 37256
rect 17957 37247 18015 37253
rect 17957 37244 17969 37247
rect 17920 37216 17969 37244
rect 17920 37204 17926 37216
rect 17957 37213 17969 37216
rect 18003 37213 18015 37247
rect 18230 37244 18236 37256
rect 18191 37216 18236 37244
rect 17957 37207 18015 37213
rect 18230 37204 18236 37216
rect 18288 37204 18294 37256
rect 18414 37204 18420 37256
rect 18472 37253 18478 37256
rect 18472 37247 18487 37253
rect 18475 37213 18487 37247
rect 18472 37207 18487 37213
rect 19613 37247 19671 37253
rect 19613 37213 19625 37247
rect 19659 37213 19671 37247
rect 19613 37207 19671 37213
rect 18472 37204 18478 37207
rect 14826 37176 14832 37188
rect 14787 37148 14832 37176
rect 14826 37136 14832 37148
rect 14884 37136 14890 37188
rect 16025 37179 16083 37185
rect 16025 37176 16037 37179
rect 15028 37148 16037 37176
rect 15028 37108 15056 37148
rect 16025 37145 16037 37148
rect 16071 37145 16083 37179
rect 16025 37139 16083 37145
rect 16577 37179 16635 37185
rect 16577 37145 16589 37179
rect 16623 37176 16635 37179
rect 17310 37176 17316 37188
rect 16623 37148 17316 37176
rect 16623 37145 16635 37148
rect 16577 37139 16635 37145
rect 17310 37136 17316 37148
rect 17368 37136 17374 37188
rect 18248 37176 18276 37204
rect 19628 37176 19656 37207
rect 19978 37204 19984 37256
rect 20036 37244 20042 37256
rect 20809 37247 20867 37253
rect 20809 37244 20821 37247
rect 20036 37216 20821 37244
rect 20036 37204 20042 37216
rect 20809 37213 20821 37216
rect 20855 37213 20867 37247
rect 20990 37244 20996 37256
rect 20951 37216 20996 37244
rect 20809 37207 20867 37213
rect 20990 37204 20996 37216
rect 21048 37204 21054 37256
rect 21542 37204 21548 37256
rect 21600 37244 21606 37256
rect 21637 37247 21695 37253
rect 21637 37244 21649 37247
rect 21600 37216 21649 37244
rect 21600 37204 21606 37216
rect 21637 37213 21649 37216
rect 21683 37213 21695 37247
rect 21637 37207 21695 37213
rect 22833 37247 22891 37253
rect 22833 37213 22845 37247
rect 22879 37213 22891 37247
rect 23014 37244 23020 37256
rect 22975 37216 23020 37244
rect 22833 37207 22891 37213
rect 18248 37148 19656 37176
rect 14200 37080 15056 37108
rect 15197 37111 15255 37117
rect 15197 37077 15209 37111
rect 15243 37108 15255 37111
rect 15838 37108 15844 37120
rect 15243 37080 15844 37108
rect 15243 37077 15255 37080
rect 15197 37071 15255 37077
rect 15838 37068 15844 37080
rect 15896 37068 15902 37120
rect 16942 37068 16948 37120
rect 17000 37108 17006 37120
rect 17678 37108 17684 37120
rect 17000 37080 17684 37108
rect 17000 37068 17006 37080
rect 17678 37068 17684 37080
rect 17736 37068 17742 37120
rect 22848 37108 22876 37207
rect 23014 37204 23020 37216
rect 23072 37204 23078 37256
rect 24026 37204 24032 37256
rect 24084 37244 24090 37256
rect 24397 37247 24455 37253
rect 24397 37244 24409 37247
rect 24084 37216 24409 37244
rect 24084 37204 24090 37216
rect 24397 37213 24409 37216
rect 24443 37213 24455 37247
rect 24397 37207 24455 37213
rect 24581 37247 24639 37253
rect 24581 37213 24593 37247
rect 24627 37213 24639 37247
rect 24581 37207 24639 37213
rect 24949 37247 25007 37253
rect 24949 37213 24961 37247
rect 24995 37244 25007 37247
rect 25041 37247 25099 37253
rect 25041 37244 25053 37247
rect 24995 37216 25053 37244
rect 24995 37213 25007 37216
rect 24949 37207 25007 37213
rect 25041 37213 25053 37216
rect 25087 37213 25099 37247
rect 25958 37244 25964 37256
rect 25919 37216 25964 37244
rect 25041 37207 25099 37213
rect 23382 37136 23388 37188
rect 23440 37176 23446 37188
rect 23477 37179 23535 37185
rect 23477 37176 23489 37179
rect 23440 37148 23489 37176
rect 23440 37136 23446 37148
rect 23477 37145 23489 37148
rect 23523 37176 23535 37179
rect 24596 37176 24624 37207
rect 25958 37204 25964 37216
rect 26016 37204 26022 37256
rect 26050 37204 26056 37256
rect 26108 37244 26114 37256
rect 26252 37253 26280 37284
rect 26145 37247 26203 37253
rect 26145 37244 26157 37247
rect 26108 37216 26157 37244
rect 26108 37204 26114 37216
rect 26145 37213 26157 37216
rect 26191 37213 26203 37247
rect 26145 37207 26203 37213
rect 26237 37247 26295 37253
rect 26237 37213 26249 37247
rect 26283 37213 26295 37247
rect 26237 37207 26295 37213
rect 26697 37247 26755 37253
rect 26697 37213 26709 37247
rect 26743 37213 26755 37247
rect 26697 37207 26755 37213
rect 23523 37148 24624 37176
rect 23523 37145 23535 37148
rect 23477 37139 23535 37145
rect 24762 37136 24768 37188
rect 24820 37176 24826 37188
rect 26712 37176 26740 37207
rect 26786 37204 26792 37256
rect 26844 37244 26850 37256
rect 26881 37247 26939 37253
rect 26881 37244 26893 37247
rect 26844 37216 26893 37244
rect 26844 37204 26850 37216
rect 26881 37213 26893 37216
rect 26927 37213 26939 37247
rect 26881 37207 26939 37213
rect 27341 37247 27399 37253
rect 27341 37213 27353 37247
rect 27387 37244 27399 37247
rect 27430 37244 27436 37256
rect 27387 37216 27436 37244
rect 27387 37213 27399 37216
rect 27341 37207 27399 37213
rect 27430 37204 27436 37216
rect 27488 37204 27494 37256
rect 27724 37253 27752 37284
rect 27982 37272 27988 37284
rect 28040 37272 28046 37324
rect 28828 37312 28856 37420
rect 29012 37380 29040 37420
rect 29178 37408 29184 37460
rect 29236 37448 29242 37460
rect 29822 37448 29828 37460
rect 29236 37420 29828 37448
rect 29236 37408 29242 37420
rect 29822 37408 29828 37420
rect 29880 37408 29886 37460
rect 29730 37380 29736 37392
rect 29012 37352 29736 37380
rect 29730 37340 29736 37352
rect 29788 37340 29794 37392
rect 28736 37284 28856 37312
rect 27709 37247 27767 37253
rect 27709 37213 27721 37247
rect 27755 37213 27767 37247
rect 27709 37207 27767 37213
rect 28537 37247 28595 37253
rect 28537 37213 28549 37247
rect 28583 37244 28595 37247
rect 28736 37244 28764 37284
rect 28583 37216 28764 37244
rect 28583 37213 28595 37216
rect 28537 37207 28595 37213
rect 28810 37204 28816 37256
rect 28868 37244 28874 37256
rect 28868 37216 28913 37244
rect 28868 37204 28874 37216
rect 28994 37204 29000 37256
rect 29052 37253 29058 37256
rect 29052 37247 29067 37253
rect 29055 37213 29067 37247
rect 29052 37207 29067 37213
rect 29052 37204 29058 37207
rect 27525 37179 27583 37185
rect 27525 37176 27537 37179
rect 24820 37148 26740 37176
rect 26804 37148 27537 37176
rect 24820 37136 24826 37148
rect 23687 37111 23745 37117
rect 23687 37108 23699 37111
rect 22848 37080 23699 37108
rect 23687 37077 23699 37080
rect 23733 37108 23745 37111
rect 24026 37108 24032 37120
rect 23733 37080 24032 37108
rect 23733 37077 23745 37080
rect 23687 37071 23745 37077
rect 24026 37068 24032 37080
rect 24084 37068 24090 37120
rect 24857 37111 24915 37117
rect 24857 37077 24869 37111
rect 24903 37108 24915 37111
rect 25590 37108 25596 37120
rect 24903 37080 25596 37108
rect 24903 37077 24915 37080
rect 24857 37071 24915 37077
rect 25590 37068 25596 37080
rect 25648 37108 25654 37120
rect 26804 37108 26832 37148
rect 27525 37145 27537 37148
rect 27571 37145 27583 37179
rect 27525 37139 27583 37145
rect 27614 37136 27620 37188
rect 27672 37176 27678 37188
rect 27672 37148 27765 37176
rect 27672 37136 27678 37148
rect 27798 37136 27804 37188
rect 27856 37176 27862 37188
rect 29549 37179 29607 37185
rect 29549 37176 29561 37179
rect 27856 37148 29561 37176
rect 27856 37136 27862 37148
rect 29549 37145 29561 37148
rect 29595 37145 29607 37179
rect 29549 37139 29607 37145
rect 30098 37136 30104 37188
rect 30156 37176 30162 37188
rect 32320 37176 33120 37190
rect 30156 37148 33120 37176
rect 30156 37136 30162 37148
rect 25648 37080 26832 37108
rect 25648 37068 25654 37080
rect 27154 37068 27160 37120
rect 27212 37108 27218 37120
rect 27632 37108 27660 37136
rect 32320 37134 33120 37148
rect 27212 37080 27660 37108
rect 28353 37111 28411 37117
rect 27212 37068 27218 37080
rect 28353 37077 28365 37111
rect 28399 37108 28411 37111
rect 28948 37108 28954 37120
rect 28399 37080 28954 37108
rect 28399 37077 28411 37080
rect 28353 37071 28411 37077
rect 28948 37068 28954 37080
rect 29006 37068 29012 37120
rect 29638 37068 29644 37120
rect 29696 37108 29702 37120
rect 30837 37111 30895 37117
rect 30837 37108 30849 37111
rect 29696 37080 30849 37108
rect 29696 37068 29702 37080
rect 30837 37077 30849 37080
rect 30883 37077 30895 37111
rect 30837 37071 30895 37077
rect 1104 37018 32016 37040
rect 1104 36966 7288 37018
rect 7340 36966 17592 37018
rect 17644 36966 27896 37018
rect 27948 36966 32016 37018
rect 1104 36944 32016 36966
rect 1397 36907 1455 36913
rect 1397 36873 1409 36907
rect 1443 36904 1455 36907
rect 1486 36904 1492 36916
rect 1443 36876 1492 36904
rect 1443 36873 1455 36876
rect 1397 36867 1455 36873
rect 1486 36864 1492 36876
rect 1544 36864 1550 36916
rect 3786 36904 3792 36916
rect 2516 36876 3792 36904
rect 2516 36777 2544 36876
rect 3786 36864 3792 36876
rect 3844 36864 3850 36916
rect 4338 36864 4344 36916
rect 4396 36904 4402 36916
rect 5261 36907 5319 36913
rect 5261 36904 5273 36907
rect 4396 36876 5273 36904
rect 4396 36864 4402 36876
rect 5261 36873 5273 36876
rect 5307 36873 5319 36907
rect 8021 36907 8079 36913
rect 8021 36904 8033 36907
rect 5261 36867 5319 36873
rect 6380 36876 8033 36904
rect 4985 36839 5043 36845
rect 4985 36836 4997 36839
rect 2792 36808 4108 36836
rect 2792 36777 2820 36808
rect 1581 36771 1639 36777
rect 1581 36737 1593 36771
rect 1627 36768 1639 36771
rect 2317 36771 2375 36777
rect 2317 36768 2329 36771
rect 1627 36740 2329 36768
rect 1627 36737 1639 36740
rect 1581 36731 1639 36737
rect 2317 36737 2329 36740
rect 2363 36737 2375 36771
rect 2317 36731 2375 36737
rect 2501 36771 2559 36777
rect 2501 36737 2513 36771
rect 2547 36737 2559 36771
rect 2501 36731 2559 36737
rect 2777 36771 2835 36777
rect 2777 36737 2789 36771
rect 2823 36737 2835 36771
rect 2777 36731 2835 36737
rect 2866 36728 2872 36780
rect 2924 36768 2930 36780
rect 2961 36771 3019 36777
rect 2961 36768 2973 36771
rect 2924 36740 2973 36768
rect 2924 36728 2930 36740
rect 2961 36737 2973 36740
rect 3007 36737 3019 36771
rect 3786 36768 3792 36780
rect 3747 36740 3792 36768
rect 2961 36731 3019 36737
rect 3786 36728 3792 36740
rect 3844 36728 3850 36780
rect 4080 36777 4108 36808
rect 4356 36808 4997 36836
rect 4356 36780 4384 36808
rect 4985 36805 4997 36808
rect 5031 36805 5043 36839
rect 4985 36799 5043 36805
rect 4065 36771 4123 36777
rect 4065 36737 4077 36771
rect 4111 36768 4123 36771
rect 4154 36768 4160 36780
rect 4111 36740 4160 36768
rect 4111 36737 4123 36740
rect 4065 36731 4123 36737
rect 4154 36728 4160 36740
rect 4212 36728 4218 36780
rect 4249 36771 4307 36777
rect 4249 36737 4261 36771
rect 4295 36768 4307 36771
rect 4338 36768 4344 36780
rect 4295 36740 4344 36768
rect 4295 36737 4307 36740
rect 4249 36731 4307 36737
rect 4338 36728 4344 36740
rect 4396 36728 4402 36780
rect 4614 36728 4620 36780
rect 4672 36768 4678 36780
rect 4709 36771 4767 36777
rect 4709 36768 4721 36771
rect 4672 36740 4721 36768
rect 4672 36728 4678 36740
rect 4709 36737 4721 36740
rect 4755 36737 4767 36771
rect 4709 36731 4767 36737
rect 4893 36771 4951 36777
rect 4893 36737 4905 36771
rect 4939 36737 4951 36771
rect 4893 36731 4951 36737
rect 5077 36771 5135 36777
rect 5077 36737 5089 36771
rect 5123 36768 5135 36771
rect 5626 36768 5632 36780
rect 5123 36740 5632 36768
rect 5123 36737 5135 36740
rect 5077 36731 5135 36737
rect 1857 36703 1915 36709
rect 1857 36669 1869 36703
rect 1903 36700 1915 36703
rect 3234 36700 3240 36712
rect 1903 36672 3240 36700
rect 1903 36669 1915 36672
rect 1857 36663 1915 36669
rect 3234 36660 3240 36672
rect 3292 36660 3298 36712
rect 4908 36700 4936 36731
rect 5626 36728 5632 36740
rect 5684 36728 5690 36780
rect 5350 36700 5356 36712
rect 4908 36672 5356 36700
rect 5350 36660 5356 36672
rect 5408 36700 5414 36712
rect 6380 36700 6408 36876
rect 8021 36873 8033 36876
rect 8067 36904 8079 36907
rect 8386 36904 8392 36916
rect 8067 36876 8392 36904
rect 8067 36873 8079 36876
rect 8021 36867 8079 36873
rect 8386 36864 8392 36876
rect 8444 36864 8450 36916
rect 9033 36907 9091 36913
rect 9033 36873 9045 36907
rect 9079 36904 9091 36907
rect 9079 36876 10272 36904
rect 9079 36873 9091 36876
rect 9033 36867 9091 36873
rect 6822 36796 6828 36848
rect 6880 36836 6886 36848
rect 9214 36836 9220 36848
rect 6880 36808 7144 36836
rect 6880 36796 6886 36808
rect 6546 36768 6552 36780
rect 6507 36740 6552 36768
rect 6546 36728 6552 36740
rect 6604 36728 6610 36780
rect 6822 36700 6828 36712
rect 5408 36672 6408 36700
rect 6783 36672 6828 36700
rect 5408 36660 5414 36672
rect 6822 36660 6828 36672
rect 6880 36660 6886 36712
rect 3326 36592 3332 36644
rect 3384 36632 3390 36644
rect 7006 36632 7012 36644
rect 3384 36604 7012 36632
rect 3384 36592 3390 36604
rect 7006 36592 7012 36604
rect 7064 36592 7070 36644
rect 7116 36632 7144 36808
rect 8036 36808 9220 36836
rect 8036 36777 8064 36808
rect 9214 36796 9220 36808
rect 9272 36836 9278 36848
rect 9769 36839 9827 36845
rect 9769 36836 9781 36839
rect 9272 36808 9781 36836
rect 9272 36796 9278 36808
rect 9769 36805 9781 36808
rect 9815 36805 9827 36839
rect 10244 36836 10272 36876
rect 10318 36864 10324 36916
rect 10376 36904 10382 36916
rect 11793 36907 11851 36913
rect 11793 36904 11805 36907
rect 10376 36876 11805 36904
rect 10376 36864 10382 36876
rect 11793 36873 11805 36876
rect 11839 36873 11851 36907
rect 11793 36867 11851 36873
rect 12250 36864 12256 36916
rect 12308 36904 12314 36916
rect 14366 36904 14372 36916
rect 12308 36876 14372 36904
rect 12308 36864 12314 36876
rect 14366 36864 14372 36876
rect 14424 36864 14430 36916
rect 14550 36864 14556 36916
rect 14608 36904 14614 36916
rect 14645 36907 14703 36913
rect 14645 36904 14657 36907
rect 14608 36876 14657 36904
rect 14608 36864 14614 36876
rect 14645 36873 14657 36876
rect 14691 36873 14703 36907
rect 15746 36904 15752 36916
rect 15707 36876 15752 36904
rect 14645 36867 14703 36873
rect 15746 36864 15752 36876
rect 15804 36864 15810 36916
rect 15838 36864 15844 36916
rect 15896 36904 15902 36916
rect 16853 36907 16911 36913
rect 15896 36876 15941 36904
rect 15896 36864 15902 36876
rect 16853 36873 16865 36907
rect 16899 36904 16911 36907
rect 18506 36904 18512 36916
rect 16899 36876 18512 36904
rect 16899 36873 16911 36876
rect 16853 36867 16911 36873
rect 18506 36864 18512 36876
rect 18564 36864 18570 36916
rect 18601 36907 18659 36913
rect 18601 36873 18613 36907
rect 18647 36904 18659 36907
rect 19058 36904 19064 36916
rect 18647 36876 19064 36904
rect 18647 36873 18659 36876
rect 18601 36867 18659 36873
rect 19058 36864 19064 36876
rect 19116 36864 19122 36916
rect 19705 36907 19763 36913
rect 19705 36873 19717 36907
rect 19751 36904 19763 36907
rect 19978 36904 19984 36916
rect 19751 36876 19984 36904
rect 19751 36873 19763 36876
rect 19705 36867 19763 36873
rect 19978 36864 19984 36876
rect 20036 36864 20042 36916
rect 20441 36907 20499 36913
rect 20441 36873 20453 36907
rect 20487 36904 20499 36907
rect 20898 36904 20904 36916
rect 20487 36876 20904 36904
rect 20487 36873 20499 36876
rect 20441 36867 20499 36873
rect 20898 36864 20904 36876
rect 20956 36904 20962 36916
rect 21174 36904 21180 36916
rect 20956 36876 21180 36904
rect 20956 36864 20962 36876
rect 21174 36864 21180 36876
rect 21232 36864 21238 36916
rect 27338 36904 27344 36916
rect 25516 36876 27344 36904
rect 11149 36839 11207 36845
rect 10244 36808 10548 36836
rect 9769 36799 9827 36805
rect 7837 36771 7895 36777
rect 7837 36737 7849 36771
rect 7883 36737 7895 36771
rect 7837 36731 7895 36737
rect 8021 36771 8079 36777
rect 8021 36737 8033 36771
rect 8067 36737 8079 36771
rect 8662 36768 8668 36780
rect 8623 36740 8668 36768
rect 8021 36731 8079 36737
rect 7852 36700 7880 36731
rect 8662 36728 8668 36740
rect 8720 36728 8726 36780
rect 8849 36771 8907 36777
rect 8849 36737 8861 36771
rect 8895 36768 8907 36771
rect 9033 36771 9091 36777
rect 9033 36768 9045 36771
rect 8895 36740 9045 36768
rect 8895 36737 8907 36740
rect 8849 36731 8907 36737
rect 9033 36737 9045 36740
rect 9079 36737 9091 36771
rect 9582 36768 9588 36780
rect 9543 36740 9588 36768
rect 9033 36731 9091 36737
rect 9582 36728 9588 36740
rect 9640 36728 9646 36780
rect 10520 36777 10548 36808
rect 11149 36805 11161 36839
rect 11195 36836 11207 36839
rect 11885 36839 11943 36845
rect 11885 36836 11897 36839
rect 11195 36808 11897 36836
rect 11195 36805 11207 36808
rect 11149 36799 11207 36805
rect 11885 36805 11897 36808
rect 11931 36805 11943 36839
rect 11885 36799 11943 36805
rect 12161 36839 12219 36845
rect 12161 36805 12173 36839
rect 12207 36836 12219 36839
rect 15286 36836 15292 36848
rect 12207 36808 15292 36836
rect 12207 36805 12219 36808
rect 12161 36799 12219 36805
rect 15286 36796 15292 36808
rect 15344 36796 15350 36848
rect 23109 36839 23167 36845
rect 23109 36836 23121 36839
rect 15672 36808 16988 36836
rect 10137 36771 10195 36777
rect 10137 36737 10149 36771
rect 10183 36768 10195 36771
rect 10229 36771 10287 36777
rect 10229 36768 10241 36771
rect 10183 36740 10241 36768
rect 10183 36737 10195 36740
rect 10137 36731 10195 36737
rect 10229 36737 10241 36740
rect 10275 36737 10287 36771
rect 10229 36731 10287 36737
rect 10505 36771 10563 36777
rect 10505 36737 10517 36771
rect 10551 36768 10563 36771
rect 11054 36768 11060 36780
rect 10551 36740 11060 36768
rect 10551 36737 10563 36740
rect 10505 36731 10563 36737
rect 11054 36728 11060 36740
rect 11112 36728 11118 36780
rect 11517 36771 11575 36777
rect 11517 36737 11529 36771
rect 11563 36768 11575 36771
rect 11606 36768 11612 36780
rect 11563 36740 11612 36768
rect 11563 36737 11575 36740
rect 11517 36731 11575 36737
rect 11606 36728 11612 36740
rect 11664 36728 11670 36780
rect 11701 36771 11759 36777
rect 11701 36737 11713 36771
rect 11747 36768 11759 36771
rect 11790 36768 11796 36780
rect 11747 36740 11796 36768
rect 11747 36737 11759 36740
rect 11701 36731 11759 36737
rect 11790 36728 11796 36740
rect 11848 36728 11854 36780
rect 12526 36728 12532 36780
rect 12584 36768 12590 36780
rect 12805 36771 12863 36777
rect 12805 36768 12817 36771
rect 12584 36740 12817 36768
rect 12584 36728 12590 36740
rect 12805 36737 12817 36740
rect 12851 36737 12863 36771
rect 13078 36768 13084 36780
rect 13039 36740 13084 36768
rect 12805 36731 12863 36737
rect 13078 36728 13084 36740
rect 13136 36728 13142 36780
rect 13262 36768 13268 36780
rect 13223 36740 13268 36768
rect 13262 36728 13268 36740
rect 13320 36768 13326 36780
rect 13320 36740 13400 36768
rect 13320 36728 13326 36740
rect 9122 36700 9128 36712
rect 7852 36672 9128 36700
rect 9122 36660 9128 36672
rect 9180 36660 9186 36712
rect 9306 36660 9312 36712
rect 9364 36700 9370 36712
rect 9401 36703 9459 36709
rect 9401 36700 9413 36703
rect 9364 36672 9413 36700
rect 9364 36660 9370 36672
rect 9401 36669 9413 36672
rect 9447 36700 9459 36703
rect 13372 36700 13400 36740
rect 13446 36728 13452 36780
rect 13504 36768 13510 36780
rect 14093 36771 14151 36777
rect 14093 36768 14105 36771
rect 13504 36740 14105 36768
rect 13504 36728 13510 36740
rect 14093 36737 14105 36740
rect 14139 36737 14151 36771
rect 14274 36768 14280 36780
rect 14235 36740 14280 36768
rect 14093 36731 14151 36737
rect 14274 36728 14280 36740
rect 14332 36728 14338 36780
rect 14369 36771 14427 36777
rect 14369 36737 14381 36771
rect 14415 36737 14427 36771
rect 14369 36731 14427 36737
rect 14384 36700 14412 36731
rect 14458 36728 14464 36780
rect 14516 36768 14522 36780
rect 14918 36768 14924 36780
rect 14516 36740 14924 36768
rect 14516 36728 14522 36740
rect 14918 36728 14924 36740
rect 14976 36768 14982 36780
rect 15672 36768 15700 36808
rect 16960 36780 16988 36808
rect 17236 36808 23121 36836
rect 16666 36768 16672 36780
rect 14976 36740 15700 36768
rect 16627 36740 16672 36768
rect 14976 36728 14982 36740
rect 16666 36728 16672 36740
rect 16724 36728 16730 36780
rect 16942 36768 16948 36780
rect 16903 36740 16948 36768
rect 16942 36728 16948 36740
rect 17000 36728 17006 36780
rect 9447 36672 12434 36700
rect 13372 36672 14412 36700
rect 9447 36669 9459 36672
rect 9401 36663 9459 36669
rect 8849 36635 8907 36641
rect 8849 36632 8861 36635
rect 7116 36604 8861 36632
rect 8849 36601 8861 36604
rect 8895 36601 8907 36635
rect 9140 36632 9168 36660
rect 10137 36635 10195 36641
rect 10137 36632 10149 36635
rect 9140 36604 10149 36632
rect 8849 36595 8907 36601
rect 10137 36601 10149 36604
rect 10183 36601 10195 36635
rect 10137 36595 10195 36601
rect 10226 36592 10232 36644
rect 10284 36632 10290 36644
rect 10505 36635 10563 36641
rect 10505 36632 10517 36635
rect 10284 36604 10517 36632
rect 10284 36592 10290 36604
rect 10505 36601 10517 36604
rect 10551 36601 10563 36635
rect 12406 36632 12434 36672
rect 14550 36660 14556 36712
rect 14608 36700 14614 36712
rect 15654 36700 15660 36712
rect 14608 36672 15660 36700
rect 14608 36660 14614 36672
rect 15654 36660 15660 36672
rect 15712 36660 15718 36712
rect 16025 36703 16083 36709
rect 16025 36669 16037 36703
rect 16071 36700 16083 36703
rect 17034 36700 17040 36712
rect 16071 36672 17040 36700
rect 16071 36669 16083 36672
rect 16025 36663 16083 36669
rect 17034 36660 17040 36672
rect 17092 36660 17098 36712
rect 17236 36632 17264 36808
rect 23109 36805 23121 36808
rect 23155 36836 23167 36839
rect 23382 36836 23388 36848
rect 23155 36808 23388 36836
rect 23155 36805 23167 36808
rect 23109 36799 23167 36805
rect 23382 36796 23388 36808
rect 23440 36796 23446 36848
rect 17589 36771 17647 36777
rect 17589 36737 17601 36771
rect 17635 36768 17647 36771
rect 17770 36768 17776 36780
rect 17635 36740 17776 36768
rect 17635 36737 17647 36740
rect 17589 36731 17647 36737
rect 17770 36728 17776 36740
rect 17828 36728 17834 36780
rect 18785 36771 18843 36777
rect 18785 36768 18797 36771
rect 18156 36740 18797 36768
rect 17494 36660 17500 36712
rect 17552 36700 17558 36712
rect 17865 36703 17923 36709
rect 17865 36700 17877 36703
rect 17552 36672 17877 36700
rect 17552 36660 17558 36672
rect 17865 36669 17877 36672
rect 17911 36700 17923 36703
rect 18046 36700 18052 36712
rect 17911 36672 18052 36700
rect 17911 36669 17923 36672
rect 17865 36663 17923 36669
rect 18046 36660 18052 36672
rect 18104 36660 18110 36712
rect 12406 36604 17264 36632
rect 10505 36595 10563 36601
rect 17678 36592 17684 36644
rect 17736 36632 17742 36644
rect 18156 36632 18184 36740
rect 18785 36737 18797 36740
rect 18831 36737 18843 36771
rect 18785 36731 18843 36737
rect 19061 36771 19119 36777
rect 19061 36737 19073 36771
rect 19107 36737 19119 36771
rect 19242 36768 19248 36780
rect 19203 36740 19248 36768
rect 19061 36731 19119 36737
rect 18230 36660 18236 36712
rect 18288 36700 18294 36712
rect 19076 36700 19104 36731
rect 19242 36728 19248 36740
rect 19300 36728 19306 36780
rect 19518 36728 19524 36780
rect 19576 36768 19582 36780
rect 19889 36771 19947 36777
rect 19889 36768 19901 36771
rect 19576 36740 19901 36768
rect 19576 36728 19582 36740
rect 19889 36737 19901 36740
rect 19935 36737 19947 36771
rect 19889 36731 19947 36737
rect 20165 36771 20223 36777
rect 20165 36737 20177 36771
rect 20211 36737 20223 36771
rect 20165 36731 20223 36737
rect 20349 36771 20407 36777
rect 20349 36737 20361 36771
rect 20395 36768 20407 36771
rect 20441 36771 20499 36777
rect 20441 36768 20453 36771
rect 20395 36740 20453 36768
rect 20395 36737 20407 36740
rect 20349 36731 20407 36737
rect 20441 36737 20453 36740
rect 20487 36737 20499 36771
rect 20441 36731 20499 36737
rect 20903 36771 20961 36777
rect 20903 36737 20915 36771
rect 20949 36737 20961 36771
rect 20903 36731 20961 36737
rect 20180 36700 20208 36731
rect 18288 36672 20208 36700
rect 20916 36700 20944 36731
rect 21174 36728 21180 36780
rect 21232 36768 21238 36780
rect 21821 36771 21879 36777
rect 21821 36768 21833 36771
rect 21232 36740 21833 36768
rect 21232 36728 21238 36740
rect 21821 36737 21833 36740
rect 21867 36737 21879 36771
rect 21821 36731 21879 36737
rect 22646 36728 22652 36780
rect 22704 36768 22710 36780
rect 22925 36771 22983 36777
rect 22925 36768 22937 36771
rect 22704 36740 22937 36768
rect 22704 36728 22710 36740
rect 22925 36737 22937 36740
rect 22971 36768 22983 36771
rect 23014 36768 23020 36780
rect 22971 36740 23020 36768
rect 22971 36737 22983 36740
rect 22925 36731 22983 36737
rect 23014 36728 23020 36740
rect 23072 36728 23078 36780
rect 23400 36768 23428 36796
rect 24121 36771 24179 36777
rect 24121 36768 24133 36771
rect 23400 36740 24133 36768
rect 24121 36737 24133 36740
rect 24167 36737 24179 36771
rect 25222 36768 25228 36780
rect 25183 36740 25228 36768
rect 24121 36731 24179 36737
rect 25222 36728 25228 36740
rect 25280 36728 25286 36780
rect 25516 36777 25544 36876
rect 27338 36864 27344 36876
rect 27396 36864 27402 36916
rect 28810 36864 28816 36916
rect 28868 36904 28874 36916
rect 30193 36907 30251 36913
rect 28868 36876 30052 36904
rect 28868 36864 28874 36876
rect 30024 36848 30052 36876
rect 30193 36873 30205 36907
rect 30239 36904 30251 36907
rect 30282 36904 30288 36916
rect 30239 36876 30288 36904
rect 30239 36873 30251 36876
rect 30193 36867 30251 36873
rect 30282 36864 30288 36876
rect 30340 36864 30346 36916
rect 28994 36836 29000 36848
rect 27264 36808 29000 36836
rect 25501 36771 25559 36777
rect 25501 36737 25513 36771
rect 25547 36737 25559 36771
rect 26142 36768 26148 36780
rect 26103 36740 26148 36768
rect 25501 36731 25559 36737
rect 26142 36728 26148 36740
rect 26200 36728 26206 36780
rect 26421 36771 26479 36777
rect 26421 36737 26433 36771
rect 26467 36768 26479 36771
rect 27154 36768 27160 36780
rect 26467 36740 27160 36768
rect 26467 36737 26479 36740
rect 26421 36731 26479 36737
rect 27154 36728 27160 36740
rect 27212 36728 27218 36780
rect 27264 36777 27292 36808
rect 28994 36796 29000 36808
rect 29052 36796 29058 36848
rect 30006 36796 30012 36848
rect 30064 36836 30070 36848
rect 30064 36808 30696 36836
rect 30064 36796 30070 36808
rect 27249 36771 27307 36777
rect 27249 36737 27261 36771
rect 27295 36737 27307 36771
rect 27505 36771 27563 36777
rect 27505 36768 27517 36771
rect 27249 36731 27307 36737
rect 27356 36740 27517 36768
rect 22370 36700 22376 36712
rect 20916 36672 22376 36700
rect 18288 36660 18294 36672
rect 22370 36660 22376 36672
rect 22428 36660 22434 36712
rect 24026 36660 24032 36712
rect 24084 36700 24090 36712
rect 26786 36700 26792 36712
rect 24084 36672 26792 36700
rect 24084 36660 24090 36672
rect 26786 36660 26792 36672
rect 26844 36660 26850 36712
rect 27356 36700 27384 36740
rect 27505 36737 27517 36740
rect 27551 36737 27563 36771
rect 29270 36768 29276 36780
rect 29231 36740 29276 36768
rect 27505 36731 27563 36737
rect 29270 36728 29276 36740
rect 29328 36728 29334 36780
rect 29730 36728 29736 36780
rect 29788 36768 29794 36780
rect 30668 36777 30696 36808
rect 30377 36771 30435 36777
rect 30377 36768 30389 36771
rect 29788 36740 30389 36768
rect 29788 36728 29794 36740
rect 30377 36737 30389 36740
rect 30423 36737 30435 36771
rect 30377 36731 30435 36737
rect 30653 36771 30711 36777
rect 30653 36737 30665 36771
rect 30699 36737 30711 36771
rect 30653 36731 30711 36737
rect 30837 36771 30895 36777
rect 30837 36737 30849 36771
rect 30883 36768 30895 36771
rect 31294 36768 31300 36780
rect 30883 36740 31300 36768
rect 30883 36737 30895 36740
rect 30837 36731 30895 36737
rect 29549 36703 29607 36709
rect 29549 36700 29561 36703
rect 27264 36672 27384 36700
rect 28552 36672 29561 36700
rect 17736 36604 18184 36632
rect 18509 36635 18567 36641
rect 17736 36592 17742 36604
rect 18509 36601 18521 36635
rect 18555 36632 18567 36635
rect 19242 36632 19248 36644
rect 18555 36604 19248 36632
rect 18555 36601 18567 36604
rect 18509 36595 18567 36601
rect 19242 36592 19248 36604
rect 19300 36592 19306 36644
rect 21358 36592 21364 36644
rect 21416 36632 21422 36644
rect 22281 36635 22339 36641
rect 22281 36632 22293 36635
rect 21416 36604 22293 36632
rect 21416 36592 21422 36604
rect 22281 36601 22293 36604
rect 22327 36601 22339 36635
rect 22281 36595 22339 36601
rect 24305 36635 24363 36641
rect 24305 36601 24317 36635
rect 24351 36632 24363 36635
rect 25590 36632 25596 36644
rect 24351 36604 25596 36632
rect 24351 36601 24363 36604
rect 24305 36595 24363 36601
rect 25590 36592 25596 36604
rect 25648 36592 25654 36644
rect 25961 36635 26019 36641
rect 25961 36601 25973 36635
rect 26007 36632 26019 36635
rect 27264 36632 27292 36672
rect 26007 36604 27292 36632
rect 26007 36601 26019 36604
rect 25961 36595 26019 36601
rect 1765 36567 1823 36573
rect 1765 36533 1777 36567
rect 1811 36564 1823 36567
rect 2222 36564 2228 36576
rect 1811 36536 2228 36564
rect 1811 36533 1823 36536
rect 1765 36527 1823 36533
rect 2222 36524 2228 36536
rect 2280 36524 2286 36576
rect 2406 36524 2412 36576
rect 2464 36564 2470 36576
rect 3605 36567 3663 36573
rect 3605 36564 3617 36567
rect 2464 36536 3617 36564
rect 2464 36524 2470 36536
rect 3605 36533 3617 36536
rect 3651 36533 3663 36567
rect 6362 36564 6368 36576
rect 6323 36536 6368 36564
rect 3605 36527 3663 36533
rect 6362 36524 6368 36536
rect 6420 36524 6426 36576
rect 6733 36567 6791 36573
rect 6733 36533 6745 36567
rect 6779 36564 6791 36567
rect 8110 36564 8116 36576
rect 6779 36536 8116 36564
rect 6779 36533 6791 36536
rect 6733 36527 6791 36533
rect 8110 36524 8116 36536
rect 8168 36524 8174 36576
rect 8386 36524 8392 36576
rect 8444 36564 8450 36576
rect 11149 36567 11207 36573
rect 11149 36564 11161 36567
rect 8444 36536 11161 36564
rect 8444 36524 8450 36536
rect 11149 36533 11161 36536
rect 11195 36533 11207 36567
rect 11149 36527 11207 36533
rect 11698 36524 11704 36576
rect 11756 36564 11762 36576
rect 12069 36567 12127 36573
rect 12069 36564 12081 36567
rect 11756 36536 12081 36564
rect 11756 36524 11762 36536
rect 12069 36533 12081 36536
rect 12115 36564 12127 36567
rect 12161 36567 12219 36573
rect 12161 36564 12173 36567
rect 12115 36536 12173 36564
rect 12115 36533 12127 36536
rect 12069 36527 12127 36533
rect 12161 36533 12173 36536
rect 12207 36533 12219 36567
rect 12161 36527 12219 36533
rect 12621 36567 12679 36573
rect 12621 36533 12633 36567
rect 12667 36564 12679 36567
rect 13538 36564 13544 36576
rect 12667 36536 13544 36564
rect 12667 36533 12679 36536
rect 12621 36527 12679 36533
rect 13538 36524 13544 36536
rect 13596 36524 13602 36576
rect 15378 36564 15384 36576
rect 15339 36536 15384 36564
rect 15378 36524 15384 36536
rect 15436 36524 15442 36576
rect 15746 36524 15752 36576
rect 15804 36564 15810 36576
rect 16669 36567 16727 36573
rect 16669 36564 16681 36567
rect 15804 36536 16681 36564
rect 15804 36524 15810 36536
rect 16669 36533 16681 36536
rect 16715 36533 16727 36567
rect 17402 36564 17408 36576
rect 17363 36536 17408 36564
rect 16669 36527 16727 36533
rect 17402 36524 17408 36536
rect 17460 36524 17466 36576
rect 17773 36567 17831 36573
rect 17773 36533 17785 36567
rect 17819 36564 17831 36567
rect 19150 36564 19156 36576
rect 17819 36536 19156 36564
rect 17819 36533 17831 36536
rect 17773 36527 17831 36533
rect 19150 36524 19156 36536
rect 19208 36524 19214 36576
rect 19702 36524 19708 36576
rect 19760 36564 19766 36576
rect 20993 36567 21051 36573
rect 20993 36564 21005 36567
rect 19760 36536 21005 36564
rect 19760 36524 19766 36536
rect 20993 36533 21005 36536
rect 21039 36533 21051 36567
rect 20993 36527 21051 36533
rect 21174 36524 21180 36576
rect 21232 36564 21238 36576
rect 21910 36564 21916 36576
rect 21232 36536 21916 36564
rect 21232 36524 21238 36536
rect 21910 36524 21916 36536
rect 21968 36524 21974 36576
rect 24670 36524 24676 36576
rect 24728 36564 24734 36576
rect 25041 36567 25099 36573
rect 25041 36564 25053 36567
rect 24728 36536 25053 36564
rect 24728 36524 24734 36536
rect 25041 36533 25053 36536
rect 25087 36533 25099 36567
rect 25041 36527 25099 36533
rect 25409 36567 25467 36573
rect 25409 36533 25421 36567
rect 25455 36564 25467 36567
rect 26050 36564 26056 36576
rect 25455 36536 26056 36564
rect 25455 36533 25467 36536
rect 25409 36527 25467 36533
rect 26050 36524 26056 36536
rect 26108 36524 26114 36576
rect 26329 36567 26387 36573
rect 26329 36533 26341 36567
rect 26375 36564 26387 36567
rect 26786 36564 26792 36576
rect 26375 36536 26792 36564
rect 26375 36533 26387 36536
rect 26329 36527 26387 36533
rect 26786 36524 26792 36536
rect 26844 36524 26850 36576
rect 27430 36524 27436 36576
rect 27488 36564 27494 36576
rect 28552 36564 28580 36672
rect 29549 36669 29561 36672
rect 29595 36700 29607 36703
rect 30852 36700 30880 36731
rect 31294 36728 31300 36740
rect 31352 36728 31358 36780
rect 29595 36672 30880 36700
rect 29595 36669 29607 36672
rect 29549 36663 29607 36669
rect 28902 36592 28908 36644
rect 28960 36632 28966 36644
rect 29457 36635 29515 36641
rect 29457 36632 29469 36635
rect 28960 36604 29469 36632
rect 28960 36592 28966 36604
rect 29457 36601 29469 36604
rect 29503 36632 29515 36635
rect 31018 36632 31024 36644
rect 29503 36604 31024 36632
rect 29503 36601 29515 36604
rect 29457 36595 29515 36601
rect 31018 36592 31024 36604
rect 31076 36592 31082 36644
rect 27488 36536 28580 36564
rect 27488 36524 27494 36536
rect 28626 36524 28632 36576
rect 28684 36564 28690 36576
rect 29089 36567 29147 36573
rect 28684 36536 28729 36564
rect 28684 36524 28690 36536
rect 29089 36533 29101 36567
rect 29135 36564 29147 36567
rect 29546 36564 29552 36576
rect 29135 36536 29552 36564
rect 29135 36533 29147 36536
rect 29089 36527 29147 36533
rect 29546 36524 29552 36536
rect 29604 36524 29610 36576
rect 1104 36474 32016 36496
rect 1104 36422 2136 36474
rect 2188 36422 12440 36474
rect 12492 36422 22744 36474
rect 22796 36422 32016 36474
rect 1104 36400 32016 36422
rect 2498 36320 2504 36372
rect 2556 36360 2562 36372
rect 4614 36360 4620 36372
rect 2556 36332 4620 36360
rect 2556 36320 2562 36332
rect 4614 36320 4620 36332
rect 4672 36320 4678 36372
rect 6270 36320 6276 36372
rect 6328 36360 6334 36372
rect 7929 36363 7987 36369
rect 6328 36332 7328 36360
rect 6328 36320 6334 36332
rect 1581 36295 1639 36301
rect 1581 36261 1593 36295
rect 1627 36292 1639 36295
rect 2590 36292 2596 36304
rect 1627 36264 2596 36292
rect 1627 36261 1639 36264
rect 1581 36255 1639 36261
rect 2590 36252 2596 36264
rect 2648 36252 2654 36304
rect 2792 36196 4200 36224
rect 2792 36165 2820 36196
rect 4172 36168 4200 36196
rect 5442 36184 5448 36236
rect 5500 36224 5506 36236
rect 5537 36227 5595 36233
rect 5537 36224 5549 36227
rect 5500 36196 5549 36224
rect 5500 36184 5506 36196
rect 5537 36193 5549 36196
rect 5583 36193 5595 36227
rect 7300 36224 7328 36332
rect 7929 36329 7941 36363
rect 7975 36360 7987 36363
rect 8021 36363 8079 36369
rect 8021 36360 8033 36363
rect 7975 36332 8033 36360
rect 7975 36329 7987 36332
rect 7929 36323 7987 36329
rect 8021 36329 8033 36332
rect 8067 36329 8079 36363
rect 8386 36360 8392 36372
rect 8347 36332 8392 36360
rect 8021 36323 8079 36329
rect 8386 36320 8392 36332
rect 8444 36320 8450 36372
rect 9122 36320 9128 36372
rect 9180 36360 9186 36372
rect 9677 36363 9735 36369
rect 9677 36360 9689 36363
rect 9180 36332 9689 36360
rect 9180 36320 9186 36332
rect 9677 36329 9689 36332
rect 9723 36329 9735 36363
rect 9677 36323 9735 36329
rect 10318 36320 10324 36372
rect 10376 36360 10382 36372
rect 10686 36360 10692 36372
rect 10376 36332 10692 36360
rect 10376 36320 10382 36332
rect 10686 36320 10692 36332
rect 10744 36320 10750 36372
rect 10778 36320 10784 36372
rect 10836 36360 10842 36372
rect 10873 36363 10931 36369
rect 10873 36360 10885 36363
rect 10836 36332 10885 36360
rect 10836 36320 10842 36332
rect 10873 36329 10885 36332
rect 10919 36329 10931 36363
rect 10873 36323 10931 36329
rect 11054 36320 11060 36372
rect 11112 36360 11118 36372
rect 11517 36363 11575 36369
rect 11517 36360 11529 36363
rect 11112 36332 11529 36360
rect 11112 36320 11118 36332
rect 11517 36329 11529 36332
rect 11563 36329 11575 36363
rect 22186 36360 22192 36372
rect 11517 36323 11575 36329
rect 11716 36332 22192 36360
rect 7377 36295 7435 36301
rect 7377 36261 7389 36295
rect 7423 36292 7435 36295
rect 11606 36292 11612 36304
rect 7423 36264 11612 36292
rect 7423 36261 7435 36264
rect 7377 36255 7435 36261
rect 11606 36252 11612 36264
rect 11664 36252 11670 36304
rect 9306 36224 9312 36236
rect 7300 36196 8064 36224
rect 9267 36196 9312 36224
rect 5537 36187 5595 36193
rect 1397 36159 1455 36165
rect 1397 36125 1409 36159
rect 1443 36125 1455 36159
rect 1397 36119 1455 36125
rect 2501 36159 2559 36165
rect 2501 36125 2513 36159
rect 2547 36125 2559 36159
rect 2501 36119 2559 36125
rect 2777 36159 2835 36165
rect 2777 36125 2789 36159
rect 2823 36125 2835 36159
rect 2777 36119 2835 36125
rect 2961 36159 3019 36165
rect 2961 36125 2973 36159
rect 3007 36156 3019 36159
rect 3234 36156 3240 36168
rect 3007 36128 3240 36156
rect 3007 36125 3019 36128
rect 2961 36119 3019 36125
rect 1412 36020 1440 36119
rect 2516 36088 2544 36119
rect 3234 36116 3240 36128
rect 3292 36116 3298 36168
rect 3786 36116 3792 36168
rect 3844 36156 3850 36168
rect 3973 36159 4031 36165
rect 3973 36156 3985 36159
rect 3844 36128 3985 36156
rect 3844 36116 3850 36128
rect 3973 36125 3985 36128
rect 4019 36125 4031 36159
rect 3973 36119 4031 36125
rect 4154 36116 4160 36168
rect 4212 36156 4218 36168
rect 4249 36159 4307 36165
rect 4249 36156 4261 36159
rect 4212 36128 4261 36156
rect 4212 36116 4218 36128
rect 4249 36125 4261 36128
rect 4295 36125 4307 36159
rect 4249 36119 4307 36125
rect 4433 36159 4491 36165
rect 4433 36125 4445 36159
rect 4479 36156 4491 36159
rect 4706 36156 4712 36168
rect 4479 36128 4712 36156
rect 4479 36125 4491 36128
rect 4433 36119 4491 36125
rect 4706 36116 4712 36128
rect 4764 36156 4770 36168
rect 5166 36156 5172 36168
rect 4764 36128 5172 36156
rect 4764 36116 4770 36128
rect 5166 36116 5172 36128
rect 5224 36116 5230 36168
rect 5804 36159 5862 36165
rect 5804 36125 5816 36159
rect 5850 36156 5862 36159
rect 6638 36156 6644 36168
rect 5850 36128 6644 36156
rect 5850 36125 5862 36128
rect 5804 36119 5862 36125
rect 6638 36116 6644 36128
rect 6696 36116 6702 36168
rect 8036 36165 8064 36196
rect 9306 36184 9312 36196
rect 9364 36184 9370 36236
rect 9582 36184 9588 36236
rect 9640 36224 9646 36236
rect 10962 36224 10968 36236
rect 9640 36196 10824 36224
rect 10923 36196 10968 36224
rect 9640 36184 9646 36196
rect 7561 36159 7619 36165
rect 7561 36125 7573 36159
rect 7607 36125 7619 36159
rect 7561 36119 7619 36125
rect 8021 36159 8079 36165
rect 8021 36125 8033 36159
rect 8067 36125 8079 36159
rect 8021 36119 8079 36125
rect 8205 36159 8263 36165
rect 8205 36125 8217 36159
rect 8251 36156 8263 36159
rect 9398 36156 9404 36168
rect 8251 36128 9404 36156
rect 8251 36125 8263 36128
rect 8205 36119 8263 36125
rect 3804 36088 3832 36116
rect 2516 36060 3832 36088
rect 7576 36088 7604 36119
rect 9398 36116 9404 36128
rect 9456 36116 9462 36168
rect 9493 36159 9551 36165
rect 9493 36125 9505 36159
rect 9539 36156 9551 36159
rect 9674 36156 9680 36168
rect 9539 36128 9680 36156
rect 9539 36125 9551 36128
rect 9493 36119 9551 36125
rect 9674 36116 9680 36128
rect 9732 36116 9738 36168
rect 10686 36156 10692 36168
rect 10647 36128 10692 36156
rect 10686 36116 10692 36128
rect 10744 36116 10750 36168
rect 10796 36156 10824 36196
rect 10962 36184 10968 36196
rect 11020 36184 11026 36236
rect 11422 36156 11428 36168
rect 10796 36128 11428 36156
rect 11422 36116 11428 36128
rect 11480 36116 11486 36168
rect 11609 36159 11667 36165
rect 11609 36125 11621 36159
rect 11655 36156 11667 36159
rect 11716 36156 11744 36332
rect 22186 36320 22192 36332
rect 22244 36320 22250 36372
rect 23661 36363 23719 36369
rect 23661 36329 23673 36363
rect 23707 36360 23719 36363
rect 24762 36360 24768 36372
rect 23707 36332 24768 36360
rect 23707 36329 23719 36332
rect 23661 36323 23719 36329
rect 24762 36320 24768 36332
rect 24820 36320 24826 36372
rect 26142 36320 26148 36372
rect 26200 36360 26206 36372
rect 27617 36363 27675 36369
rect 27617 36360 27629 36363
rect 26200 36332 27629 36360
rect 26200 36320 26206 36332
rect 27617 36329 27629 36332
rect 27663 36329 27675 36363
rect 28902 36360 28908 36372
rect 27617 36323 27675 36329
rect 27724 36332 28908 36360
rect 13262 36252 13268 36304
rect 13320 36292 13326 36304
rect 13541 36295 13599 36301
rect 13541 36292 13553 36295
rect 13320 36264 13553 36292
rect 13320 36252 13326 36264
rect 13541 36261 13553 36264
rect 13587 36261 13599 36295
rect 13541 36255 13599 36261
rect 14274 36252 14280 36304
rect 14332 36292 14338 36304
rect 14829 36295 14887 36301
rect 14829 36292 14841 36295
rect 14332 36264 14841 36292
rect 14332 36252 14338 36264
rect 14829 36261 14841 36264
rect 14875 36261 14887 36295
rect 14829 36255 14887 36261
rect 15194 36252 15200 36304
rect 15252 36292 15258 36304
rect 16485 36295 16543 36301
rect 15252 36264 16344 36292
rect 15252 36252 15258 36264
rect 16316 36224 16344 36264
rect 16485 36261 16497 36295
rect 16531 36292 16543 36295
rect 16666 36292 16672 36304
rect 16531 36264 16672 36292
rect 16531 36261 16543 36264
rect 16485 36255 16543 36261
rect 16666 36252 16672 36264
rect 16724 36252 16730 36304
rect 17770 36292 17776 36304
rect 17731 36264 17776 36292
rect 17770 36252 17776 36264
rect 17828 36252 17834 36304
rect 27157 36295 27215 36301
rect 27157 36261 27169 36295
rect 27203 36292 27215 36295
rect 27338 36292 27344 36304
rect 27203 36264 27344 36292
rect 27203 36261 27215 36264
rect 27157 36255 27215 36261
rect 27338 36252 27344 36264
rect 27396 36252 27402 36304
rect 17494 36224 17500 36236
rect 16316 36196 16712 36224
rect 11655 36128 11744 36156
rect 12161 36159 12219 36165
rect 11655 36125 11667 36128
rect 11609 36119 11667 36125
rect 12161 36125 12173 36159
rect 12207 36156 12219 36159
rect 13170 36156 13176 36168
rect 12207 36128 13176 36156
rect 12207 36125 12219 36128
rect 12161 36119 12219 36125
rect 7576 36060 11008 36088
rect 1044 35992 1440 36020
rect 1044 35748 1072 35992
rect 2038 35980 2044 36032
rect 2096 36020 2102 36032
rect 2317 36023 2375 36029
rect 2317 36020 2329 36023
rect 2096 35992 2329 36020
rect 2096 35980 2102 35992
rect 2317 35989 2329 35992
rect 2363 35989 2375 36023
rect 2317 35983 2375 35989
rect 2958 35980 2964 36032
rect 3016 36020 3022 36032
rect 3789 36023 3847 36029
rect 3789 36020 3801 36023
rect 3016 35992 3801 36020
rect 3016 35980 3022 35992
rect 3789 35989 3801 35992
rect 3835 35989 3847 36023
rect 3789 35983 3847 35989
rect 4614 35980 4620 36032
rect 4672 36020 4678 36032
rect 6917 36023 6975 36029
rect 6917 36020 6929 36023
rect 4672 35992 6929 36020
rect 4672 35980 4678 35992
rect 6917 35989 6929 35992
rect 6963 36020 6975 36023
rect 7006 36020 7012 36032
rect 6963 35992 7012 36020
rect 6963 35989 6975 35992
rect 6917 35983 6975 35989
rect 7006 35980 7012 35992
rect 7064 35980 7070 36032
rect 7929 36023 7987 36029
rect 7929 35989 7941 36023
rect 7975 36020 7987 36023
rect 10318 36020 10324 36032
rect 7975 35992 10324 36020
rect 7975 35989 7987 35992
rect 7929 35983 7987 35989
rect 10318 35980 10324 35992
rect 10376 35980 10382 36032
rect 10502 36020 10508 36032
rect 10463 35992 10508 36020
rect 10502 35980 10508 35992
rect 10560 35980 10566 36032
rect 10980 36020 11008 36060
rect 11054 36048 11060 36100
rect 11112 36088 11118 36100
rect 11624 36088 11652 36119
rect 13170 36116 13176 36128
rect 13228 36156 13234 36168
rect 13998 36156 14004 36168
rect 13228 36128 14004 36156
rect 13228 36116 13234 36128
rect 13998 36116 14004 36128
rect 14056 36116 14062 36168
rect 14550 36156 14556 36168
rect 14511 36128 14556 36156
rect 14550 36116 14556 36128
rect 14608 36116 14614 36168
rect 14642 36116 14648 36168
rect 14700 36156 14706 36168
rect 14737 36159 14795 36165
rect 14737 36156 14749 36159
rect 14700 36128 14749 36156
rect 14700 36116 14706 36128
rect 14737 36125 14749 36128
rect 14783 36125 14795 36159
rect 15746 36156 15752 36168
rect 15707 36128 15752 36156
rect 14737 36119 14795 36125
rect 15746 36116 15752 36128
rect 15804 36116 15810 36168
rect 16025 36159 16083 36165
rect 16025 36125 16037 36159
rect 16071 36156 16083 36159
rect 16574 36156 16580 36168
rect 16071 36128 16580 36156
rect 16071 36125 16083 36128
rect 16025 36119 16083 36125
rect 16574 36116 16580 36128
rect 16632 36116 16638 36168
rect 16684 36165 16712 36196
rect 16776 36196 17500 36224
rect 16776 36165 16804 36196
rect 17494 36184 17500 36196
rect 17552 36184 17558 36236
rect 19518 36224 19524 36236
rect 18064 36196 19524 36224
rect 16669 36159 16727 36165
rect 16669 36125 16681 36159
rect 16715 36125 16727 36159
rect 16669 36119 16727 36125
rect 16761 36159 16819 36165
rect 16761 36125 16773 36159
rect 16807 36125 16819 36159
rect 16942 36156 16948 36168
rect 16903 36128 16948 36156
rect 16761 36119 16819 36125
rect 16942 36116 16948 36128
rect 17000 36116 17006 36168
rect 17034 36116 17040 36168
rect 17092 36156 17098 36168
rect 17092 36128 17137 36156
rect 17092 36116 17098 36128
rect 17862 36116 17868 36168
rect 17920 36156 17926 36168
rect 17957 36159 18015 36165
rect 17957 36156 17969 36159
rect 17920 36128 17969 36156
rect 17920 36116 17926 36128
rect 17957 36125 17969 36128
rect 18003 36156 18015 36159
rect 18064 36156 18092 36196
rect 19518 36184 19524 36196
rect 19576 36184 19582 36236
rect 22664 36196 23796 36224
rect 18230 36156 18236 36168
rect 18003 36128 18092 36156
rect 18191 36128 18236 36156
rect 18003 36125 18015 36128
rect 17957 36119 18015 36125
rect 18230 36116 18236 36128
rect 18288 36116 18294 36168
rect 18322 36116 18328 36168
rect 18380 36156 18386 36168
rect 18417 36159 18475 36165
rect 18417 36156 18429 36159
rect 18380 36128 18429 36156
rect 18380 36116 18386 36128
rect 18417 36125 18429 36128
rect 18463 36125 18475 36159
rect 18417 36119 18475 36125
rect 19429 36159 19487 36165
rect 19429 36125 19441 36159
rect 19475 36156 19487 36159
rect 19536 36156 19564 36184
rect 22664 36168 22692 36196
rect 19475 36128 19564 36156
rect 19705 36159 19763 36165
rect 19475 36125 19487 36128
rect 19429 36119 19487 36125
rect 19705 36125 19717 36159
rect 19751 36125 19763 36159
rect 19705 36119 19763 36125
rect 19889 36159 19947 36165
rect 19889 36125 19901 36159
rect 19935 36156 19947 36159
rect 19978 36156 19984 36168
rect 19935 36128 19984 36156
rect 19935 36125 19947 36128
rect 19889 36119 19947 36125
rect 11112 36060 11652 36088
rect 12428 36091 12486 36097
rect 11112 36048 11118 36060
rect 12428 36057 12440 36091
rect 12474 36088 12486 36091
rect 13354 36088 13360 36100
rect 12474 36060 13360 36088
rect 12474 36057 12486 36060
rect 12428 36051 12486 36057
rect 13354 36048 13360 36060
rect 13412 36048 13418 36100
rect 15933 36091 15991 36097
rect 15933 36057 15945 36091
rect 15979 36088 15991 36091
rect 17052 36088 17080 36116
rect 15979 36060 17080 36088
rect 18248 36088 18276 36116
rect 19720 36088 19748 36119
rect 19978 36116 19984 36128
rect 20036 36116 20042 36168
rect 20806 36156 20812 36168
rect 20719 36128 20812 36156
rect 20806 36116 20812 36128
rect 20864 36156 20870 36168
rect 22554 36156 22560 36168
rect 20864 36128 22560 36156
rect 20864 36116 20870 36128
rect 22554 36116 22560 36128
rect 22612 36116 22618 36168
rect 22646 36116 22652 36168
rect 22704 36156 22710 36168
rect 22704 36128 22749 36156
rect 22704 36116 22710 36128
rect 23474 36116 23480 36168
rect 23532 36156 23538 36168
rect 23768 36165 23796 36196
rect 24946 36184 24952 36236
rect 25004 36224 25010 36236
rect 25774 36224 25780 36236
rect 25004 36196 25780 36224
rect 25004 36184 25010 36196
rect 25774 36184 25780 36196
rect 25832 36184 25838 36236
rect 26786 36184 26792 36236
rect 26844 36224 26850 36236
rect 27724 36224 27752 36332
rect 28902 36320 28908 36332
rect 28960 36320 28966 36372
rect 29546 36224 29552 36236
rect 26844 36196 27752 36224
rect 29507 36196 29552 36224
rect 26844 36184 26850 36196
rect 29546 36184 29552 36196
rect 29604 36184 29610 36236
rect 23569 36159 23627 36165
rect 23569 36156 23581 36159
rect 23532 36128 23581 36156
rect 23532 36116 23538 36128
rect 23569 36125 23581 36128
rect 23615 36125 23627 36159
rect 23569 36119 23627 36125
rect 23753 36159 23811 36165
rect 23753 36125 23765 36159
rect 23799 36125 23811 36159
rect 23753 36119 23811 36125
rect 24581 36159 24639 36165
rect 24581 36125 24593 36159
rect 24627 36125 24639 36159
rect 24854 36156 24860 36168
rect 24815 36128 24860 36156
rect 24581 36119 24639 36125
rect 18248 36060 19748 36088
rect 21076 36091 21134 36097
rect 15979 36057 15991 36060
rect 15933 36051 15991 36057
rect 21076 36057 21088 36091
rect 21122 36088 21134 36091
rect 21910 36088 21916 36100
rect 21122 36060 21916 36088
rect 21122 36057 21134 36060
rect 21076 36051 21134 36057
rect 21910 36048 21916 36060
rect 21968 36048 21974 36100
rect 22278 36048 22284 36100
rect 22336 36088 22342 36100
rect 22925 36091 22983 36097
rect 22925 36088 22937 36091
rect 22336 36060 22937 36088
rect 22336 36048 22342 36060
rect 22925 36057 22937 36060
rect 22971 36057 22983 36091
rect 22925 36051 22983 36057
rect 23198 36048 23204 36100
rect 23256 36088 23262 36100
rect 24397 36091 24455 36097
rect 24397 36088 24409 36091
rect 23256 36060 24409 36088
rect 23256 36048 23262 36060
rect 24397 36057 24409 36060
rect 24443 36057 24455 36091
rect 24596 36088 24624 36119
rect 24854 36116 24860 36128
rect 24912 36116 24918 36168
rect 25041 36159 25099 36165
rect 25041 36125 25053 36159
rect 25087 36156 25099 36159
rect 25087 36128 25268 36156
rect 25087 36125 25099 36128
rect 25041 36119 25099 36125
rect 25130 36088 25136 36100
rect 24596 36060 25136 36088
rect 24397 36051 24455 36057
rect 25130 36048 25136 36060
rect 25188 36048 25194 36100
rect 12066 36020 12072 36032
rect 10980 35992 12072 36020
rect 12066 35980 12072 35992
rect 12124 35980 12130 36032
rect 15565 36023 15623 36029
rect 15565 35989 15577 36023
rect 15611 36020 15623 36023
rect 15838 36020 15844 36032
rect 15611 35992 15844 36020
rect 15611 35989 15623 35992
rect 15565 35983 15623 35989
rect 15838 35980 15844 35992
rect 15896 35980 15902 36032
rect 16022 35980 16028 36032
rect 16080 36020 16086 36032
rect 19150 36020 19156 36032
rect 16080 35992 19156 36020
rect 16080 35980 16086 35992
rect 19150 35980 19156 35992
rect 19208 35980 19214 36032
rect 19245 36023 19303 36029
rect 19245 35989 19257 36023
rect 19291 36020 19303 36023
rect 19518 36020 19524 36032
rect 19291 35992 19524 36020
rect 19291 35989 19303 35992
rect 19245 35983 19303 35989
rect 19518 35980 19524 35992
rect 19576 35980 19582 36032
rect 21542 35980 21548 36032
rect 21600 36020 21606 36032
rect 22189 36023 22247 36029
rect 22189 36020 22201 36023
rect 21600 35992 22201 36020
rect 21600 35980 21606 35992
rect 22189 35989 22201 35992
rect 22235 35989 22247 36023
rect 22189 35983 22247 35989
rect 23842 35980 23848 36032
rect 23900 36020 23906 36032
rect 25240 36020 25268 36128
rect 27154 36116 27160 36168
rect 27212 36156 27218 36168
rect 27801 36159 27859 36165
rect 27801 36156 27813 36159
rect 27212 36128 27813 36156
rect 27212 36116 27218 36128
rect 27801 36125 27813 36128
rect 27847 36125 27859 36159
rect 27801 36119 27859 36125
rect 28077 36159 28135 36165
rect 28077 36125 28089 36159
rect 28123 36125 28135 36159
rect 28261 36159 28319 36165
rect 28261 36156 28273 36159
rect 28077 36119 28135 36125
rect 28184 36128 28273 36156
rect 26050 36097 26056 36100
rect 26044 36051 26056 36097
rect 26108 36088 26114 36100
rect 26108 36060 26144 36088
rect 26050 36048 26056 36051
rect 26108 36048 26114 36060
rect 27430 36048 27436 36100
rect 27488 36088 27494 36100
rect 28092 36088 28120 36119
rect 27488 36060 28120 36088
rect 27488 36048 27494 36060
rect 23900 35992 25268 36020
rect 23900 35980 23906 35992
rect 26510 35980 26516 36032
rect 26568 36020 26574 36032
rect 28184 36020 28212 36128
rect 28261 36125 28273 36128
rect 28307 36156 28319 36159
rect 28534 36156 28540 36168
rect 28307 36128 28540 36156
rect 28307 36125 28319 36128
rect 28261 36119 28319 36125
rect 28534 36116 28540 36128
rect 28592 36116 28598 36168
rect 28626 36116 28632 36168
rect 28684 36156 28690 36168
rect 29805 36159 29863 36165
rect 29805 36156 29817 36159
rect 28684 36128 29817 36156
rect 28684 36116 28690 36128
rect 29805 36125 29817 36128
rect 29851 36125 29863 36159
rect 29805 36119 29863 36125
rect 28813 36091 28871 36097
rect 28813 36057 28825 36091
rect 28859 36057 28871 36091
rect 28813 36051 28871 36057
rect 26568 35992 28212 36020
rect 26568 35980 26574 35992
rect 28258 35980 28264 36032
rect 28316 36020 28322 36032
rect 28828 36020 28856 36051
rect 28316 35992 28856 36020
rect 28316 35980 28322 35992
rect 30834 35980 30840 36032
rect 30892 36020 30898 36032
rect 30929 36023 30987 36029
rect 30929 36020 30941 36023
rect 30892 35992 30941 36020
rect 30892 35980 30898 35992
rect 30929 35989 30941 35992
rect 30975 35989 30987 36023
rect 30929 35983 30987 35989
rect 1104 35930 32016 35952
rect 1104 35878 7288 35930
rect 7340 35878 17592 35930
rect 17644 35878 27896 35930
rect 27948 35878 32016 35930
rect 1104 35856 32016 35878
rect 2777 35819 2835 35825
rect 2777 35785 2789 35819
rect 2823 35816 2835 35819
rect 3234 35816 3240 35828
rect 2823 35788 3240 35816
rect 2823 35785 2835 35788
rect 2777 35779 2835 35785
rect 3234 35776 3240 35788
rect 3292 35776 3298 35828
rect 10594 35816 10600 35828
rect 3436 35788 10600 35816
rect 768 35720 1072 35748
rect 768 35476 796 35720
rect 2222 35708 2228 35760
rect 2280 35748 2286 35760
rect 3326 35748 3332 35760
rect 2280 35720 3332 35748
rect 2280 35708 2286 35720
rect 3326 35708 3332 35720
rect 3384 35708 3390 35760
rect 3436 35757 3464 35788
rect 10594 35776 10600 35788
rect 10652 35776 10658 35828
rect 11514 35776 11520 35828
rect 11572 35816 11578 35828
rect 14921 35819 14979 35825
rect 11572 35788 14872 35816
rect 11572 35776 11578 35788
rect 3421 35751 3479 35757
rect 3421 35717 3433 35751
rect 3467 35717 3479 35751
rect 3421 35711 3479 35717
rect 6365 35751 6423 35757
rect 6365 35717 6377 35751
rect 6411 35748 6423 35751
rect 6454 35748 6460 35760
rect 6411 35720 6460 35748
rect 6411 35717 6423 35720
rect 6365 35711 6423 35717
rect 6454 35708 6460 35720
rect 6512 35708 6518 35760
rect 9858 35748 9864 35760
rect 7668 35720 9864 35748
rect 1394 35680 1400 35692
rect 1355 35652 1400 35680
rect 1394 35640 1400 35652
rect 1452 35640 1458 35692
rect 1670 35689 1676 35692
rect 1664 35643 1676 35689
rect 1728 35680 1734 35692
rect 6549 35683 6607 35689
rect 1728 35652 1764 35680
rect 1670 35640 1676 35643
rect 1728 35640 1734 35652
rect 6549 35649 6561 35683
rect 6595 35649 6607 35683
rect 6549 35643 6607 35649
rect 6825 35683 6883 35689
rect 6825 35649 6837 35683
rect 6871 35649 6883 35683
rect 7006 35680 7012 35692
rect 6967 35652 7012 35680
rect 6825 35643 6883 35649
rect 6564 35544 6592 35643
rect 6840 35612 6868 35643
rect 7006 35640 7012 35652
rect 7064 35640 7070 35692
rect 7668 35689 7696 35720
rect 9858 35708 9864 35720
rect 9916 35708 9922 35760
rect 9950 35708 9956 35760
rect 10008 35748 10014 35760
rect 13354 35748 13360 35760
rect 10008 35720 12434 35748
rect 13315 35720 13360 35748
rect 10008 35708 10014 35720
rect 7653 35683 7711 35689
rect 7653 35649 7665 35683
rect 7699 35649 7711 35683
rect 7653 35643 7711 35649
rect 7920 35683 7978 35689
rect 7920 35649 7932 35683
rect 7966 35680 7978 35683
rect 8938 35680 8944 35692
rect 7966 35652 8944 35680
rect 7966 35649 7978 35652
rect 7920 35643 7978 35649
rect 8938 35640 8944 35652
rect 8996 35640 9002 35692
rect 9674 35640 9680 35692
rect 9732 35680 9738 35692
rect 10781 35683 10839 35689
rect 10781 35680 10793 35683
rect 9732 35652 10793 35680
rect 9732 35640 9738 35652
rect 10781 35649 10793 35652
rect 10827 35680 10839 35683
rect 10870 35680 10876 35692
rect 10827 35652 10876 35680
rect 10827 35649 10839 35652
rect 10781 35643 10839 35649
rect 10870 35640 10876 35652
rect 10928 35640 10934 35692
rect 10965 35683 11023 35689
rect 10965 35649 10977 35683
rect 11011 35680 11023 35683
rect 11054 35680 11060 35692
rect 11011 35652 11060 35680
rect 11011 35649 11023 35652
rect 10965 35643 11023 35649
rect 11054 35640 11060 35652
rect 11112 35640 11118 35692
rect 11606 35640 11612 35692
rect 11664 35680 11670 35692
rect 11773 35683 11831 35689
rect 11773 35680 11785 35683
rect 11664 35652 11785 35680
rect 11664 35640 11670 35652
rect 11773 35649 11785 35652
rect 11819 35649 11831 35683
rect 12406 35680 12434 35720
rect 13354 35708 13360 35720
rect 13412 35708 13418 35760
rect 13446 35708 13452 35760
rect 13504 35748 13510 35760
rect 14553 35751 14611 35757
rect 14553 35748 14565 35751
rect 13504 35720 14565 35748
rect 13504 35708 13510 35720
rect 14553 35717 14565 35720
rect 14599 35717 14611 35751
rect 14553 35711 14611 35717
rect 14642 35708 14648 35760
rect 14700 35748 14706 35760
rect 14753 35751 14811 35757
rect 14753 35748 14765 35751
rect 14700 35720 14765 35748
rect 14700 35708 14706 35720
rect 14753 35717 14765 35720
rect 14799 35717 14811 35751
rect 14753 35711 14811 35717
rect 13538 35680 13544 35692
rect 12406 35652 13400 35680
rect 13499 35652 13544 35680
rect 11773 35643 11831 35649
rect 6914 35612 6920 35624
rect 6840 35584 6920 35612
rect 6914 35572 6920 35584
rect 6972 35572 6978 35624
rect 9030 35572 9036 35624
rect 9088 35612 9094 35624
rect 9493 35615 9551 35621
rect 9493 35612 9505 35615
rect 9088 35584 9505 35612
rect 9088 35572 9094 35584
rect 9493 35581 9505 35584
rect 9539 35581 9551 35615
rect 9493 35575 9551 35581
rect 9582 35572 9588 35624
rect 9640 35612 9646 35624
rect 9769 35615 9827 35621
rect 9769 35612 9781 35615
rect 9640 35584 9781 35612
rect 9640 35572 9646 35584
rect 9769 35581 9781 35584
rect 9815 35581 9827 35615
rect 11514 35612 11520 35624
rect 11475 35584 11520 35612
rect 9769 35575 9827 35581
rect 11514 35572 11520 35584
rect 11572 35572 11578 35624
rect 7006 35544 7012 35556
rect 6564 35516 7012 35544
rect 7006 35504 7012 35516
rect 7064 35504 7070 35556
rect 10042 35504 10048 35556
rect 10100 35544 10106 35556
rect 10873 35547 10931 35553
rect 10873 35544 10885 35547
rect 10100 35516 10885 35544
rect 10100 35504 10106 35516
rect 10873 35513 10885 35516
rect 10919 35513 10931 35547
rect 13372 35544 13400 35652
rect 13538 35640 13544 35652
rect 13596 35640 13602 35692
rect 13722 35680 13728 35692
rect 13683 35652 13728 35680
rect 13722 35640 13728 35652
rect 13780 35640 13786 35692
rect 14844 35680 14872 35788
rect 14921 35785 14933 35819
rect 14967 35785 14979 35819
rect 20806 35816 20812 35828
rect 14921 35779 14979 35785
rect 15488 35788 20812 35816
rect 14936 35748 14964 35779
rect 15102 35748 15108 35760
rect 14936 35720 15108 35748
rect 15102 35708 15108 35720
rect 15160 35708 15166 35760
rect 15488 35680 15516 35788
rect 20806 35776 20812 35788
rect 20864 35776 20870 35828
rect 22066 35788 32352 35816
rect 15838 35748 15844 35760
rect 15799 35720 15844 35748
rect 15838 35708 15844 35720
rect 15896 35708 15902 35760
rect 22066 35748 22094 35788
rect 24946 35748 24952 35760
rect 16868 35720 18736 35748
rect 16868 35692 16896 35720
rect 14844 35652 15516 35680
rect 15562 35640 15568 35692
rect 15620 35680 15626 35692
rect 15749 35683 15807 35689
rect 15749 35680 15761 35683
rect 15620 35652 15761 35680
rect 15620 35640 15626 35652
rect 15749 35649 15761 35652
rect 15795 35649 15807 35683
rect 16850 35680 16856 35692
rect 16811 35652 16856 35680
rect 15749 35643 15807 35649
rect 16850 35640 16856 35652
rect 16908 35640 16914 35692
rect 17120 35683 17178 35689
rect 17120 35649 17132 35683
rect 17166 35680 17178 35683
rect 17402 35680 17408 35692
rect 17166 35652 17408 35680
rect 17166 35649 17178 35652
rect 17120 35643 17178 35649
rect 17402 35640 17408 35652
rect 17460 35640 17466 35692
rect 18708 35689 18736 35720
rect 18800 35720 22094 35748
rect 24412 35720 24952 35748
rect 18693 35683 18751 35689
rect 18693 35649 18705 35683
rect 18739 35649 18751 35683
rect 18693 35643 18751 35649
rect 13817 35615 13875 35621
rect 13817 35581 13829 35615
rect 13863 35612 13875 35615
rect 15654 35612 15660 35624
rect 13863 35584 15660 35612
rect 13863 35581 13875 35584
rect 13817 35575 13875 35581
rect 15654 35572 15660 35584
rect 15712 35572 15718 35624
rect 15930 35612 15936 35624
rect 15891 35584 15936 35612
rect 15930 35572 15936 35584
rect 15988 35572 15994 35624
rect 18800 35612 18828 35720
rect 18960 35683 19018 35689
rect 18960 35649 18972 35683
rect 19006 35680 19018 35683
rect 19242 35680 19248 35692
rect 19006 35652 19248 35680
rect 19006 35649 19018 35652
rect 18960 35643 19018 35649
rect 19242 35640 19248 35652
rect 19300 35640 19306 35692
rect 20898 35680 20904 35692
rect 20859 35652 20904 35680
rect 20898 35640 20904 35652
rect 20956 35640 20962 35692
rect 20993 35683 21051 35689
rect 20993 35649 21005 35683
rect 21039 35649 21051 35683
rect 20993 35643 21051 35649
rect 21085 35683 21143 35689
rect 21085 35649 21097 35683
rect 21131 35680 21143 35683
rect 21542 35680 21548 35692
rect 21131 35652 21548 35680
rect 21131 35649 21143 35652
rect 21085 35643 21143 35649
rect 17880 35584 18828 35612
rect 21008 35612 21036 35643
rect 21542 35640 21548 35652
rect 21600 35640 21606 35692
rect 21726 35640 21732 35692
rect 21784 35680 21790 35692
rect 21821 35683 21879 35689
rect 21821 35680 21833 35683
rect 21784 35652 21833 35680
rect 21784 35640 21790 35652
rect 21821 35649 21833 35652
rect 21867 35649 21879 35683
rect 21821 35643 21879 35649
rect 22732 35683 22790 35689
rect 22732 35649 22744 35683
rect 22778 35680 22790 35683
rect 23014 35680 23020 35692
rect 22778 35652 23020 35680
rect 22778 35649 22790 35652
rect 22732 35643 22790 35649
rect 23014 35640 23020 35652
rect 23072 35640 23078 35692
rect 24412 35689 24440 35720
rect 24946 35708 24952 35720
rect 25004 35708 25010 35760
rect 25038 35708 25044 35760
rect 25096 35748 25102 35760
rect 25096 35720 27292 35748
rect 25096 35708 25102 35720
rect 24670 35689 24676 35692
rect 24397 35683 24455 35689
rect 24397 35649 24409 35683
rect 24443 35649 24455 35683
rect 24664 35680 24676 35689
rect 24631 35652 24676 35680
rect 24397 35643 24455 35649
rect 24664 35643 24676 35652
rect 24670 35640 24676 35643
rect 24728 35640 24734 35692
rect 26421 35683 26479 35689
rect 26421 35649 26433 35683
rect 26467 35680 26479 35683
rect 26602 35680 26608 35692
rect 26467 35652 26608 35680
rect 26467 35649 26479 35652
rect 26421 35643 26479 35649
rect 26602 35640 26608 35652
rect 26660 35640 26666 35692
rect 27154 35680 27160 35692
rect 27115 35652 27160 35680
rect 27154 35640 27160 35652
rect 27212 35640 27218 35692
rect 21174 35612 21180 35624
rect 21008 35584 21180 35612
rect 13372 35516 15516 35544
rect 10873 35507 10931 35513
rect 768 35448 888 35476
rect 0 35340 800 35354
rect 860 35340 888 35448
rect 3786 35436 3792 35488
rect 3844 35476 3850 35488
rect 4709 35479 4767 35485
rect 4709 35476 4721 35479
rect 3844 35448 4721 35476
rect 3844 35436 3850 35448
rect 4709 35445 4721 35448
rect 4755 35445 4767 35479
rect 4709 35439 4767 35445
rect 9033 35479 9091 35485
rect 9033 35445 9045 35479
rect 9079 35476 9091 35479
rect 9214 35476 9220 35488
rect 9079 35448 9220 35476
rect 9079 35445 9091 35448
rect 9033 35439 9091 35445
rect 9214 35436 9220 35448
rect 9272 35436 9278 35488
rect 12894 35476 12900 35488
rect 12855 35448 12900 35476
rect 12894 35436 12900 35448
rect 12952 35436 12958 35488
rect 14737 35479 14795 35485
rect 14737 35445 14749 35479
rect 14783 35476 14795 35479
rect 15194 35476 15200 35488
rect 14783 35448 15200 35476
rect 14783 35445 14795 35448
rect 14737 35439 14795 35445
rect 15194 35436 15200 35448
rect 15252 35436 15258 35488
rect 15286 35436 15292 35488
rect 15344 35476 15350 35488
rect 15381 35479 15439 35485
rect 15381 35476 15393 35479
rect 15344 35448 15393 35476
rect 15344 35436 15350 35448
rect 15381 35445 15393 35448
rect 15427 35445 15439 35479
rect 15488 35476 15516 35516
rect 17880 35476 17908 35584
rect 21174 35572 21180 35584
rect 21232 35572 21238 35624
rect 21634 35572 21640 35624
rect 21692 35612 21698 35624
rect 22465 35615 22523 35621
rect 22465 35612 22477 35615
rect 21692 35584 22477 35612
rect 21692 35572 21698 35584
rect 22465 35581 22477 35584
rect 22511 35581 22523 35615
rect 22465 35575 22523 35581
rect 21542 35504 21548 35556
rect 21600 35544 21606 35556
rect 21913 35547 21971 35553
rect 21913 35544 21925 35547
rect 21600 35516 21925 35544
rect 21600 35504 21606 35516
rect 21913 35513 21925 35516
rect 21959 35513 21971 35547
rect 23842 35544 23848 35556
rect 23803 35516 23848 35544
rect 21913 35507 21971 35513
rect 23842 35504 23848 35516
rect 23900 35504 23906 35556
rect 26237 35547 26295 35553
rect 26237 35544 26249 35547
rect 25332 35516 26249 35544
rect 18230 35476 18236 35488
rect 15488 35448 17908 35476
rect 18191 35448 18236 35476
rect 15381 35439 15439 35445
rect 18230 35436 18236 35448
rect 18288 35436 18294 35488
rect 18690 35436 18696 35488
rect 18748 35476 18754 35488
rect 19978 35476 19984 35488
rect 18748 35448 19984 35476
rect 18748 35436 18754 35448
rect 19978 35436 19984 35448
rect 20036 35476 20042 35488
rect 20073 35479 20131 35485
rect 20073 35476 20085 35479
rect 20036 35448 20085 35476
rect 20036 35436 20042 35448
rect 20073 35445 20085 35448
rect 20119 35445 20131 35479
rect 20073 35439 20131 35445
rect 21269 35479 21327 35485
rect 21269 35445 21281 35479
rect 21315 35476 21327 35479
rect 21634 35476 21640 35488
rect 21315 35448 21640 35476
rect 21315 35445 21327 35448
rect 21269 35439 21327 35445
rect 21634 35436 21640 35448
rect 21692 35436 21698 35488
rect 22370 35436 22376 35488
rect 22428 35476 22434 35488
rect 25038 35476 25044 35488
rect 22428 35448 25044 35476
rect 22428 35436 22434 35448
rect 25038 35436 25044 35448
rect 25096 35436 25102 35488
rect 25130 35436 25136 35488
rect 25188 35476 25194 35488
rect 25332 35476 25360 35516
rect 26237 35513 26249 35516
rect 26283 35544 26295 35547
rect 27172 35544 27200 35640
rect 27264 35612 27292 35720
rect 27338 35708 27344 35760
rect 27396 35748 27402 35760
rect 27396 35720 27660 35748
rect 27396 35708 27402 35720
rect 27430 35680 27436 35692
rect 27391 35652 27436 35680
rect 27430 35640 27436 35652
rect 27488 35640 27494 35692
rect 27632 35689 27660 35720
rect 28534 35708 28540 35760
rect 28592 35748 28598 35760
rect 30162 35751 30220 35757
rect 30162 35748 30174 35751
rect 28592 35720 30174 35748
rect 28592 35708 28598 35720
rect 30162 35717 30174 35720
rect 30208 35717 30220 35751
rect 30162 35711 30220 35717
rect 27617 35683 27675 35689
rect 27617 35649 27629 35683
rect 27663 35649 27675 35683
rect 28166 35680 28172 35692
rect 28127 35652 28172 35680
rect 27617 35643 27675 35649
rect 28166 35640 28172 35652
rect 28224 35640 28230 35692
rect 28997 35683 29055 35689
rect 28997 35649 29009 35683
rect 29043 35649 29055 35683
rect 29270 35680 29276 35692
rect 29231 35652 29276 35680
rect 28997 35643 29055 35649
rect 28442 35612 28448 35624
rect 27264 35584 28448 35612
rect 28442 35572 28448 35584
rect 28500 35572 28506 35624
rect 29012 35612 29040 35643
rect 29270 35640 29276 35652
rect 29328 35640 29334 35692
rect 29454 35680 29460 35692
rect 29415 35652 29460 35680
rect 29454 35640 29460 35652
rect 29512 35640 29518 35692
rect 29730 35612 29736 35624
rect 29012 35584 29736 35612
rect 29730 35572 29736 35584
rect 29788 35572 29794 35624
rect 29917 35615 29975 35621
rect 29917 35581 29929 35615
rect 29963 35581 29975 35615
rect 29917 35575 29975 35581
rect 26283 35516 27200 35544
rect 26283 35513 26295 35516
rect 26237 35507 26295 35513
rect 27246 35504 27252 35556
rect 27304 35544 27310 35556
rect 27304 35516 28856 35544
rect 27304 35504 27310 35516
rect 25774 35476 25780 35488
rect 25188 35448 25360 35476
rect 25735 35448 25780 35476
rect 25188 35436 25194 35448
rect 25774 35436 25780 35448
rect 25832 35436 25838 35488
rect 26326 35436 26332 35488
rect 26384 35476 26390 35488
rect 26973 35479 27031 35485
rect 26973 35476 26985 35479
rect 26384 35448 26985 35476
rect 26384 35436 26390 35448
rect 26973 35445 26985 35448
rect 27019 35445 27031 35479
rect 26973 35439 27031 35445
rect 28074 35436 28080 35488
rect 28132 35476 28138 35488
rect 28258 35476 28264 35488
rect 28132 35448 28264 35476
rect 28132 35436 28138 35448
rect 28258 35436 28264 35448
rect 28316 35436 28322 35488
rect 28828 35485 28856 35516
rect 28994 35504 29000 35556
rect 29052 35544 29058 35556
rect 29546 35544 29552 35556
rect 29052 35516 29552 35544
rect 29052 35504 29058 35516
rect 29546 35504 29552 35516
rect 29604 35544 29610 35556
rect 29932 35544 29960 35575
rect 29604 35516 29960 35544
rect 29604 35504 29610 35516
rect 28813 35479 28871 35485
rect 28813 35445 28825 35479
rect 28859 35445 28871 35479
rect 31294 35476 31300 35488
rect 31255 35448 31300 35476
rect 28813 35439 28871 35445
rect 31294 35436 31300 35448
rect 31352 35436 31358 35488
rect 32324 35476 32352 35788
rect 32232 35448 32352 35476
rect 0 35312 888 35340
rect 1104 35386 32016 35408
rect 1104 35334 2136 35386
rect 2188 35334 12440 35386
rect 12492 35334 22744 35386
rect 22796 35334 32016 35386
rect 1104 35312 32016 35334
rect 32232 35340 32260 35448
rect 32320 35340 33120 35354
rect 32232 35312 33120 35340
rect 0 35298 800 35312
rect 32320 35298 33120 35312
rect 1670 35232 1676 35284
rect 1728 35272 1734 35284
rect 1857 35275 1915 35281
rect 1857 35272 1869 35275
rect 1728 35244 1869 35272
rect 1728 35232 1734 35244
rect 1857 35241 1869 35244
rect 1903 35241 1915 35275
rect 2222 35272 2228 35284
rect 2183 35244 2228 35272
rect 1857 35235 1915 35241
rect 2222 35232 2228 35244
rect 2280 35272 2286 35284
rect 3145 35275 3203 35281
rect 3145 35272 3157 35275
rect 2280 35244 3157 35272
rect 2280 35232 2286 35244
rect 3145 35241 3157 35244
rect 3191 35241 3203 35275
rect 5074 35272 5080 35284
rect 3145 35235 3203 35241
rect 3804 35244 5080 35272
rect 3804 35204 3832 35244
rect 5074 35232 5080 35244
rect 5132 35232 5138 35284
rect 6457 35275 6515 35281
rect 6457 35241 6469 35275
rect 6503 35272 6515 35275
rect 6546 35272 6552 35284
rect 6503 35244 6552 35272
rect 6503 35241 6515 35244
rect 6457 35235 6515 35241
rect 6546 35232 6552 35244
rect 6604 35232 6610 35284
rect 8938 35272 8944 35284
rect 8899 35244 8944 35272
rect 8938 35232 8944 35244
rect 8996 35232 9002 35284
rect 12069 35275 12127 35281
rect 12069 35241 12081 35275
rect 12115 35272 12127 35275
rect 12894 35272 12900 35284
rect 12115 35244 12900 35272
rect 12115 35241 12127 35244
rect 12069 35235 12127 35241
rect 12894 35232 12900 35244
rect 12952 35232 12958 35284
rect 14918 35272 14924 35284
rect 14879 35244 14924 35272
rect 14918 35232 14924 35244
rect 14976 35232 14982 35284
rect 15562 35272 15568 35284
rect 15523 35244 15568 35272
rect 15562 35232 15568 35244
rect 15620 35232 15626 35284
rect 16942 35232 16948 35284
rect 17000 35272 17006 35284
rect 17129 35275 17187 35281
rect 17129 35272 17141 35275
rect 17000 35244 17141 35272
rect 17000 35232 17006 35244
rect 17129 35241 17141 35244
rect 17175 35241 17187 35275
rect 17129 35235 17187 35241
rect 17589 35275 17647 35281
rect 17589 35241 17601 35275
rect 17635 35272 17647 35275
rect 17862 35272 17868 35284
rect 17635 35244 17868 35272
rect 17635 35241 17647 35244
rect 17589 35235 17647 35241
rect 17862 35232 17868 35244
rect 17920 35232 17926 35284
rect 18049 35275 18107 35281
rect 18049 35241 18061 35275
rect 18095 35272 18107 35275
rect 19242 35272 19248 35284
rect 18095 35244 18828 35272
rect 19203 35244 19248 35272
rect 18095 35241 18107 35244
rect 18049 35235 18107 35241
rect 5169 35207 5227 35213
rect 5169 35204 5181 35207
rect 2332 35176 3832 35204
rect 4816 35176 5181 35204
rect 2332 35145 2360 35176
rect 2317 35139 2375 35145
rect 2317 35105 2329 35139
rect 2363 35105 2375 35139
rect 2317 35099 2375 35105
rect 2682 35096 2688 35148
rect 2740 35136 2746 35148
rect 3786 35136 3792 35148
rect 2740 35108 3792 35136
rect 2740 35096 2746 35108
rect 3786 35096 3792 35108
rect 3844 35096 3850 35148
rect 2038 35068 2044 35080
rect 1999 35040 2044 35068
rect 2038 35028 2044 35040
rect 2096 35028 2102 35080
rect 2958 35068 2964 35080
rect 2919 35040 2964 35068
rect 2958 35028 2964 35040
rect 3016 35028 3022 35080
rect 3237 35071 3295 35077
rect 3237 35037 3249 35071
rect 3283 35068 3295 35071
rect 4338 35068 4344 35080
rect 3283 35040 4344 35068
rect 3283 35037 3295 35040
rect 3237 35031 3295 35037
rect 4338 35028 4344 35040
rect 4396 35068 4402 35080
rect 4816 35068 4844 35176
rect 5169 35173 5181 35176
rect 5215 35173 5227 35207
rect 5169 35167 5227 35173
rect 8110 35164 8116 35216
rect 8168 35204 8174 35216
rect 9309 35207 9367 35213
rect 9309 35204 9321 35207
rect 8168 35176 9321 35204
rect 8168 35164 8174 35176
rect 9309 35173 9321 35176
rect 9355 35173 9367 35207
rect 9309 35167 9367 35173
rect 10962 35164 10968 35216
rect 11020 35204 11026 35216
rect 11701 35207 11759 35213
rect 11701 35204 11713 35207
rect 11020 35176 11713 35204
rect 11020 35164 11026 35176
rect 11701 35173 11713 35176
rect 11747 35173 11759 35207
rect 13538 35204 13544 35216
rect 13451 35176 13544 35204
rect 11701 35167 11759 35173
rect 13538 35164 13544 35176
rect 13596 35204 13602 35216
rect 16022 35204 16028 35216
rect 13596 35176 16028 35204
rect 13596 35164 13602 35176
rect 16022 35164 16028 35176
rect 16080 35164 16086 35216
rect 17405 35207 17463 35213
rect 17405 35173 17417 35207
rect 17451 35204 17463 35207
rect 18690 35204 18696 35216
rect 17451 35176 18696 35204
rect 17451 35173 17463 35176
rect 17405 35167 17463 35173
rect 18690 35164 18696 35176
rect 18748 35164 18754 35216
rect 18800 35204 18828 35244
rect 19242 35232 19248 35244
rect 19300 35232 19306 35284
rect 19334 35232 19340 35284
rect 19392 35272 19398 35284
rect 19392 35244 21956 35272
rect 19392 35232 19398 35244
rect 19426 35204 19432 35216
rect 18800 35176 19432 35204
rect 19426 35164 19432 35176
rect 19484 35164 19490 35216
rect 19613 35207 19671 35213
rect 19613 35173 19625 35207
rect 19659 35204 19671 35207
rect 20806 35204 20812 35216
rect 19659 35176 20812 35204
rect 19659 35173 19671 35176
rect 19613 35167 19671 35173
rect 20806 35164 20812 35176
rect 20864 35164 20870 35216
rect 21450 35164 21456 35216
rect 21508 35204 21514 35216
rect 21928 35204 21956 35244
rect 22002 35232 22008 35284
rect 22060 35272 22066 35284
rect 22094 35272 22100 35284
rect 22060 35244 22100 35272
rect 22060 35232 22066 35244
rect 22094 35232 22100 35244
rect 22152 35232 22158 35284
rect 23014 35272 23020 35284
rect 22975 35244 23020 35272
rect 23014 35232 23020 35244
rect 23072 35232 23078 35284
rect 24949 35275 25007 35281
rect 24949 35241 24961 35275
rect 24995 35272 25007 35275
rect 25222 35272 25228 35284
rect 24995 35244 25228 35272
rect 24995 35241 25007 35244
rect 24949 35235 25007 35241
rect 25222 35232 25228 35244
rect 25280 35232 25286 35284
rect 26050 35272 26056 35284
rect 26011 35244 26056 35272
rect 26050 35232 26056 35244
rect 26108 35232 26114 35284
rect 26142 35232 26148 35284
rect 26200 35272 26206 35284
rect 26421 35275 26479 35281
rect 26421 35272 26433 35275
rect 26200 35244 26433 35272
rect 26200 35232 26206 35244
rect 26421 35241 26433 35244
rect 26467 35272 26479 35275
rect 28997 35275 29055 35281
rect 26467 35244 28580 35272
rect 26467 35241 26479 35244
rect 26421 35235 26479 35241
rect 22646 35204 22652 35216
rect 21508 35176 21864 35204
rect 21928 35176 22652 35204
rect 21508 35164 21514 35176
rect 7006 35136 7012 35148
rect 6656 35108 7012 35136
rect 6656 35077 6684 35108
rect 7006 35096 7012 35108
rect 7064 35136 7070 35148
rect 9401 35139 9459 35145
rect 9401 35136 9413 35139
rect 7064 35108 7788 35136
rect 7064 35096 7070 35108
rect 4396 35040 4844 35068
rect 6641 35071 6699 35077
rect 4396 35028 4402 35040
rect 6641 35037 6653 35071
rect 6687 35037 6699 35071
rect 6914 35068 6920 35080
rect 6875 35040 6920 35068
rect 6641 35031 6699 35037
rect 6914 35028 6920 35040
rect 6972 35028 6978 35080
rect 7098 35068 7104 35080
rect 7059 35040 7104 35068
rect 7098 35028 7104 35040
rect 7156 35028 7162 35080
rect 7760 35077 7788 35108
rect 8312 35108 9413 35136
rect 8312 35080 8340 35108
rect 9401 35105 9413 35108
rect 9447 35105 9459 35139
rect 11882 35136 11888 35148
rect 9401 35099 9459 35105
rect 10888 35108 11888 35136
rect 7745 35071 7803 35077
rect 7745 35037 7757 35071
rect 7791 35068 7803 35071
rect 7926 35068 7932 35080
rect 7791 35040 7932 35068
rect 7791 35037 7803 35040
rect 7745 35031 7803 35037
rect 7926 35028 7932 35040
rect 7984 35028 7990 35080
rect 8021 35071 8079 35077
rect 8021 35037 8033 35071
rect 8067 35037 8079 35071
rect 8021 35031 8079 35037
rect 8205 35071 8263 35077
rect 8205 35037 8217 35071
rect 8251 35068 8263 35071
rect 8294 35068 8300 35080
rect 8251 35040 8300 35068
rect 8251 35037 8263 35040
rect 8205 35031 8263 35037
rect 1946 34960 1952 35012
rect 2004 35000 2010 35012
rect 4034 35003 4092 35009
rect 4034 35000 4046 35003
rect 2004 34972 4046 35000
rect 2004 34960 2010 34972
rect 4034 34969 4046 34972
rect 4080 34969 4092 35003
rect 6932 35000 6960 35028
rect 8036 35000 8064 35031
rect 8294 35028 8300 35040
rect 8352 35028 8358 35080
rect 9122 35068 9128 35080
rect 9083 35040 9128 35068
rect 9122 35028 9128 35040
rect 9180 35028 9186 35080
rect 9858 35068 9864 35080
rect 9771 35040 9864 35068
rect 9858 35028 9864 35040
rect 9916 35068 9922 35080
rect 10888 35068 10916 35108
rect 11882 35096 11888 35108
rect 11940 35096 11946 35148
rect 14550 35136 14556 35148
rect 14511 35108 14556 35136
rect 14550 35096 14556 35108
rect 14608 35096 14614 35148
rect 20898 35136 20904 35148
rect 14660 35108 17678 35136
rect 14660 35068 14688 35108
rect 9916 35040 10916 35068
rect 10980 35040 14688 35068
rect 14737 35071 14795 35077
rect 9916 35028 9922 35040
rect 9398 35000 9404 35012
rect 6932 34972 9404 35000
rect 4034 34963 4092 34969
rect 9398 34960 9404 34972
rect 9456 35000 9462 35012
rect 9582 35000 9588 35012
rect 9456 34972 9588 35000
rect 9456 34960 9462 34972
rect 9582 34960 9588 34972
rect 9640 34960 9646 35012
rect 10128 35003 10186 35009
rect 10128 34969 10140 35003
rect 10174 35000 10186 35003
rect 10502 35000 10508 35012
rect 10174 34972 10508 35000
rect 10174 34969 10186 34972
rect 10128 34963 10186 34969
rect 10502 34960 10508 34972
rect 10560 34960 10566 35012
rect 10778 34960 10784 35012
rect 10836 35000 10842 35012
rect 10980 35000 11008 35040
rect 14737 35037 14749 35071
rect 14783 35037 14795 35071
rect 15378 35068 15384 35080
rect 15339 35040 15384 35068
rect 14737 35031 14795 35037
rect 13354 35000 13360 35012
rect 10836 34972 11008 35000
rect 13315 34972 13360 35000
rect 10836 34960 10842 34972
rect 13354 34960 13360 34972
rect 13412 34960 13418 35012
rect 14642 34960 14648 35012
rect 14700 35000 14706 35012
rect 14752 35000 14780 35031
rect 15378 35028 15384 35040
rect 15436 35028 15442 35080
rect 16577 35071 16635 35077
rect 16577 35037 16589 35071
rect 16623 35037 16635 35071
rect 16577 35031 16635 35037
rect 16390 35000 16396 35012
rect 14700 34972 14780 35000
rect 14844 34972 16396 35000
rect 14700 34960 14706 34972
rect 2774 34932 2780 34944
rect 2735 34904 2780 34932
rect 2774 34892 2780 34904
rect 2832 34892 2838 34944
rect 6914 34892 6920 34944
rect 6972 34932 6978 34944
rect 7466 34932 7472 34944
rect 6972 34904 7472 34932
rect 6972 34892 6978 34904
rect 7466 34892 7472 34904
rect 7524 34892 7530 34944
rect 7561 34935 7619 34941
rect 7561 34901 7573 34935
rect 7607 34932 7619 34935
rect 7742 34932 7748 34944
rect 7607 34904 7748 34932
rect 7607 34901 7619 34904
rect 7561 34895 7619 34901
rect 7742 34892 7748 34904
rect 7800 34892 7806 34944
rect 11054 34892 11060 34944
rect 11112 34932 11118 34944
rect 11241 34935 11299 34941
rect 11241 34932 11253 34935
rect 11112 34904 11253 34932
rect 11112 34892 11118 34904
rect 11241 34901 11253 34904
rect 11287 34932 11299 34935
rect 12069 34935 12127 34941
rect 12069 34932 12081 34935
rect 11287 34904 12081 34932
rect 11287 34901 11299 34904
rect 11241 34895 11299 34901
rect 12069 34901 12081 34904
rect 12115 34901 12127 34935
rect 12250 34932 12256 34944
rect 12211 34904 12256 34932
rect 12069 34895 12127 34901
rect 12250 34892 12256 34904
rect 12308 34892 12314 34944
rect 13078 34892 13084 34944
rect 13136 34932 13142 34944
rect 14844 34932 14872 34972
rect 16390 34960 16396 34972
rect 16448 34960 16454 35012
rect 13136 34904 14872 34932
rect 13136 34892 13142 34904
rect 15378 34892 15384 34944
rect 15436 34932 15442 34944
rect 16482 34932 16488 34944
rect 15436 34904 16488 34932
rect 15436 34892 15442 34904
rect 16482 34892 16488 34904
rect 16540 34892 16546 34944
rect 16592 34932 16620 35031
rect 16666 35028 16672 35080
rect 16724 35068 16730 35080
rect 16761 35071 16819 35077
rect 16761 35068 16773 35071
rect 16724 35040 16773 35068
rect 16724 35028 16730 35040
rect 16761 35037 16773 35040
rect 16807 35037 16819 35071
rect 16761 35031 16819 35037
rect 16945 35071 17003 35077
rect 16945 35037 16957 35071
rect 16991 35068 17003 35071
rect 17126 35068 17132 35080
rect 16991 35040 17132 35068
rect 16991 35037 17003 35040
rect 16945 35031 17003 35037
rect 17126 35028 17132 35040
rect 17184 35028 17190 35080
rect 17650 35062 17678 35108
rect 19352 35108 20904 35136
rect 17773 35071 17831 35077
rect 17773 35062 17785 35071
rect 17650 35037 17785 35062
rect 17819 35037 17831 35071
rect 17650 35034 17831 35037
rect 17773 35031 17831 35034
rect 17954 35028 17960 35080
rect 18012 35068 18018 35080
rect 18693 35071 18751 35077
rect 18693 35068 18705 35071
rect 18012 35040 18705 35068
rect 18012 35028 18018 35040
rect 18693 35037 18705 35040
rect 18739 35068 18751 35071
rect 18874 35068 18880 35080
rect 18739 35040 18880 35068
rect 18739 35037 18751 35040
rect 18693 35031 18751 35037
rect 18874 35028 18880 35040
rect 18932 35068 18938 35080
rect 19352 35068 19380 35108
rect 20898 35096 20904 35108
rect 20956 35096 20962 35148
rect 21836 35136 21864 35176
rect 22646 35164 22652 35176
rect 22704 35164 22710 35216
rect 23106 35164 23112 35216
rect 23164 35204 23170 35216
rect 23385 35207 23443 35213
rect 23385 35204 23397 35207
rect 23164 35176 23397 35204
rect 23164 35164 23170 35176
rect 23385 35173 23397 35176
rect 23431 35204 23443 35207
rect 26160 35204 26188 35232
rect 23431 35176 26188 35204
rect 23431 35173 23443 35176
rect 23385 35167 23443 35173
rect 26234 35164 26240 35216
rect 26292 35204 26298 35216
rect 27246 35204 27252 35216
rect 26292 35176 27252 35204
rect 26292 35164 26298 35176
rect 27246 35164 27252 35176
rect 27304 35164 27310 35216
rect 28552 35204 28580 35244
rect 28997 35241 29009 35275
rect 29043 35272 29055 35275
rect 29178 35272 29184 35284
rect 29043 35244 29184 35272
rect 29043 35241 29055 35244
rect 28997 35235 29055 35241
rect 29178 35232 29184 35244
rect 29236 35272 29242 35284
rect 29454 35272 29460 35284
rect 29236 35244 29460 35272
rect 29236 35232 29242 35244
rect 29454 35232 29460 35244
rect 29512 35232 29518 35284
rect 29089 35207 29147 35213
rect 29089 35204 29101 35207
rect 28552 35176 29101 35204
rect 29089 35173 29101 35176
rect 29135 35173 29147 35207
rect 29089 35167 29147 35173
rect 29270 35164 29276 35216
rect 29328 35204 29334 35216
rect 29328 35176 30604 35204
rect 29328 35164 29334 35176
rect 21913 35139 21971 35145
rect 21913 35136 21925 35139
rect 21836 35108 21925 35136
rect 21913 35105 21925 35108
rect 21959 35105 21971 35139
rect 21913 35099 21971 35105
rect 25958 35096 25964 35148
rect 26016 35136 26022 35148
rect 26016 35108 27568 35136
rect 26016 35096 26022 35108
rect 18932 35040 19380 35068
rect 19429 35071 19487 35077
rect 18932 35028 18938 35040
rect 19429 35037 19441 35071
rect 19475 35068 19487 35071
rect 19518 35068 19524 35080
rect 19475 35040 19524 35068
rect 19475 35037 19487 35040
rect 19429 35031 19487 35037
rect 19518 35028 19524 35040
rect 19576 35028 19582 35080
rect 19705 35071 19763 35077
rect 19705 35037 19717 35071
rect 19751 35037 19763 35071
rect 20162 35068 20168 35080
rect 20123 35040 20168 35068
rect 19705 35031 19763 35037
rect 16853 35003 16911 35009
rect 16853 34969 16865 35003
rect 16899 35000 16911 35003
rect 17405 35003 17463 35009
rect 17405 35000 17417 35003
rect 16899 34972 17417 35000
rect 16899 34969 16911 34972
rect 16853 34963 16911 34969
rect 17405 34969 17417 34972
rect 17451 34969 17463 35003
rect 17405 34963 17463 34969
rect 17494 34960 17500 35012
rect 17552 35000 17558 35012
rect 18049 35003 18107 35009
rect 18049 35000 18061 35003
rect 17552 34972 18061 35000
rect 17552 34960 17558 34972
rect 18049 34969 18061 34972
rect 18095 34969 18107 35003
rect 19720 35000 19748 35031
rect 20162 35028 20168 35040
rect 20220 35028 20226 35080
rect 20809 35071 20867 35077
rect 20809 35068 20821 35071
rect 20272 35040 20821 35068
rect 18049 34963 18107 34969
rect 18248 34972 19748 35000
rect 18248 34944 18276 34972
rect 18230 34932 18236 34944
rect 16592 34904 18236 34932
rect 18230 34892 18236 34904
rect 18288 34892 18294 34944
rect 18509 34935 18567 34941
rect 18509 34901 18521 34935
rect 18555 34932 18567 34935
rect 19150 34932 19156 34944
rect 18555 34904 19156 34932
rect 18555 34901 18567 34904
rect 18509 34895 18567 34901
rect 19150 34892 19156 34904
rect 19208 34892 19214 34944
rect 20070 34892 20076 34944
rect 20128 34932 20134 34944
rect 20272 34941 20300 35040
rect 20809 35037 20821 35040
rect 20855 35037 20867 35071
rect 21174 35068 21180 35080
rect 21135 35040 21180 35068
rect 20809 35031 20867 35037
rect 20824 35000 20852 35031
rect 21174 35028 21180 35040
rect 21232 35028 21238 35080
rect 21358 35028 21364 35080
rect 21416 35068 21422 35080
rect 21545 35071 21603 35077
rect 21545 35068 21557 35071
rect 21416 35040 21557 35068
rect 21416 35028 21422 35040
rect 21545 35037 21557 35040
rect 21591 35037 21603 35071
rect 21545 35031 21603 35037
rect 21634 35028 21640 35080
rect 21692 35068 21698 35080
rect 22097 35071 22155 35077
rect 22097 35068 22109 35071
rect 21692 35040 22109 35068
rect 21692 35028 21698 35040
rect 22097 35037 22109 35040
rect 22143 35037 22155 35071
rect 23198 35068 23204 35080
rect 23159 35040 23204 35068
rect 22097 35031 22155 35037
rect 23198 35028 23204 35040
rect 23256 35028 23262 35080
rect 23477 35071 23535 35077
rect 23477 35037 23489 35071
rect 23523 35068 23535 35071
rect 23658 35068 23664 35080
rect 23523 35040 23664 35068
rect 23523 35037 23535 35040
rect 23477 35031 23535 35037
rect 23658 35028 23664 35040
rect 23716 35028 23722 35080
rect 25130 35068 25136 35080
rect 25091 35040 25136 35068
rect 25130 35028 25136 35040
rect 25188 35028 25194 35080
rect 25409 35071 25467 35077
rect 25409 35037 25421 35071
rect 25455 35037 25467 35071
rect 25409 35031 25467 35037
rect 22278 35000 22284 35012
rect 20824 34972 22284 35000
rect 22278 34960 22284 34972
rect 22336 34960 22342 35012
rect 24854 34960 24860 35012
rect 24912 35000 24918 35012
rect 25222 35000 25228 35012
rect 24912 34972 25228 35000
rect 24912 34960 24918 34972
rect 25222 34960 25228 34972
rect 25280 35000 25286 35012
rect 25424 35000 25452 35031
rect 25498 35028 25504 35080
rect 25556 35068 25562 35080
rect 25593 35071 25651 35077
rect 25593 35068 25605 35071
rect 25556 35040 25605 35068
rect 25556 35028 25562 35040
rect 25593 35037 25605 35040
rect 25639 35068 25651 35071
rect 25774 35068 25780 35080
rect 25639 35040 25780 35068
rect 25639 35037 25651 35040
rect 25593 35031 25651 35037
rect 25774 35028 25780 35040
rect 25832 35028 25838 35080
rect 26237 35071 26295 35077
rect 26237 35037 26249 35071
rect 26283 35068 26295 35071
rect 26326 35068 26332 35080
rect 26283 35040 26332 35068
rect 26283 35037 26295 35040
rect 26237 35031 26295 35037
rect 26326 35028 26332 35040
rect 26384 35028 26390 35080
rect 26510 35068 26516 35080
rect 26471 35040 26516 35068
rect 26510 35028 26516 35040
rect 26568 35028 26574 35080
rect 26786 35028 26792 35080
rect 26844 35068 26850 35080
rect 27157 35071 27215 35077
rect 27157 35068 27169 35071
rect 26844 35040 27169 35068
rect 26844 35028 26850 35040
rect 27157 35037 27169 35040
rect 27203 35037 27215 35071
rect 27157 35031 27215 35037
rect 27430 35000 27436 35012
rect 25280 34972 27436 35000
rect 25280 34960 25286 34972
rect 27430 34960 27436 34972
rect 27488 34960 27494 35012
rect 27540 35000 27568 35108
rect 28718 35096 28724 35148
rect 28776 35136 28782 35148
rect 30285 35139 30343 35145
rect 30285 35136 30297 35139
rect 28776 35108 30297 35136
rect 28776 35096 28782 35108
rect 30285 35105 30297 35108
rect 30331 35105 30343 35139
rect 30285 35099 30343 35105
rect 27617 35071 27675 35077
rect 27617 35037 27629 35071
rect 27663 35068 27675 35071
rect 28994 35068 29000 35080
rect 27663 35040 29000 35068
rect 27663 35037 27675 35040
rect 27617 35031 27675 35037
rect 28994 35028 29000 35040
rect 29052 35028 29058 35080
rect 29089 35071 29147 35077
rect 29089 35037 29101 35071
rect 29135 35068 29147 35071
rect 29825 35071 29883 35077
rect 29825 35068 29837 35071
rect 29135 35040 29837 35068
rect 29135 35037 29147 35040
rect 29089 35031 29147 35037
rect 29825 35037 29837 35040
rect 29871 35037 29883 35071
rect 29825 35031 29883 35037
rect 30190 35028 30196 35080
rect 30248 35068 30254 35080
rect 30469 35071 30527 35077
rect 30469 35068 30481 35071
rect 30248 35040 30481 35068
rect 30248 35028 30254 35040
rect 30469 35037 30481 35040
rect 30515 35037 30527 35071
rect 30576 35068 30604 35176
rect 30745 35071 30803 35077
rect 30745 35068 30757 35071
rect 30576 35040 30757 35068
rect 30469 35031 30527 35037
rect 30745 35037 30757 35040
rect 30791 35037 30803 35071
rect 30745 35031 30803 35037
rect 30926 35028 30932 35080
rect 30984 35068 30990 35080
rect 31294 35068 31300 35080
rect 30984 35040 31300 35068
rect 30984 35028 30990 35040
rect 31294 35028 31300 35040
rect 31352 35028 31358 35080
rect 27862 35003 27920 35009
rect 27862 35000 27874 35003
rect 27540 34972 27874 35000
rect 27862 34969 27874 34972
rect 27908 34969 27920 35003
rect 27862 34963 27920 34969
rect 28074 34960 28080 35012
rect 28132 35000 28138 35012
rect 29641 35003 29699 35009
rect 29641 35000 29653 35003
rect 28132 34972 29653 35000
rect 28132 34960 28138 34972
rect 29641 34969 29653 34972
rect 29687 34969 29699 35003
rect 29641 34963 29699 34969
rect 20257 34935 20315 34941
rect 20257 34932 20269 34935
rect 20128 34904 20269 34932
rect 20128 34892 20134 34904
rect 20257 34901 20269 34904
rect 20303 34901 20315 34935
rect 20257 34895 20315 34901
rect 20346 34892 20352 34944
rect 20404 34932 20410 34944
rect 25314 34932 25320 34944
rect 20404 34904 25320 34932
rect 20404 34892 20410 34904
rect 25314 34892 25320 34904
rect 25372 34892 25378 34944
rect 26973 34935 27031 34941
rect 26973 34901 26985 34935
rect 27019 34932 27031 34935
rect 27154 34932 27160 34944
rect 27019 34904 27160 34932
rect 27019 34901 27031 34904
rect 26973 34895 27031 34901
rect 27154 34892 27160 34904
rect 27212 34892 27218 34944
rect 1104 34842 32016 34864
rect 1104 34790 7288 34842
rect 7340 34790 17592 34842
rect 17644 34790 27896 34842
rect 27948 34790 32016 34842
rect 1104 34768 32016 34790
rect 3697 34731 3755 34737
rect 3697 34697 3709 34731
rect 3743 34728 3755 34731
rect 5166 34728 5172 34740
rect 3743 34700 5028 34728
rect 5127 34700 5172 34728
rect 3743 34697 3755 34700
rect 3697 34691 3755 34697
rect 2774 34620 2780 34672
rect 2832 34660 2838 34672
rect 4034 34663 4092 34669
rect 4034 34660 4046 34663
rect 2832 34632 4046 34660
rect 2832 34620 2838 34632
rect 4034 34629 4046 34632
rect 4080 34629 4092 34663
rect 5000 34660 5028 34700
rect 5166 34688 5172 34700
rect 5224 34688 5230 34740
rect 5629 34731 5687 34737
rect 5629 34697 5641 34731
rect 5675 34728 5687 34731
rect 7006 34728 7012 34740
rect 5675 34700 7012 34728
rect 5675 34697 5687 34700
rect 5629 34691 5687 34697
rect 7006 34688 7012 34700
rect 7064 34688 7070 34740
rect 7098 34688 7104 34740
rect 7156 34728 7162 34740
rect 7745 34731 7803 34737
rect 7745 34728 7757 34731
rect 7156 34700 7757 34728
rect 7156 34688 7162 34700
rect 7745 34697 7757 34700
rect 7791 34728 7803 34731
rect 8018 34728 8024 34740
rect 7791 34700 8024 34728
rect 7791 34697 7803 34700
rect 7745 34691 7803 34697
rect 8018 34688 8024 34700
rect 8076 34688 8082 34740
rect 8389 34731 8447 34737
rect 8389 34697 8401 34731
rect 8435 34728 8447 34731
rect 10410 34728 10416 34740
rect 8435 34700 10416 34728
rect 8435 34697 8447 34700
rect 8389 34691 8447 34697
rect 10410 34688 10416 34700
rect 10468 34728 10474 34740
rect 10778 34728 10784 34740
rect 10468 34700 10784 34728
rect 10468 34688 10474 34700
rect 10778 34688 10784 34700
rect 10836 34688 10842 34740
rect 10962 34688 10968 34740
rect 11020 34728 11026 34740
rect 11793 34731 11851 34737
rect 11793 34728 11805 34731
rect 11020 34700 11805 34728
rect 11020 34688 11026 34700
rect 11793 34697 11805 34700
rect 11839 34697 11851 34731
rect 11793 34691 11851 34697
rect 11882 34688 11888 34740
rect 11940 34728 11946 34740
rect 14185 34731 14243 34737
rect 11940 34700 11985 34728
rect 11940 34688 11946 34700
rect 14185 34697 14197 34731
rect 14231 34728 14243 34731
rect 14550 34728 14556 34740
rect 14231 34700 14556 34728
rect 14231 34697 14243 34700
rect 14185 34691 14243 34697
rect 14550 34688 14556 34700
rect 14608 34688 14614 34740
rect 14737 34731 14795 34737
rect 14737 34697 14749 34731
rect 14783 34728 14795 34731
rect 15378 34728 15384 34740
rect 14783 34700 15384 34728
rect 14783 34697 14795 34700
rect 14737 34691 14795 34697
rect 15378 34688 15384 34700
rect 15436 34688 15442 34740
rect 15562 34688 15568 34740
rect 15620 34728 15626 34740
rect 17405 34731 17463 34737
rect 17405 34728 17417 34731
rect 15620 34700 17417 34728
rect 15620 34688 15626 34700
rect 17405 34697 17417 34700
rect 17451 34697 17463 34731
rect 17405 34691 17463 34697
rect 18417 34731 18475 34737
rect 18417 34697 18429 34731
rect 18463 34728 18475 34731
rect 20070 34728 20076 34740
rect 18463 34700 20076 34728
rect 18463 34697 18475 34700
rect 18417 34691 18475 34697
rect 20070 34688 20076 34700
rect 20128 34688 20134 34740
rect 21634 34688 21640 34740
rect 21692 34728 21698 34740
rect 22097 34731 22155 34737
rect 22097 34728 22109 34731
rect 21692 34700 22109 34728
rect 21692 34688 21698 34700
rect 22097 34697 22109 34700
rect 22143 34697 22155 34731
rect 28166 34728 28172 34740
rect 22097 34691 22155 34697
rect 23032 34700 28172 34728
rect 5000 34632 5672 34660
rect 4034 34623 4092 34629
rect 5644 34604 5672 34632
rect 6362 34620 6368 34672
rect 6420 34660 6426 34672
rect 6610 34663 6668 34669
rect 6610 34660 6622 34663
rect 6420 34632 6622 34660
rect 6420 34620 6426 34632
rect 6610 34629 6622 34632
rect 6656 34629 6668 34663
rect 6610 34623 6668 34629
rect 8202 34620 8208 34672
rect 8260 34660 8266 34672
rect 8297 34663 8355 34669
rect 8297 34660 8309 34663
rect 8260 34632 8309 34660
rect 8260 34620 8266 34632
rect 8297 34629 8309 34632
rect 8343 34660 8355 34663
rect 8570 34660 8576 34672
rect 8343 34632 8576 34660
rect 8343 34629 8355 34632
rect 8297 34623 8355 34629
rect 8570 34620 8576 34632
rect 8628 34620 8634 34672
rect 9858 34660 9864 34672
rect 8956 34632 9864 34660
rect 1397 34595 1455 34601
rect 1397 34561 1409 34595
rect 1443 34561 1455 34595
rect 1397 34555 1455 34561
rect 3053 34595 3111 34601
rect 3053 34561 3065 34595
rect 3099 34592 3111 34595
rect 5074 34592 5080 34604
rect 3099 34564 5080 34592
rect 3099 34561 3111 34564
rect 3053 34555 3111 34561
rect 1412 34388 1440 34555
rect 5074 34552 5080 34564
rect 5132 34552 5138 34604
rect 5626 34552 5632 34604
rect 5684 34552 5690 34604
rect 5810 34592 5816 34604
rect 5771 34564 5816 34592
rect 5810 34552 5816 34564
rect 5868 34552 5874 34604
rect 8956 34601 8984 34632
rect 9858 34620 9864 34632
rect 9916 34620 9922 34672
rect 11698 34660 11704 34672
rect 11659 34632 11704 34660
rect 11698 34620 11704 34632
rect 11756 34620 11762 34672
rect 12069 34663 12127 34669
rect 12069 34629 12081 34663
rect 12115 34660 12127 34663
rect 12250 34660 12256 34672
rect 12115 34632 12256 34660
rect 12115 34629 12127 34632
rect 12069 34623 12127 34629
rect 12250 34620 12256 34632
rect 12308 34620 12314 34672
rect 15286 34620 15292 34672
rect 15344 34660 15350 34672
rect 15344 34632 15608 34660
rect 15344 34620 15350 34632
rect 8941 34595 8999 34601
rect 8941 34561 8953 34595
rect 8987 34561 8999 34595
rect 8941 34555 8999 34561
rect 9208 34595 9266 34601
rect 9208 34561 9220 34595
rect 9254 34592 9266 34595
rect 10042 34592 10048 34604
rect 9254 34564 10048 34592
rect 9254 34561 9266 34564
rect 9208 34555 9266 34561
rect 10042 34552 10048 34564
rect 10100 34552 10106 34604
rect 13173 34595 13231 34601
rect 13173 34561 13185 34595
rect 13219 34592 13231 34595
rect 13538 34592 13544 34604
rect 13219 34564 13544 34592
rect 13219 34561 13231 34564
rect 13173 34555 13231 34561
rect 13538 34552 13544 34564
rect 13596 34552 13602 34604
rect 14001 34595 14059 34601
rect 14001 34561 14013 34595
rect 14047 34561 14059 34595
rect 14182 34592 14188 34604
rect 14143 34564 14188 34592
rect 14001 34555 14059 34561
rect 3329 34527 3387 34533
rect 3329 34493 3341 34527
rect 3375 34524 3387 34527
rect 3697 34527 3755 34533
rect 3697 34524 3709 34527
rect 3375 34496 3709 34524
rect 3375 34493 3387 34496
rect 3329 34487 3387 34493
rect 3697 34493 3709 34496
rect 3743 34493 3755 34527
rect 3697 34487 3755 34493
rect 3789 34527 3847 34533
rect 3789 34493 3801 34527
rect 3835 34493 3847 34527
rect 6362 34524 6368 34536
rect 6323 34496 6368 34524
rect 3789 34487 3847 34493
rect 2682 34416 2688 34468
rect 2740 34456 2746 34468
rect 3804 34456 3832 34487
rect 6362 34484 6368 34496
rect 6420 34484 6426 34536
rect 11517 34527 11575 34533
rect 11517 34493 11529 34527
rect 11563 34524 11575 34527
rect 12342 34524 12348 34536
rect 11563 34496 12348 34524
rect 11563 34493 11575 34496
rect 11517 34487 11575 34493
rect 12342 34484 12348 34496
rect 12400 34484 12406 34536
rect 13262 34484 13268 34536
rect 13320 34524 13326 34536
rect 13357 34527 13415 34533
rect 13357 34524 13369 34527
rect 13320 34496 13369 34524
rect 13320 34484 13326 34496
rect 13357 34493 13369 34496
rect 13403 34493 13415 34527
rect 13357 34487 13415 34493
rect 13446 34484 13452 34536
rect 13504 34524 13510 34536
rect 14016 34524 14044 34555
rect 14182 34552 14188 34564
rect 14240 34552 14246 34604
rect 14642 34592 14648 34604
rect 14603 34564 14648 34592
rect 14642 34552 14648 34564
rect 14700 34552 14706 34604
rect 14829 34595 14887 34601
rect 14829 34561 14841 34595
rect 14875 34592 14887 34595
rect 15194 34592 15200 34604
rect 14875 34564 15200 34592
rect 14875 34561 14887 34564
rect 14829 34555 14887 34561
rect 14844 34524 14872 34555
rect 15194 34552 15200 34564
rect 15252 34552 15258 34604
rect 15470 34592 15476 34604
rect 15431 34564 15476 34592
rect 15470 34552 15476 34564
rect 15528 34552 15534 34604
rect 15580 34592 15608 34632
rect 15654 34620 15660 34672
rect 15712 34660 15718 34672
rect 19521 34663 19579 34669
rect 15712 34632 19472 34660
rect 15712 34620 15718 34632
rect 16761 34595 16819 34601
rect 15580 34564 16712 34592
rect 13504 34496 13549 34524
rect 14016 34496 14872 34524
rect 13504 34484 13510 34496
rect 14918 34484 14924 34536
rect 14976 34524 14982 34536
rect 15657 34527 15715 34533
rect 15657 34524 15669 34527
rect 14976 34496 15669 34524
rect 14976 34484 14982 34496
rect 15657 34493 15669 34496
rect 15703 34493 15715 34527
rect 15657 34487 15715 34493
rect 15749 34527 15807 34533
rect 15749 34493 15761 34527
rect 15795 34524 15807 34527
rect 16298 34524 16304 34536
rect 15795 34496 16304 34524
rect 15795 34493 15807 34496
rect 15749 34487 15807 34493
rect 16298 34484 16304 34496
rect 16356 34484 16362 34536
rect 16390 34484 16396 34536
rect 16448 34524 16454 34536
rect 16684 34524 16712 34564
rect 16761 34561 16773 34595
rect 16807 34592 16819 34595
rect 17494 34592 17500 34604
rect 16807 34564 17500 34592
rect 16807 34561 16819 34564
rect 16761 34555 16819 34561
rect 17494 34552 17500 34564
rect 17552 34552 17558 34604
rect 17589 34595 17647 34601
rect 17589 34561 17601 34595
rect 17635 34592 17647 34595
rect 17954 34592 17960 34604
rect 17635 34564 17960 34592
rect 17635 34561 17647 34564
rect 17589 34555 17647 34561
rect 17954 34552 17960 34564
rect 18012 34552 18018 34604
rect 18233 34595 18291 34601
rect 18233 34561 18245 34595
rect 18279 34592 18291 34595
rect 18322 34592 18328 34604
rect 18279 34564 18328 34592
rect 18279 34561 18291 34564
rect 18233 34555 18291 34561
rect 18322 34552 18328 34564
rect 18380 34552 18386 34604
rect 18506 34592 18512 34604
rect 18467 34564 18512 34592
rect 18506 34552 18512 34564
rect 18564 34552 18570 34604
rect 19444 34592 19472 34632
rect 19521 34629 19533 34663
rect 19567 34660 19579 34663
rect 19978 34660 19984 34672
rect 19567 34632 19984 34660
rect 19567 34629 19579 34632
rect 19521 34623 19579 34629
rect 19978 34620 19984 34632
rect 20036 34660 20042 34672
rect 20622 34660 20628 34672
rect 20036 34632 20628 34660
rect 20036 34620 20042 34632
rect 20622 34620 20628 34632
rect 20680 34620 20686 34672
rect 22649 34663 22707 34669
rect 22649 34660 22661 34663
rect 20732 34632 22661 34660
rect 20732 34592 20760 34632
rect 22649 34629 22661 34632
rect 22695 34629 22707 34663
rect 22649 34623 22707 34629
rect 19444 34564 20760 34592
rect 20898 34552 20904 34604
rect 20956 34592 20962 34604
rect 22281 34595 22339 34601
rect 22281 34592 22293 34595
rect 20956 34564 22293 34592
rect 20956 34552 20962 34564
rect 22281 34561 22293 34564
rect 22327 34561 22339 34595
rect 22281 34555 22339 34561
rect 22462 34552 22468 34604
rect 22520 34592 22526 34604
rect 22925 34595 22983 34601
rect 22925 34592 22937 34595
rect 22520 34564 22937 34592
rect 22520 34552 22526 34564
rect 22925 34561 22937 34564
rect 22971 34561 22983 34595
rect 22925 34555 22983 34561
rect 21174 34524 21180 34536
rect 16448 34496 16620 34524
rect 16684 34496 21180 34524
rect 16448 34484 16454 34496
rect 2740 34428 3832 34456
rect 12989 34459 13047 34465
rect 2740 34416 2746 34428
rect 12989 34425 13001 34459
rect 13035 34456 13047 34459
rect 15930 34456 15936 34468
rect 13035 34428 15936 34456
rect 13035 34425 13047 34428
rect 12989 34419 13047 34425
rect 15930 34416 15936 34428
rect 15988 34416 15994 34468
rect 16592 34456 16620 34496
rect 21174 34484 21180 34496
rect 21232 34484 21238 34536
rect 23032 34524 23060 34700
rect 28166 34688 28172 34700
rect 28224 34688 28230 34740
rect 30374 34728 30380 34740
rect 29104 34700 30380 34728
rect 25958 34660 25964 34672
rect 23492 34632 25360 34660
rect 25919 34632 25964 34660
rect 23106 34552 23112 34604
rect 23164 34592 23170 34604
rect 23164 34564 23209 34592
rect 23164 34552 23170 34564
rect 23198 34524 23204 34536
rect 21284 34496 23060 34524
rect 23159 34496 23204 34524
rect 16945 34459 17003 34465
rect 16945 34456 16957 34459
rect 16592 34428 16957 34456
rect 16945 34425 16957 34428
rect 16991 34425 17003 34459
rect 16945 34419 17003 34425
rect 17310 34416 17316 34468
rect 17368 34456 17374 34468
rect 21284 34456 21312 34496
rect 23198 34484 23204 34496
rect 23256 34524 23262 34536
rect 23492 34524 23520 34632
rect 23658 34592 23664 34604
rect 23619 34564 23664 34592
rect 23658 34552 23664 34564
rect 23716 34552 23722 34604
rect 24857 34595 24915 34601
rect 24857 34561 24869 34595
rect 24903 34592 24915 34595
rect 25038 34592 25044 34604
rect 24903 34564 25044 34592
rect 24903 34561 24915 34564
rect 24857 34555 24915 34561
rect 25038 34552 25044 34564
rect 25096 34552 25102 34604
rect 25133 34595 25191 34601
rect 25133 34561 25145 34595
rect 25179 34592 25191 34595
rect 25222 34592 25228 34604
rect 25179 34564 25228 34592
rect 25179 34561 25191 34564
rect 25133 34555 25191 34561
rect 25222 34552 25228 34564
rect 25280 34552 25286 34604
rect 25332 34601 25360 34632
rect 25958 34620 25964 34632
rect 26016 34620 26022 34672
rect 28902 34660 28908 34672
rect 26436 34632 28908 34660
rect 25317 34595 25375 34601
rect 25317 34561 25329 34595
rect 25363 34592 25375 34595
rect 25774 34592 25780 34604
rect 25363 34564 25780 34592
rect 25363 34561 25375 34564
rect 25317 34555 25375 34561
rect 25774 34552 25780 34564
rect 25832 34552 25838 34604
rect 26145 34595 26203 34601
rect 26145 34561 26157 34595
rect 26191 34592 26203 34595
rect 26234 34592 26240 34604
rect 26191 34564 26240 34592
rect 26191 34561 26203 34564
rect 26145 34555 26203 34561
rect 26234 34552 26240 34564
rect 26292 34552 26298 34604
rect 26436 34590 26464 34632
rect 28902 34620 28908 34632
rect 28960 34620 28966 34672
rect 26344 34562 26464 34590
rect 26344 34533 26372 34562
rect 27338 34552 27344 34604
rect 27396 34590 27402 34604
rect 27433 34595 27491 34601
rect 27433 34590 27445 34595
rect 27396 34562 27445 34590
rect 27396 34552 27402 34562
rect 27433 34561 27445 34562
rect 27479 34561 27491 34595
rect 28353 34595 28411 34601
rect 28353 34592 28365 34595
rect 27433 34555 27491 34561
rect 27632 34564 28365 34592
rect 23256 34496 23520 34524
rect 26329 34527 26387 34533
rect 23256 34484 23262 34496
rect 26329 34493 26341 34527
rect 26375 34493 26387 34527
rect 26329 34487 26387 34493
rect 26421 34527 26479 34533
rect 26421 34493 26433 34527
rect 26467 34493 26479 34527
rect 26421 34487 26479 34493
rect 27157 34527 27215 34533
rect 27157 34493 27169 34527
rect 27203 34524 27215 34527
rect 27632 34524 27660 34564
rect 28353 34561 28365 34564
rect 28399 34561 28411 34595
rect 28353 34555 28411 34561
rect 28442 34552 28448 34604
rect 28500 34592 28506 34604
rect 28537 34595 28595 34601
rect 28537 34592 28549 34595
rect 28500 34564 28549 34592
rect 28500 34552 28506 34564
rect 28537 34561 28549 34564
rect 28583 34561 28595 34595
rect 28537 34555 28595 34561
rect 29104 34524 29132 34700
rect 30374 34688 30380 34700
rect 30432 34728 30438 34740
rect 30834 34728 30840 34740
rect 30432 34700 30840 34728
rect 30432 34688 30438 34700
rect 30834 34688 30840 34700
rect 30892 34728 30898 34740
rect 30892 34700 31156 34728
rect 30892 34688 30898 34700
rect 29472 34632 30972 34660
rect 29270 34552 29276 34604
rect 29328 34592 29334 34604
rect 29472 34601 29500 34632
rect 29457 34595 29515 34601
rect 29457 34592 29469 34595
rect 29328 34564 29469 34592
rect 29328 34552 29334 34564
rect 29457 34561 29469 34564
rect 29503 34561 29515 34595
rect 29457 34555 29515 34561
rect 29730 34552 29736 34604
rect 29788 34592 29794 34604
rect 30190 34592 30196 34604
rect 29788 34564 30196 34592
rect 29788 34552 29794 34564
rect 30190 34552 30196 34564
rect 30248 34592 30254 34604
rect 30944 34601 30972 34632
rect 31128 34601 31156 34700
rect 30653 34595 30711 34601
rect 30653 34592 30665 34595
rect 30248 34564 30665 34592
rect 30248 34552 30254 34564
rect 30653 34561 30665 34564
rect 30699 34561 30711 34595
rect 30653 34555 30711 34561
rect 30929 34595 30987 34601
rect 30929 34561 30941 34595
rect 30975 34561 30987 34595
rect 30929 34555 30987 34561
rect 31113 34595 31171 34601
rect 31113 34561 31125 34595
rect 31159 34561 31171 34595
rect 31113 34555 31171 34561
rect 27203 34496 27660 34524
rect 27724 34496 29132 34524
rect 29181 34527 29239 34533
rect 27203 34493 27215 34496
rect 27157 34487 27215 34493
rect 22186 34456 22192 34468
rect 17368 34428 21312 34456
rect 22066 34428 22192 34456
rect 17368 34416 17374 34428
rect 1578 34388 1584 34400
rect 860 34360 1440 34388
rect 1539 34360 1584 34388
rect 860 33980 888 34360
rect 1578 34348 1584 34360
rect 1636 34348 1642 34400
rect 2866 34388 2872 34400
rect 2827 34360 2872 34388
rect 2866 34348 2872 34360
rect 2924 34348 2930 34400
rect 3142 34348 3148 34400
rect 3200 34388 3206 34400
rect 3237 34391 3295 34397
rect 3237 34388 3249 34391
rect 3200 34360 3249 34388
rect 3200 34348 3206 34360
rect 3237 34357 3249 34360
rect 3283 34357 3295 34391
rect 3237 34351 3295 34357
rect 10321 34391 10379 34397
rect 10321 34357 10333 34391
rect 10367 34388 10379 34391
rect 10410 34388 10416 34400
rect 10367 34360 10416 34388
rect 10367 34357 10379 34360
rect 10321 34351 10379 34357
rect 10410 34348 10416 34360
rect 10468 34348 10474 34400
rect 15289 34391 15347 34397
rect 15289 34357 15301 34391
rect 15335 34388 15347 34391
rect 15378 34388 15384 34400
rect 15335 34360 15384 34388
rect 15335 34357 15347 34360
rect 15289 34351 15347 34357
rect 15378 34348 15384 34360
rect 15436 34348 15442 34400
rect 18233 34391 18291 34397
rect 18233 34357 18245 34391
rect 18279 34388 18291 34391
rect 18414 34388 18420 34400
rect 18279 34360 18420 34388
rect 18279 34357 18291 34360
rect 18233 34351 18291 34357
rect 18414 34348 18420 34360
rect 18472 34348 18478 34400
rect 19334 34348 19340 34400
rect 19392 34388 19398 34400
rect 20530 34388 20536 34400
rect 19392 34360 20536 34388
rect 19392 34348 19398 34360
rect 20530 34348 20536 34360
rect 20588 34388 20594 34400
rect 20809 34391 20867 34397
rect 20809 34388 20821 34391
rect 20588 34360 20821 34388
rect 20588 34348 20594 34360
rect 20809 34357 20821 34360
rect 20855 34388 20867 34391
rect 22066 34388 22094 34428
rect 22186 34416 22192 34428
rect 22244 34416 22250 34468
rect 22649 34459 22707 34465
rect 22649 34425 22661 34459
rect 22695 34456 22707 34459
rect 23842 34456 23848 34468
rect 22695 34428 23848 34456
rect 22695 34425 22707 34428
rect 22649 34419 22707 34425
rect 23842 34416 23848 34428
rect 23900 34416 23906 34468
rect 26436 34456 26464 34487
rect 27724 34456 27752 34496
rect 29181 34493 29193 34527
rect 29227 34493 29239 34527
rect 29181 34487 29239 34493
rect 26436 34428 27752 34456
rect 28353 34459 28411 34465
rect 28353 34425 28365 34459
rect 28399 34456 28411 34459
rect 28721 34459 28779 34465
rect 28721 34456 28733 34459
rect 28399 34428 28733 34456
rect 28399 34425 28411 34428
rect 28353 34419 28411 34425
rect 28721 34425 28733 34428
rect 28767 34456 28779 34459
rect 29196 34456 29224 34487
rect 29546 34484 29552 34536
rect 29604 34524 29610 34536
rect 30469 34527 30527 34533
rect 30469 34524 30481 34527
rect 29604 34496 30481 34524
rect 29604 34484 29610 34496
rect 30469 34493 30481 34496
rect 30515 34493 30527 34527
rect 30469 34487 30527 34493
rect 29822 34456 29828 34468
rect 28767 34428 29828 34456
rect 28767 34425 28779 34428
rect 28721 34419 28779 34425
rect 29822 34416 29828 34428
rect 29880 34456 29886 34468
rect 30742 34456 30748 34468
rect 29880 34428 30748 34456
rect 29880 34416 29886 34428
rect 30742 34416 30748 34428
rect 30800 34416 30806 34468
rect 20855 34360 22094 34388
rect 20855 34357 20867 34360
rect 20809 34351 20867 34357
rect 22370 34348 22376 34400
rect 22428 34388 22434 34400
rect 22741 34391 22799 34397
rect 22741 34388 22753 34391
rect 22428 34360 22753 34388
rect 22428 34348 22434 34360
rect 22741 34357 22753 34360
rect 22787 34357 22799 34391
rect 22741 34351 22799 34357
rect 23566 34348 23572 34400
rect 23624 34388 23630 34400
rect 23753 34391 23811 34397
rect 23753 34388 23765 34391
rect 23624 34360 23765 34388
rect 23624 34348 23630 34360
rect 23753 34357 23765 34360
rect 23799 34357 23811 34391
rect 23753 34351 23811 34357
rect 24673 34391 24731 34397
rect 24673 34357 24685 34391
rect 24719 34388 24731 34391
rect 24762 34388 24768 34400
rect 24719 34360 24768 34388
rect 24719 34357 24731 34360
rect 24673 34351 24731 34357
rect 24762 34348 24768 34360
rect 24820 34348 24826 34400
rect 1104 34298 32016 34320
rect 1104 34246 2136 34298
rect 2188 34246 12440 34298
rect 12492 34246 22744 34298
rect 22796 34246 32016 34298
rect 1104 34224 32016 34246
rect 1857 34187 1915 34193
rect 1857 34153 1869 34187
rect 1903 34184 1915 34187
rect 1946 34184 1952 34196
rect 1903 34156 1952 34184
rect 1903 34153 1915 34156
rect 1857 34147 1915 34153
rect 1946 34144 1952 34156
rect 2004 34144 2010 34196
rect 2222 34184 2228 34196
rect 2183 34156 2228 34184
rect 2222 34144 2228 34156
rect 2280 34144 2286 34196
rect 5718 34144 5724 34196
rect 5776 34184 5782 34196
rect 5905 34187 5963 34193
rect 5905 34184 5917 34187
rect 5776 34156 5917 34184
rect 5776 34144 5782 34156
rect 5905 34153 5917 34156
rect 5951 34184 5963 34187
rect 6822 34184 6828 34196
rect 5951 34156 6828 34184
rect 5951 34153 5963 34156
rect 5905 34147 5963 34153
rect 6822 34144 6828 34156
rect 6880 34144 6886 34196
rect 8941 34187 8999 34193
rect 8941 34153 8953 34187
rect 8987 34184 8999 34187
rect 9122 34184 9128 34196
rect 8987 34156 9128 34184
rect 8987 34153 8999 34156
rect 8941 34147 8999 34153
rect 9122 34144 9128 34156
rect 9180 34144 9186 34196
rect 10042 34184 10048 34196
rect 10003 34156 10048 34184
rect 10042 34144 10048 34156
rect 10100 34144 10106 34196
rect 10686 34144 10692 34196
rect 10744 34184 10750 34196
rect 11701 34187 11759 34193
rect 11701 34184 11713 34187
rect 10744 34156 11713 34184
rect 10744 34144 10750 34156
rect 11701 34153 11713 34156
rect 11747 34153 11759 34187
rect 11701 34147 11759 34153
rect 14645 34187 14703 34193
rect 14645 34153 14657 34187
rect 14691 34184 14703 34187
rect 14918 34184 14924 34196
rect 14691 34156 14924 34184
rect 14691 34153 14703 34156
rect 14645 34147 14703 34153
rect 14918 34144 14924 34156
rect 14976 34144 14982 34196
rect 15197 34187 15255 34193
rect 15197 34153 15209 34187
rect 15243 34184 15255 34187
rect 15470 34184 15476 34196
rect 15243 34156 15476 34184
rect 15243 34153 15255 34156
rect 15197 34147 15255 34153
rect 15470 34144 15476 34156
rect 15528 34144 15534 34196
rect 18601 34187 18659 34193
rect 18601 34153 18613 34187
rect 18647 34184 18659 34187
rect 20717 34187 20775 34193
rect 18647 34156 20668 34184
rect 18647 34153 18659 34156
rect 18601 34147 18659 34153
rect 17681 34119 17739 34125
rect 17681 34116 17693 34119
rect 11992 34088 17693 34116
rect 2317 34051 2375 34057
rect 2317 34017 2329 34051
rect 2363 34048 2375 34051
rect 2498 34048 2504 34060
rect 2363 34020 2504 34048
rect 2363 34017 2375 34020
rect 2317 34011 2375 34017
rect 2498 34008 2504 34020
rect 2556 34008 2562 34060
rect 2774 34008 2780 34060
rect 2832 34048 2838 34060
rect 3142 34048 3148 34060
rect 2832 34020 3148 34048
rect 2832 34008 2838 34020
rect 3142 34008 3148 34020
rect 3200 34008 3206 34060
rect 6362 34008 6368 34060
rect 6420 34048 6426 34060
rect 6917 34051 6975 34057
rect 6917 34048 6929 34051
rect 6420 34020 6929 34048
rect 6420 34008 6426 34020
rect 6917 34017 6929 34020
rect 6963 34017 6975 34051
rect 6917 34011 6975 34017
rect 8110 34008 8116 34060
rect 8168 34048 8174 34060
rect 10413 34051 10471 34057
rect 10413 34048 10425 34051
rect 8168 34020 10425 34048
rect 8168 34008 8174 34020
rect 10413 34017 10425 34020
rect 10459 34017 10471 34051
rect 10413 34011 10471 34017
rect 768 33952 888 33980
rect 2041 33983 2099 33989
rect 768 33708 796 33952
rect 2041 33949 2053 33983
rect 2087 33949 2099 33983
rect 2958 33980 2964 33992
rect 2919 33952 2964 33980
rect 2041 33943 2099 33949
rect 2056 33912 2084 33943
rect 2958 33940 2964 33952
rect 3016 33940 3022 33992
rect 3234 33980 3240 33992
rect 3195 33952 3240 33980
rect 3234 33940 3240 33952
rect 3292 33940 3298 33992
rect 4430 33940 4436 33992
rect 4488 33980 4494 33992
rect 4525 33983 4583 33989
rect 4525 33980 4537 33983
rect 4488 33952 4537 33980
rect 4488 33940 4494 33952
rect 4525 33949 4537 33952
rect 4571 33980 4583 33983
rect 6380 33980 6408 34008
rect 11992 33992 12020 34088
rect 17681 34085 17693 34088
rect 17727 34116 17739 34119
rect 18506 34116 18512 34128
rect 17727 34088 18512 34116
rect 17727 34085 17739 34088
rect 17681 34079 17739 34085
rect 18506 34076 18512 34088
rect 18564 34076 18570 34128
rect 20640 34116 20668 34156
rect 20717 34153 20729 34187
rect 20763 34184 20775 34187
rect 21726 34184 21732 34196
rect 20763 34156 21732 34184
rect 20763 34153 20775 34156
rect 20717 34147 20775 34153
rect 21726 34144 21732 34156
rect 21784 34144 21790 34196
rect 23477 34187 23535 34193
rect 23477 34153 23489 34187
rect 23523 34184 23535 34187
rect 23658 34184 23664 34196
rect 23523 34156 23664 34184
rect 23523 34153 23535 34156
rect 23477 34147 23535 34153
rect 23658 34144 23664 34156
rect 23716 34144 23722 34196
rect 25774 34184 25780 34196
rect 25735 34156 25780 34184
rect 25774 34144 25780 34156
rect 25832 34144 25838 34196
rect 28994 34184 29000 34196
rect 26344 34156 29000 34184
rect 20806 34116 20812 34128
rect 20640 34088 20812 34116
rect 20806 34076 20812 34088
rect 20864 34116 20870 34128
rect 21545 34119 21603 34125
rect 21545 34116 21557 34119
rect 20864 34088 21557 34116
rect 20864 34076 20870 34088
rect 21545 34085 21557 34088
rect 21591 34085 21603 34119
rect 21545 34079 21603 34085
rect 14737 34051 14795 34057
rect 14737 34017 14749 34051
rect 14783 34048 14795 34051
rect 16298 34048 16304 34060
rect 14783 34020 15884 34048
rect 16259 34020 16304 34048
rect 14783 34017 14795 34020
rect 14737 34011 14795 34017
rect 4571 33952 6408 33980
rect 4571 33949 4583 33952
rect 4525 33943 4583 33949
rect 7926 33940 7932 33992
rect 7984 33980 7990 33992
rect 9122 33980 9128 33992
rect 7984 33952 9128 33980
rect 7984 33940 7990 33952
rect 9122 33940 9128 33952
rect 9180 33940 9186 33992
rect 9398 33980 9404 33992
rect 9359 33952 9404 33980
rect 9398 33940 9404 33952
rect 9456 33940 9462 33992
rect 9585 33983 9643 33989
rect 9585 33949 9597 33983
rect 9631 33949 9643 33983
rect 10226 33980 10232 33992
rect 10187 33952 10232 33980
rect 9585 33943 9643 33949
rect 2406 33912 2412 33924
rect 2056 33884 2412 33912
rect 2406 33872 2412 33884
rect 2464 33872 2470 33924
rect 2866 33872 2872 33924
rect 2924 33912 2930 33924
rect 4770 33915 4828 33921
rect 4770 33912 4782 33915
rect 2924 33884 4782 33912
rect 2924 33872 2930 33884
rect 4770 33881 4782 33884
rect 4816 33881 4828 33915
rect 4770 33875 4828 33881
rect 7184 33915 7242 33921
rect 7184 33881 7196 33915
rect 7230 33912 7242 33915
rect 7558 33912 7564 33924
rect 7230 33884 7564 33912
rect 7230 33881 7242 33884
rect 7184 33875 7242 33881
rect 7558 33872 7564 33884
rect 7616 33872 7622 33924
rect 9214 33872 9220 33924
rect 9272 33912 9278 33924
rect 9600 33912 9628 33943
rect 10226 33940 10232 33952
rect 10284 33940 10290 33992
rect 10505 33983 10563 33989
rect 10505 33949 10517 33983
rect 10551 33949 10563 33983
rect 11054 33980 11060 33992
rect 11015 33952 11060 33980
rect 10505 33943 10563 33949
rect 10520 33912 10548 33943
rect 11054 33940 11060 33952
rect 11112 33940 11118 33992
rect 11149 33983 11207 33989
rect 11149 33949 11161 33983
rect 11195 33980 11207 33983
rect 11882 33980 11888 33992
rect 11195 33952 11888 33980
rect 11195 33949 11207 33952
rect 11149 33943 11207 33949
rect 11882 33940 11888 33952
rect 11940 33940 11946 33992
rect 11974 33940 11980 33992
rect 12032 33980 12038 33992
rect 12986 33980 12992 33992
rect 12032 33952 12077 33980
rect 12899 33952 12992 33980
rect 12032 33940 12038 33952
rect 12986 33940 12992 33952
rect 13044 33980 13050 33992
rect 14182 33980 14188 33992
rect 13044 33952 14188 33980
rect 13044 33940 13050 33952
rect 14182 33940 14188 33952
rect 14240 33940 14246 33992
rect 14458 33980 14464 33992
rect 14419 33952 14464 33980
rect 14458 33940 14464 33952
rect 14516 33940 14522 33992
rect 15381 33983 15439 33989
rect 15381 33949 15393 33983
rect 15427 33980 15439 33983
rect 15470 33980 15476 33992
rect 15427 33952 15476 33980
rect 15427 33949 15439 33952
rect 15381 33943 15439 33949
rect 15470 33940 15476 33952
rect 15528 33940 15534 33992
rect 15654 33980 15660 33992
rect 15615 33952 15660 33980
rect 15654 33940 15660 33952
rect 15712 33940 15718 33992
rect 15856 33989 15884 34020
rect 16298 34008 16304 34020
rect 16356 34008 16362 34060
rect 18690 34048 18696 34060
rect 18651 34020 18696 34048
rect 18690 34008 18696 34020
rect 18748 34008 18754 34060
rect 26344 34057 26372 34156
rect 28994 34144 29000 34156
rect 29052 34144 29058 34196
rect 31021 34187 31079 34193
rect 31021 34184 31033 34187
rect 29104 34156 31033 34184
rect 28534 34116 28540 34128
rect 28495 34088 28540 34116
rect 28534 34076 28540 34088
rect 28592 34076 28598 34128
rect 28902 34116 28908 34128
rect 28863 34088 28908 34116
rect 28902 34076 28908 34088
rect 28960 34116 28966 34128
rect 29104 34116 29132 34156
rect 31021 34153 31033 34156
rect 31067 34153 31079 34187
rect 31021 34147 31079 34153
rect 28960 34088 29132 34116
rect 28960 34076 28966 34088
rect 21637 34051 21695 34057
rect 21637 34048 21649 34051
rect 20640 34020 21649 34048
rect 15841 33983 15899 33989
rect 15841 33949 15853 33983
rect 15887 33980 15899 33983
rect 15930 33980 15936 33992
rect 15887 33952 15936 33980
rect 15887 33949 15899 33952
rect 15841 33943 15899 33949
rect 15930 33940 15936 33952
rect 15988 33940 15994 33992
rect 16482 33980 16488 33992
rect 16443 33952 16488 33980
rect 16482 33940 16488 33952
rect 16540 33940 16546 33992
rect 18414 33980 18420 33992
rect 18375 33952 18420 33980
rect 18414 33940 18420 33952
rect 18472 33940 18478 33992
rect 19334 33980 19340 33992
rect 19295 33952 19340 33980
rect 19334 33940 19340 33952
rect 19392 33940 19398 33992
rect 20162 33940 20168 33992
rect 20220 33980 20226 33992
rect 20640 33980 20668 34020
rect 21637 34017 21649 34020
rect 21683 34017 21695 34051
rect 21637 34011 21695 34017
rect 26329 34051 26387 34057
rect 26329 34017 26341 34051
rect 26375 34017 26387 34051
rect 26329 34011 26387 34017
rect 29270 34008 29276 34060
rect 29328 34048 29334 34060
rect 29328 34020 30052 34048
rect 29328 34008 29334 34020
rect 21358 33980 21364 33992
rect 20220 33952 20668 33980
rect 21319 33952 21364 33980
rect 20220 33940 20226 33952
rect 21358 33940 21364 33952
rect 21416 33940 21422 33992
rect 22097 33983 22155 33989
rect 22097 33949 22109 33983
rect 22143 33980 22155 33983
rect 22186 33980 22192 33992
rect 22143 33952 22192 33980
rect 22143 33949 22155 33952
rect 22097 33943 22155 33949
rect 22186 33940 22192 33952
rect 22244 33940 22250 33992
rect 22370 33989 22376 33992
rect 22364 33980 22376 33989
rect 22331 33952 22376 33980
rect 22364 33943 22376 33952
rect 22370 33940 22376 33943
rect 22428 33940 22434 33992
rect 24397 33983 24455 33989
rect 24397 33949 24409 33983
rect 24443 33980 24455 33983
rect 24946 33980 24952 33992
rect 24443 33952 24952 33980
rect 24443 33949 24455 33952
rect 24397 33943 24455 33949
rect 24946 33940 24952 33952
rect 25004 33940 25010 33992
rect 25774 33940 25780 33992
rect 25832 33980 25838 33992
rect 26585 33983 26643 33989
rect 26585 33980 26597 33983
rect 25832 33952 26597 33980
rect 25832 33940 25838 33952
rect 26585 33949 26597 33952
rect 26631 33949 26643 33983
rect 28718 33980 28724 33992
rect 28679 33952 28724 33980
rect 26585 33943 26643 33949
rect 28718 33940 28724 33952
rect 28776 33940 28782 33992
rect 28997 33983 29055 33989
rect 28997 33949 29009 33983
rect 29043 33980 29055 33983
rect 29454 33980 29460 33992
rect 29043 33952 29460 33980
rect 29043 33949 29055 33952
rect 28997 33943 29055 33949
rect 29454 33940 29460 33952
rect 29512 33940 29518 33992
rect 29730 33980 29736 33992
rect 29691 33952 29736 33980
rect 29730 33940 29736 33952
rect 29788 33940 29794 33992
rect 30024 33989 30052 34020
rect 30009 33983 30067 33989
rect 30009 33949 30021 33983
rect 30055 33980 30067 33983
rect 30098 33980 30104 33992
rect 30055 33952 30104 33980
rect 30055 33949 30067 33952
rect 30009 33943 30067 33949
rect 30098 33940 30104 33952
rect 30156 33940 30162 33992
rect 30190 33940 30196 33992
rect 30248 33980 30254 33992
rect 30834 33980 30840 33992
rect 30248 33952 30293 33980
rect 30795 33952 30840 33980
rect 30248 33940 30254 33952
rect 30834 33940 30840 33952
rect 30892 33940 30898 33992
rect 31110 33980 31116 33992
rect 31071 33952 31116 33980
rect 31110 33940 31116 33952
rect 31168 33940 31174 33992
rect 11698 33912 11704 33924
rect 9272 33884 10548 33912
rect 11659 33884 11704 33912
rect 9272 33872 9278 33884
rect 11698 33872 11704 33884
rect 11756 33872 11762 33924
rect 13173 33915 13231 33921
rect 13173 33881 13185 33915
rect 13219 33912 13231 33915
rect 13354 33912 13360 33924
rect 13219 33884 13360 33912
rect 13219 33881 13231 33884
rect 13173 33875 13231 33881
rect 13354 33872 13360 33884
rect 13412 33872 13418 33924
rect 16574 33872 16580 33924
rect 16632 33912 16638 33924
rect 17497 33915 17555 33921
rect 17497 33912 17509 33915
rect 16632 33884 17509 33912
rect 16632 33872 16638 33884
rect 17497 33881 17509 33884
rect 17543 33881 17555 33915
rect 17497 33875 17555 33881
rect 19604 33915 19662 33921
rect 19604 33881 19616 33915
rect 19650 33912 19662 33915
rect 21177 33915 21235 33921
rect 21177 33912 21189 33915
rect 19650 33884 21189 33912
rect 19650 33881 19662 33884
rect 19604 33875 19662 33881
rect 21177 33881 21189 33884
rect 21223 33881 21235 33915
rect 21177 33875 21235 33881
rect 22002 33872 22008 33924
rect 22060 33912 22066 33924
rect 24670 33921 24676 33924
rect 22060 33884 24624 33912
rect 22060 33872 22066 33884
rect 2777 33847 2835 33853
rect 2777 33813 2789 33847
rect 2823 33844 2835 33847
rect 3326 33844 3332 33856
rect 2823 33816 3332 33844
rect 2823 33813 2835 33816
rect 2777 33807 2835 33813
rect 3326 33804 3332 33816
rect 3384 33804 3390 33856
rect 8294 33844 8300 33856
rect 8207 33816 8300 33844
rect 8294 33804 8300 33816
rect 8352 33844 8358 33856
rect 8938 33844 8944 33856
rect 8352 33816 8944 33844
rect 8352 33804 8358 33816
rect 8938 33804 8944 33816
rect 8996 33804 9002 33856
rect 12158 33804 12164 33856
rect 12216 33844 12222 33856
rect 13446 33844 13452 33856
rect 12216 33816 13452 33844
rect 12216 33804 12222 33816
rect 13446 33804 13452 33816
rect 13504 33804 13510 33856
rect 14274 33844 14280 33856
rect 14235 33816 14280 33844
rect 14274 33804 14280 33816
rect 14332 33804 14338 33856
rect 15746 33804 15752 33856
rect 15804 33844 15810 33856
rect 16669 33847 16727 33853
rect 16669 33844 16681 33847
rect 15804 33816 16681 33844
rect 15804 33804 15810 33816
rect 16669 33813 16681 33816
rect 16715 33813 16727 33847
rect 16669 33807 16727 33813
rect 18233 33847 18291 33853
rect 18233 33813 18245 33847
rect 18279 33844 18291 33847
rect 18782 33844 18788 33856
rect 18279 33816 18788 33844
rect 18279 33813 18291 33816
rect 18233 33807 18291 33813
rect 18782 33804 18788 33816
rect 18840 33804 18846 33856
rect 22094 33804 22100 33856
rect 22152 33844 22158 33856
rect 22370 33844 22376 33856
rect 22152 33816 22376 33844
rect 22152 33804 22158 33816
rect 22370 33804 22376 33816
rect 22428 33804 22434 33856
rect 24596 33844 24624 33884
rect 24664 33875 24676 33921
rect 24728 33912 24734 33924
rect 24728 33884 24764 33912
rect 24872 33884 26556 33912
rect 24670 33872 24676 33875
rect 24728 33872 24734 33884
rect 24872 33844 24900 33884
rect 24596 33816 24900 33844
rect 26528 33844 26556 33884
rect 26896 33884 32352 33912
rect 26896 33844 26924 33884
rect 26528 33816 26924 33844
rect 27709 33847 27767 33853
rect 27709 33813 27721 33847
rect 27755 33844 27767 33847
rect 27798 33844 27804 33856
rect 27755 33816 27804 33844
rect 27755 33813 27767 33816
rect 27709 33807 27767 33813
rect 27798 33804 27804 33816
rect 27856 33804 27862 33856
rect 28718 33804 28724 33856
rect 28776 33844 28782 33856
rect 29549 33847 29607 33853
rect 29549 33844 29561 33847
rect 28776 33816 29561 33844
rect 28776 33804 28782 33816
rect 29549 33813 29561 33816
rect 29595 33813 29607 33847
rect 29549 33807 29607 33813
rect 30190 33804 30196 33856
rect 30248 33844 30254 33856
rect 30653 33847 30711 33853
rect 30653 33844 30665 33847
rect 30248 33816 30665 33844
rect 30248 33804 30254 33816
rect 30653 33813 30665 33816
rect 30699 33813 30711 33847
rect 30653 33807 30711 33813
rect 1104 33754 32016 33776
rect 768 33680 888 33708
rect 1104 33702 7288 33754
rect 7340 33702 17592 33754
rect 17644 33702 27896 33754
rect 27948 33702 32016 33754
rect 32324 33708 32352 33884
rect 1104 33680 32016 33702
rect 32232 33680 32352 33708
rect 0 33572 800 33586
rect 860 33572 888 33680
rect 5074 33640 5080 33652
rect 5035 33612 5080 33640
rect 5074 33600 5080 33612
rect 5132 33600 5138 33652
rect 7558 33640 7564 33652
rect 7519 33612 7564 33640
rect 7558 33600 7564 33612
rect 7616 33600 7622 33652
rect 8757 33643 8815 33649
rect 8757 33609 8769 33643
rect 8803 33640 8815 33643
rect 10226 33640 10232 33652
rect 8803 33612 10232 33640
rect 8803 33609 8815 33612
rect 8757 33603 8815 33609
rect 10226 33600 10232 33612
rect 10284 33600 10290 33652
rect 11698 33600 11704 33652
rect 11756 33600 11762 33652
rect 12805 33643 12863 33649
rect 12805 33640 12817 33643
rect 12406 33612 12817 33640
rect 2682 33572 2688 33584
rect 0 33544 888 33572
rect 1412 33544 2688 33572
rect 0 33530 800 33544
rect 1412 33516 1440 33544
rect 2682 33532 2688 33544
rect 2740 33572 2746 33584
rect 4430 33572 4436 33584
rect 2740 33544 4436 33572
rect 2740 33532 2746 33544
rect 1394 33504 1400 33516
rect 1355 33476 1400 33504
rect 1394 33464 1400 33476
rect 1452 33464 1458 33516
rect 1670 33513 1676 33516
rect 1664 33467 1676 33513
rect 1728 33504 1734 33516
rect 3252 33513 3280 33544
rect 4430 33532 4436 33544
rect 4488 33532 4494 33584
rect 5442 33532 5448 33584
rect 5500 33572 5506 33584
rect 7009 33575 7067 33581
rect 7009 33572 7021 33575
rect 5500 33544 7021 33572
rect 5500 33532 5506 33544
rect 7009 33541 7021 33544
rect 7055 33541 7067 33575
rect 10410 33572 10416 33584
rect 7009 33535 7067 33541
rect 9416 33544 10416 33572
rect 3237 33507 3295 33513
rect 1728 33476 1764 33504
rect 1670 33464 1676 33467
rect 1728 33464 1734 33476
rect 3237 33473 3249 33507
rect 3283 33473 3295 33507
rect 3237 33467 3295 33473
rect 3326 33464 3332 33516
rect 3384 33504 3390 33516
rect 3493 33507 3551 33513
rect 3493 33504 3505 33507
rect 3384 33476 3505 33504
rect 3384 33464 3390 33476
rect 3493 33473 3505 33476
rect 3539 33473 3551 33507
rect 3493 33467 3551 33473
rect 5261 33507 5319 33513
rect 5261 33473 5273 33507
rect 5307 33504 5319 33507
rect 5350 33504 5356 33516
rect 5307 33476 5356 33504
rect 5307 33473 5319 33476
rect 5261 33467 5319 33473
rect 5350 33464 5356 33476
rect 5408 33464 5414 33516
rect 5537 33507 5595 33513
rect 5537 33504 5549 33507
rect 5460 33476 5549 33504
rect 4706 33328 4712 33380
rect 4764 33368 4770 33380
rect 5460 33368 5488 33476
rect 5537 33473 5549 33476
rect 5583 33473 5595 33507
rect 5718 33504 5724 33516
rect 5679 33476 5724 33504
rect 5537 33467 5595 33473
rect 5718 33464 5724 33476
rect 5776 33464 5782 33516
rect 6730 33464 6736 33516
rect 6788 33504 6794 33516
rect 6825 33507 6883 33513
rect 6825 33504 6837 33507
rect 6788 33476 6837 33504
rect 6788 33464 6794 33476
rect 6825 33473 6837 33476
rect 6871 33473 6883 33507
rect 6825 33467 6883 33473
rect 7101 33507 7159 33513
rect 7101 33473 7113 33507
rect 7147 33504 7159 33507
rect 7466 33504 7472 33516
rect 7147 33476 7472 33504
rect 7147 33473 7159 33476
rect 7101 33467 7159 33473
rect 7466 33464 7472 33476
rect 7524 33464 7530 33516
rect 7742 33504 7748 33516
rect 7703 33476 7748 33504
rect 7742 33464 7748 33476
rect 7800 33464 7806 33516
rect 8018 33504 8024 33516
rect 7979 33476 8024 33504
rect 8018 33464 8024 33476
rect 8076 33464 8082 33516
rect 8941 33507 8999 33513
rect 8941 33473 8953 33507
rect 8987 33504 8999 33507
rect 9122 33504 9128 33516
rect 8987 33476 9128 33504
rect 8987 33473 8999 33476
rect 8941 33467 8999 33473
rect 9122 33464 9128 33476
rect 9180 33464 9186 33516
rect 9217 33507 9275 33513
rect 9217 33473 9229 33507
rect 9263 33504 9275 33507
rect 9306 33504 9312 33516
rect 9263 33476 9312 33504
rect 9263 33473 9275 33476
rect 9217 33467 9275 33473
rect 9306 33464 9312 33476
rect 9364 33464 9370 33516
rect 9416 33513 9444 33544
rect 10410 33532 10416 33544
rect 10468 33532 10474 33584
rect 11517 33575 11575 33581
rect 11517 33541 11529 33575
rect 11563 33572 11575 33575
rect 11716 33572 11744 33600
rect 12406 33572 12434 33612
rect 12805 33609 12817 33612
rect 12851 33640 12863 33643
rect 12851 33612 14403 33640
rect 12851 33609 12863 33612
rect 12805 33603 12863 33609
rect 13440 33575 13498 33581
rect 11563 33544 12434 33572
rect 12544 33544 13400 33572
rect 11563 33541 11575 33544
rect 11517 33535 11575 33541
rect 9401 33507 9459 33513
rect 9401 33473 9413 33507
rect 9447 33473 9459 33507
rect 9401 33467 9459 33473
rect 10321 33507 10379 33513
rect 10321 33473 10333 33507
rect 10367 33504 10379 33507
rect 10686 33504 10692 33516
rect 10367 33476 10692 33504
rect 10367 33473 10379 33476
rect 10321 33467 10379 33473
rect 10686 33464 10692 33476
rect 10744 33464 10750 33516
rect 10965 33507 11023 33513
rect 10965 33473 10977 33507
rect 11011 33473 11023 33507
rect 11698 33504 11704 33516
rect 11659 33476 11704 33504
rect 10965 33467 11023 33473
rect 7834 33396 7840 33448
rect 7892 33436 7898 33448
rect 7929 33439 7987 33445
rect 7929 33436 7941 33439
rect 7892 33408 7941 33436
rect 7892 33396 7898 33408
rect 7929 33405 7941 33408
rect 7975 33436 7987 33439
rect 8110 33436 8116 33448
rect 7975 33408 8116 33436
rect 7975 33405 7987 33408
rect 7929 33399 7987 33405
rect 8110 33396 8116 33408
rect 8168 33396 8174 33448
rect 9950 33396 9956 33448
rect 10008 33436 10014 33448
rect 10980 33436 11008 33467
rect 11698 33464 11704 33476
rect 11756 33464 11762 33516
rect 11793 33507 11851 33513
rect 11793 33473 11805 33507
rect 11839 33504 11851 33507
rect 11974 33504 11980 33516
rect 11839 33476 11980 33504
rect 11839 33473 11851 33476
rect 11793 33467 11851 33473
rect 11974 33464 11980 33476
rect 12032 33464 12038 33516
rect 12544 33513 12572 33544
rect 12529 33507 12587 33513
rect 12529 33473 12541 33507
rect 12575 33473 12587 33507
rect 12529 33467 12587 33473
rect 12713 33507 12771 33513
rect 12713 33473 12725 33507
rect 12759 33504 12771 33507
rect 12805 33507 12863 33513
rect 12805 33504 12817 33507
rect 12759 33476 12817 33504
rect 12759 33473 12771 33476
rect 12713 33467 12771 33473
rect 12805 33473 12817 33476
rect 12851 33473 12863 33507
rect 13372 33504 13400 33544
rect 13440 33541 13452 33575
rect 13486 33572 13498 33575
rect 14274 33572 14280 33584
rect 13486 33544 14280 33572
rect 13486 33541 13498 33544
rect 13440 33535 13498 33541
rect 14274 33532 14280 33544
rect 14332 33532 14338 33584
rect 14375 33572 14403 33612
rect 15194 33600 15200 33652
rect 15252 33640 15258 33652
rect 15381 33643 15439 33649
rect 15381 33640 15393 33643
rect 15252 33612 15393 33640
rect 15252 33600 15258 33612
rect 15381 33609 15393 33612
rect 15427 33609 15439 33643
rect 15746 33640 15752 33652
rect 15707 33612 15752 33640
rect 15381 33603 15439 33609
rect 15746 33600 15752 33612
rect 15804 33600 15810 33652
rect 18414 33640 18420 33652
rect 15856 33612 18420 33640
rect 15856 33572 15884 33612
rect 18414 33600 18420 33612
rect 18472 33600 18478 33652
rect 18506 33600 18512 33652
rect 18564 33640 18570 33652
rect 20073 33643 20131 33649
rect 18564 33612 20024 33640
rect 18564 33600 18570 33612
rect 19334 33572 19340 33584
rect 14375 33544 15884 33572
rect 16868 33544 19340 33572
rect 16868 33516 16896 33544
rect 13722 33504 13728 33516
rect 13372 33476 13728 33504
rect 12805 33467 12863 33473
rect 13722 33464 13728 33476
rect 13780 33464 13786 33516
rect 15841 33507 15899 33513
rect 15841 33473 15853 33507
rect 15887 33504 15899 33507
rect 16666 33504 16672 33516
rect 15887 33476 16672 33504
rect 15887 33473 15899 33476
rect 15841 33467 15899 33473
rect 16666 33464 16672 33476
rect 16724 33464 16730 33516
rect 16850 33504 16856 33516
rect 16811 33476 16856 33504
rect 16850 33464 16856 33476
rect 16908 33464 16914 33516
rect 17120 33507 17178 33513
rect 17120 33473 17132 33507
rect 17166 33504 17178 33507
rect 17862 33504 17868 33516
rect 17166 33476 17868 33504
rect 17166 33473 17178 33476
rect 17120 33467 17178 33473
rect 17862 33464 17868 33476
rect 17920 33464 17926 33516
rect 18708 33513 18736 33544
rect 19334 33532 19340 33544
rect 19392 33532 19398 33584
rect 19996 33572 20024 33612
rect 20073 33609 20085 33643
rect 20119 33640 20131 33643
rect 20162 33640 20168 33652
rect 20119 33612 20168 33640
rect 20119 33609 20131 33612
rect 20073 33603 20131 33609
rect 20162 33600 20168 33612
rect 20220 33600 20226 33652
rect 21910 33640 21916 33652
rect 21871 33612 21916 33640
rect 21910 33600 21916 33612
rect 21968 33600 21974 33652
rect 24581 33643 24639 33649
rect 24581 33609 24593 33643
rect 24627 33640 24639 33643
rect 24670 33640 24676 33652
rect 24627 33612 24676 33640
rect 24627 33609 24639 33612
rect 24581 33603 24639 33609
rect 24670 33600 24676 33612
rect 24728 33600 24734 33652
rect 25682 33600 25688 33652
rect 25740 33649 25746 33652
rect 25740 33643 25759 33649
rect 25747 33609 25759 33643
rect 25740 33603 25759 33609
rect 25740 33600 25746 33603
rect 29086 33600 29092 33652
rect 29144 33640 29150 33652
rect 29641 33643 29699 33649
rect 29641 33640 29653 33643
rect 29144 33612 29653 33640
rect 29144 33600 29150 33612
rect 29641 33609 29653 33612
rect 29687 33640 29699 33643
rect 30006 33640 30012 33652
rect 29687 33612 30012 33640
rect 29687 33609 29699 33612
rect 29641 33603 29699 33609
rect 30006 33600 30012 33612
rect 30064 33600 30070 33652
rect 30285 33643 30343 33649
rect 30285 33609 30297 33643
rect 30331 33640 30343 33643
rect 30834 33640 30840 33652
rect 30331 33612 30840 33640
rect 30331 33609 30343 33612
rect 30285 33603 30343 33609
rect 30834 33600 30840 33612
rect 30892 33600 30898 33652
rect 20717 33575 20775 33581
rect 19996 33544 20668 33572
rect 18693 33507 18751 33513
rect 18693 33473 18705 33507
rect 18739 33473 18751 33507
rect 18693 33467 18751 33473
rect 18782 33464 18788 33516
rect 18840 33504 18846 33516
rect 18949 33507 19007 33513
rect 18949 33504 18961 33507
rect 18840 33476 18961 33504
rect 18840 33464 18846 33476
rect 18949 33473 18961 33476
rect 18995 33473 19007 33507
rect 18949 33467 19007 33473
rect 20533 33507 20591 33513
rect 20533 33473 20545 33507
rect 20579 33473 20591 33507
rect 20640 33504 20668 33544
rect 20717 33541 20729 33575
rect 20763 33572 20775 33575
rect 21542 33572 21548 33584
rect 20763 33544 21548 33572
rect 20763 33541 20775 33544
rect 20717 33535 20775 33541
rect 21542 33532 21548 33544
rect 21600 33572 21606 33584
rect 22189 33575 22247 33581
rect 22189 33572 22201 33575
rect 21600 33544 22201 33572
rect 21600 33532 21606 33544
rect 22189 33541 22201 33544
rect 22235 33541 22247 33575
rect 22189 33535 22247 33541
rect 22922 33532 22928 33584
rect 22980 33572 22986 33584
rect 23707 33575 23765 33581
rect 23707 33572 23719 33575
rect 22980 33544 23719 33572
rect 22980 33532 22986 33544
rect 23707 33541 23719 33544
rect 23753 33572 23765 33575
rect 25498 33572 25504 33584
rect 23753 33544 24072 33572
rect 23753 33541 23765 33544
rect 23707 33535 23765 33541
rect 20809 33507 20867 33513
rect 20809 33504 20821 33507
rect 20640 33476 20821 33504
rect 20533 33467 20591 33473
rect 20809 33473 20821 33476
rect 20855 33473 20867 33507
rect 20809 33467 20867 33473
rect 13170 33436 13176 33448
rect 10008 33408 11008 33436
rect 13131 33408 13176 33436
rect 10008 33396 10014 33408
rect 13170 33396 13176 33408
rect 13228 33396 13234 33448
rect 15930 33436 15936 33448
rect 15891 33408 15936 33436
rect 15930 33396 15936 33408
rect 15988 33396 15994 33448
rect 20548 33436 20576 33467
rect 20622 33436 20628 33448
rect 20548 33408 20628 33436
rect 20622 33396 20628 33408
rect 20680 33396 20686 33448
rect 20824 33436 20852 33467
rect 21174 33464 21180 33516
rect 21232 33504 21238 33516
rect 21821 33507 21879 33513
rect 21821 33504 21833 33507
rect 21232 33476 21833 33504
rect 21232 33464 21238 33476
rect 21821 33473 21833 33476
rect 21867 33473 21879 33507
rect 22830 33504 22836 33516
rect 22791 33476 22836 33504
rect 21821 33467 21879 33473
rect 22830 33464 22836 33476
rect 22888 33464 22894 33516
rect 23293 33507 23351 33513
rect 23293 33473 23305 33507
rect 23339 33504 23351 33507
rect 23842 33504 23848 33516
rect 23339 33476 23848 33504
rect 23339 33473 23351 33476
rect 23293 33467 23351 33473
rect 23842 33464 23848 33476
rect 23900 33464 23906 33516
rect 22094 33436 22100 33448
rect 20824 33408 22100 33436
rect 22094 33396 22100 33408
rect 22152 33396 22158 33448
rect 22554 33396 22560 33448
rect 22612 33436 22618 33448
rect 24044 33436 24072 33544
rect 25056 33544 25504 33572
rect 24762 33504 24768 33516
rect 24723 33476 24768 33504
rect 24762 33464 24768 33476
rect 24820 33464 24826 33516
rect 25056 33513 25084 33544
rect 25498 33532 25504 33544
rect 25556 33532 25562 33584
rect 28994 33572 29000 33584
rect 28276 33544 29000 33572
rect 25041 33507 25099 33513
rect 25041 33473 25053 33507
rect 25087 33473 25099 33507
rect 27154 33504 27160 33516
rect 27115 33476 27160 33504
rect 25041 33467 25099 33473
rect 27154 33464 27160 33476
rect 27212 33464 27218 33516
rect 27433 33507 27491 33513
rect 27433 33473 27445 33507
rect 27479 33473 27491 33507
rect 27614 33504 27620 33516
rect 27575 33476 27620 33504
rect 27433 33467 27491 33473
rect 22612 33408 23612 33436
rect 24044 33408 25912 33436
rect 22612 33396 22618 33408
rect 6546 33368 6552 33380
rect 4764 33340 6552 33368
rect 4764 33328 4770 33340
rect 6546 33328 6552 33340
rect 6604 33328 6610 33380
rect 10226 33328 10232 33380
rect 10284 33368 10290 33380
rect 11517 33371 11575 33377
rect 11517 33368 11529 33371
rect 10284 33340 11529 33368
rect 10284 33328 10290 33340
rect 11517 33337 11529 33340
rect 11563 33337 11575 33371
rect 11517 33331 11575 33337
rect 20533 33371 20591 33377
rect 20533 33337 20545 33371
rect 20579 33368 20591 33371
rect 21358 33368 21364 33380
rect 20579 33340 21364 33368
rect 20579 33337 20591 33340
rect 20533 33331 20591 33337
rect 21358 33328 21364 33340
rect 21416 33328 21422 33380
rect 21542 33328 21548 33380
rect 21600 33368 21606 33380
rect 23474 33368 23480 33380
rect 21600 33340 23480 33368
rect 21600 33328 21606 33340
rect 23474 33328 23480 33340
rect 23532 33328 23538 33380
rect 23584 33368 23612 33408
rect 24118 33368 24124 33380
rect 23584 33340 24124 33368
rect 24118 33328 24124 33340
rect 24176 33328 24182 33380
rect 25884 33377 25912 33408
rect 27062 33396 27068 33448
rect 27120 33436 27126 33448
rect 27448 33436 27476 33467
rect 27614 33464 27620 33476
rect 27672 33464 27678 33516
rect 28276 33513 28304 33544
rect 28994 33532 29000 33544
rect 29052 33572 29058 33584
rect 29270 33572 29276 33584
rect 29052 33544 29276 33572
rect 29052 33532 29058 33544
rect 29270 33532 29276 33544
rect 29328 33532 29334 33584
rect 30098 33532 30104 33584
rect 30156 33572 30162 33584
rect 32232 33572 32260 33680
rect 32320 33572 33120 33586
rect 30156 33544 30788 33572
rect 32232 33544 33120 33572
rect 30156 33532 30162 33544
rect 28534 33513 28540 33516
rect 28261 33507 28319 33513
rect 28261 33473 28273 33507
rect 28307 33473 28319 33507
rect 28261 33467 28319 33473
rect 28528 33467 28540 33513
rect 28592 33504 28598 33516
rect 28592 33476 28628 33504
rect 28534 33464 28540 33467
rect 28592 33464 28598 33476
rect 29730 33464 29736 33516
rect 29788 33504 29794 33516
rect 30760 33513 30788 33544
rect 32320 33530 33120 33544
rect 30469 33507 30527 33513
rect 30469 33504 30481 33507
rect 29788 33476 30481 33504
rect 29788 33464 29794 33476
rect 30469 33473 30481 33476
rect 30515 33473 30527 33507
rect 30469 33467 30527 33473
rect 30745 33507 30803 33513
rect 30745 33473 30757 33507
rect 30791 33473 30803 33507
rect 30745 33467 30803 33473
rect 30929 33507 30987 33513
rect 30929 33473 30941 33507
rect 30975 33473 30987 33507
rect 30929 33467 30987 33473
rect 27120 33408 27476 33436
rect 27120 33396 27126 33408
rect 29454 33396 29460 33448
rect 29512 33436 29518 33448
rect 30944 33436 30972 33467
rect 31294 33436 31300 33448
rect 29512 33408 31300 33436
rect 29512 33396 29518 33408
rect 31294 33396 31300 33408
rect 31352 33396 31358 33448
rect 24949 33371 25007 33377
rect 24949 33337 24961 33371
rect 24995 33368 25007 33371
rect 25869 33371 25927 33377
rect 24995 33340 25820 33368
rect 24995 33337 25007 33340
rect 24949 33331 25007 33337
rect 2777 33303 2835 33309
rect 2777 33269 2789 33303
rect 2823 33300 2835 33303
rect 2866 33300 2872 33312
rect 2823 33272 2872 33300
rect 2823 33269 2835 33272
rect 2777 33263 2835 33269
rect 2866 33260 2872 33272
rect 2924 33260 2930 33312
rect 4614 33300 4620 33312
rect 4575 33272 4620 33300
rect 4614 33260 4620 33272
rect 4672 33260 4678 33312
rect 6641 33303 6699 33309
rect 6641 33269 6653 33303
rect 6687 33300 6699 33303
rect 7742 33300 7748 33312
rect 6687 33272 7748 33300
rect 6687 33269 6699 33272
rect 6641 33263 6699 33269
rect 7742 33260 7748 33272
rect 7800 33260 7806 33312
rect 10134 33300 10140 33312
rect 10095 33272 10140 33300
rect 10134 33260 10140 33272
rect 10192 33260 10198 33312
rect 10778 33300 10784 33312
rect 10739 33272 10784 33300
rect 10778 33260 10784 33272
rect 10836 33260 10842 33312
rect 12526 33300 12532 33312
rect 12487 33272 12532 33300
rect 12526 33260 12532 33272
rect 12584 33260 12590 33312
rect 14550 33300 14556 33312
rect 14511 33272 14556 33300
rect 14550 33260 14556 33272
rect 14608 33260 14614 33312
rect 18230 33300 18236 33312
rect 18191 33272 18236 33300
rect 18230 33260 18236 33272
rect 18288 33260 18294 33312
rect 20162 33260 20168 33312
rect 20220 33300 20226 33312
rect 20714 33300 20720 33312
rect 20220 33272 20720 33300
rect 20220 33260 20226 33272
rect 20714 33260 20720 33272
rect 20772 33260 20778 33312
rect 22002 33300 22008 33312
rect 21963 33272 22008 33300
rect 22002 33260 22008 33272
rect 22060 33260 22066 33312
rect 22097 33303 22155 33309
rect 22097 33269 22109 33303
rect 22143 33300 22155 33303
rect 22278 33300 22284 33312
rect 22143 33272 22284 33300
rect 22143 33269 22155 33272
rect 22097 33263 22155 33269
rect 22278 33260 22284 33272
rect 22336 33260 22342 33312
rect 22649 33303 22707 33309
rect 22649 33269 22661 33303
rect 22695 33300 22707 33303
rect 23290 33300 23296 33312
rect 22695 33272 23296 33300
rect 22695 33269 22707 33272
rect 22649 33263 22707 33269
rect 23290 33260 23296 33272
rect 23348 33260 23354 33312
rect 23658 33300 23664 33312
rect 23619 33272 23664 33300
rect 23658 33260 23664 33272
rect 23716 33260 23722 33312
rect 23842 33300 23848 33312
rect 23803 33272 23848 33300
rect 23842 33260 23848 33272
rect 23900 33260 23906 33312
rect 25130 33260 25136 33312
rect 25188 33300 25194 33312
rect 25685 33303 25743 33309
rect 25685 33300 25697 33303
rect 25188 33272 25697 33300
rect 25188 33260 25194 33272
rect 25685 33269 25697 33272
rect 25731 33269 25743 33303
rect 25792 33300 25820 33340
rect 25869 33337 25881 33371
rect 25915 33337 25927 33371
rect 25869 33331 25927 33337
rect 26142 33300 26148 33312
rect 25792 33272 26148 33300
rect 25685 33263 25743 33269
rect 26142 33260 26148 33272
rect 26200 33260 26206 33312
rect 26973 33303 27031 33309
rect 26973 33269 26985 33303
rect 27019 33300 27031 33303
rect 28166 33300 28172 33312
rect 27019 33272 28172 33300
rect 27019 33269 27031 33272
rect 26973 33263 27031 33269
rect 28166 33260 28172 33272
rect 28224 33260 28230 33312
rect 1104 33210 32016 33232
rect 1104 33158 2136 33210
rect 2188 33158 12440 33210
rect 12492 33158 22744 33210
rect 22796 33158 32016 33210
rect 1104 33136 32016 33158
rect 1670 33096 1676 33108
rect 1631 33068 1676 33096
rect 1670 33056 1676 33068
rect 1728 33056 1734 33108
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 3234 33096 3240 33108
rect 2924 33068 3240 33096
rect 2924 33056 2930 33068
rect 3234 33056 3240 33068
rect 3292 33096 3298 33108
rect 3329 33099 3387 33105
rect 3329 33096 3341 33099
rect 3292 33068 3341 33096
rect 3292 33056 3298 33068
rect 3329 33065 3341 33068
rect 3375 33096 3387 33099
rect 9125 33099 9183 33105
rect 3375 33068 7880 33096
rect 3375 33065 3387 33068
rect 3329 33059 3387 33065
rect 2041 33031 2099 33037
rect 2041 32997 2053 33031
rect 2087 33028 2099 33031
rect 2774 33028 2780 33040
rect 2087 33000 2780 33028
rect 2087 32997 2099 33000
rect 2041 32991 2099 32997
rect 2774 32988 2780 33000
rect 2832 32988 2838 33040
rect 3789 33031 3847 33037
rect 3789 32997 3801 33031
rect 3835 33028 3847 33031
rect 4154 33028 4160 33040
rect 3835 33000 4160 33028
rect 3835 32997 3847 33000
rect 3789 32991 3847 32997
rect 3418 32960 3424 32972
rect 2792 32932 3424 32960
rect 1857 32895 1915 32901
rect 1857 32861 1869 32895
rect 1903 32861 1915 32895
rect 1857 32855 1915 32861
rect 2133 32895 2191 32901
rect 2133 32861 2145 32895
rect 2179 32892 2191 32895
rect 2498 32892 2504 32904
rect 2179 32864 2504 32892
rect 2179 32861 2191 32864
rect 2133 32855 2191 32861
rect 1872 32824 1900 32855
rect 2498 32852 2504 32864
rect 2556 32852 2562 32904
rect 2792 32901 2820 32932
rect 3418 32920 3424 32932
rect 3476 32960 3482 32972
rect 3804 32960 3832 32991
rect 4154 32988 4160 33000
rect 4212 33028 4218 33040
rect 5350 33028 5356 33040
rect 4212 33000 5356 33028
rect 4212 32988 4218 33000
rect 5350 32988 5356 33000
rect 5408 32988 5414 33040
rect 5537 33031 5595 33037
rect 5537 32997 5549 33031
rect 5583 33028 5595 33031
rect 7558 33028 7564 33040
rect 5583 33000 7564 33028
rect 5583 32997 5595 33000
rect 5537 32991 5595 32997
rect 7558 32988 7564 33000
rect 7616 32988 7622 33040
rect 3476 32932 3832 32960
rect 3476 32920 3482 32932
rect 4614 32920 4620 32972
rect 4672 32960 4678 32972
rect 5442 32960 5448 32972
rect 4672 32932 5448 32960
rect 4672 32920 4678 32932
rect 5442 32920 5448 32932
rect 5500 32960 5506 32972
rect 6181 32963 6239 32969
rect 6181 32960 6193 32963
rect 5500 32932 6193 32960
rect 5500 32920 5506 32932
rect 6181 32929 6193 32932
rect 6227 32929 6239 32963
rect 7852 32960 7880 33068
rect 9125 33065 9137 33099
rect 9171 33096 9183 33099
rect 11606 33096 11612 33108
rect 9171 33068 11612 33096
rect 9171 33065 9183 33068
rect 9125 33059 9183 33065
rect 11606 33056 11612 33068
rect 11664 33056 11670 33108
rect 13449 33099 13507 33105
rect 13449 33096 13461 33099
rect 12406 33068 13461 33096
rect 8294 32988 8300 33040
rect 8352 33028 8358 33040
rect 10321 33031 10379 33037
rect 10321 33028 10333 33031
rect 8352 33000 10333 33028
rect 8352 32988 8358 33000
rect 10321 32997 10333 33000
rect 10367 32997 10379 33031
rect 10321 32991 10379 32997
rect 10410 32960 10416 32972
rect 7852 32932 8340 32960
rect 10371 32932 10416 32960
rect 6181 32923 6239 32929
rect 2777 32895 2835 32901
rect 2777 32861 2789 32895
rect 2823 32861 2835 32895
rect 3050 32892 3056 32904
rect 3011 32864 3056 32892
rect 2777 32855 2835 32861
rect 3050 32852 3056 32864
rect 3108 32852 3114 32904
rect 3237 32895 3295 32901
rect 3237 32861 3249 32895
rect 3283 32892 3295 32895
rect 3329 32895 3387 32901
rect 3329 32892 3341 32895
rect 3283 32864 3341 32892
rect 3283 32861 3295 32864
rect 3237 32855 3295 32861
rect 3329 32861 3341 32864
rect 3375 32861 3387 32895
rect 3970 32892 3976 32904
rect 3931 32864 3976 32892
rect 3329 32855 3387 32861
rect 3970 32852 3976 32864
rect 4028 32852 4034 32904
rect 4433 32895 4491 32901
rect 4433 32861 4445 32895
rect 4479 32861 4491 32895
rect 4433 32855 4491 32861
rect 2593 32827 2651 32833
rect 2593 32824 2605 32827
rect 1872 32796 2605 32824
rect 2593 32793 2605 32796
rect 2639 32793 2651 32827
rect 4448 32824 4476 32855
rect 4522 32852 4528 32904
rect 4580 32892 4586 32904
rect 4706 32892 4712 32904
rect 4580 32864 4712 32892
rect 4580 32852 4586 32864
rect 4706 32852 4712 32864
rect 4764 32852 4770 32904
rect 5902 32892 5908 32904
rect 5863 32864 5908 32892
rect 5902 32852 5908 32864
rect 5960 32852 5966 32904
rect 6086 32892 6092 32904
rect 6047 32864 6092 32892
rect 6086 32852 6092 32864
rect 6144 32852 6150 32904
rect 6733 32895 6791 32901
rect 6733 32861 6745 32895
rect 6779 32892 6791 32895
rect 6822 32892 6828 32904
rect 6779 32864 6828 32892
rect 6779 32861 6791 32864
rect 6733 32855 6791 32861
rect 6822 32852 6828 32864
rect 6880 32852 6886 32904
rect 7006 32892 7012 32904
rect 6967 32864 7012 32892
rect 7006 32852 7012 32864
rect 7064 32852 7070 32904
rect 7098 32852 7104 32904
rect 7156 32892 7162 32904
rect 7929 32895 7987 32901
rect 7156 32864 7201 32892
rect 7156 32852 7162 32864
rect 7929 32861 7941 32895
rect 7975 32892 7987 32895
rect 8110 32892 8116 32904
rect 7975 32864 8116 32892
rect 7975 32861 7987 32864
rect 7929 32855 7987 32861
rect 8110 32852 8116 32864
rect 8168 32852 8174 32904
rect 8205 32895 8263 32901
rect 8205 32861 8217 32895
rect 8251 32861 8263 32895
rect 8205 32855 8263 32861
rect 5445 32827 5503 32833
rect 5445 32824 5457 32827
rect 4448 32796 5457 32824
rect 2593 32787 2651 32793
rect 5445 32793 5457 32796
rect 5491 32793 5503 32827
rect 5810 32824 5816 32836
rect 5445 32787 5503 32793
rect 5552 32796 5816 32824
rect 3970 32716 3976 32768
rect 4028 32756 4034 32768
rect 5552 32756 5580 32796
rect 5810 32784 5816 32796
rect 5868 32784 5874 32836
rect 6362 32784 6368 32836
rect 6420 32824 6426 32836
rect 6917 32827 6975 32833
rect 6917 32824 6929 32827
rect 6420 32796 6929 32824
rect 6420 32784 6426 32796
rect 6917 32793 6929 32796
rect 6963 32793 6975 32827
rect 7116 32824 7144 32852
rect 8220 32824 8248 32855
rect 7116 32796 8248 32824
rect 6917 32787 6975 32793
rect 5718 32756 5724 32768
rect 4028 32728 5580 32756
rect 5679 32728 5724 32756
rect 4028 32716 4034 32728
rect 5718 32716 5724 32728
rect 5776 32716 5782 32768
rect 7285 32759 7343 32765
rect 7285 32725 7297 32759
rect 7331 32756 7343 32759
rect 7650 32756 7656 32768
rect 7331 32728 7656 32756
rect 7331 32725 7343 32728
rect 7285 32719 7343 32725
rect 7650 32716 7656 32728
rect 7708 32716 7714 32768
rect 7745 32759 7803 32765
rect 7745 32725 7757 32759
rect 7791 32756 7803 32759
rect 8018 32756 8024 32768
rect 7791 32728 8024 32756
rect 7791 32725 7803 32728
rect 7745 32719 7803 32725
rect 8018 32716 8024 32728
rect 8076 32716 8082 32768
rect 8113 32759 8171 32765
rect 8113 32725 8125 32759
rect 8159 32756 8171 32759
rect 8312 32756 8340 32932
rect 10410 32920 10416 32932
rect 10468 32920 10474 32972
rect 11882 32920 11888 32972
rect 11940 32960 11946 32972
rect 12406 32960 12434 33068
rect 13449 33065 13461 33068
rect 13495 33065 13507 33099
rect 13449 33059 13507 33065
rect 14461 33099 14519 33105
rect 14461 33065 14473 33099
rect 14507 33096 14519 33099
rect 14918 33096 14924 33108
rect 14507 33068 14924 33096
rect 14507 33065 14519 33068
rect 14461 33059 14519 33065
rect 14918 33056 14924 33068
rect 14976 33056 14982 33108
rect 16022 33056 16028 33108
rect 16080 33096 16086 33108
rect 16485 33099 16543 33105
rect 16485 33096 16497 33099
rect 16080 33068 16497 33096
rect 16080 33056 16086 33068
rect 16485 33065 16497 33068
rect 16531 33065 16543 33099
rect 16485 33059 16543 33065
rect 17405 33099 17463 33105
rect 17405 33065 17417 33099
rect 17451 33096 17463 33099
rect 22830 33096 22836 33108
rect 17451 33068 22692 33096
rect 22791 33068 22836 33096
rect 17451 33065 17463 33068
rect 17405 33059 17463 33065
rect 17034 32988 17040 33040
rect 17092 33028 17098 33040
rect 18601 33031 18659 33037
rect 18601 33028 18613 33031
rect 17092 33000 18613 33028
rect 17092 32988 17098 33000
rect 18601 32997 18613 33000
rect 18647 32997 18659 33031
rect 18601 32991 18659 32997
rect 21726 32988 21732 33040
rect 21784 33028 21790 33040
rect 22005 33031 22063 33037
rect 22005 33028 22017 33031
rect 21784 33000 22017 33028
rect 21784 32988 21790 33000
rect 22005 32997 22017 33000
rect 22051 32997 22063 33031
rect 22664 33028 22692 33068
rect 22830 33056 22836 33068
rect 22888 33056 22894 33108
rect 23201 33099 23259 33105
rect 23201 33065 23213 33099
rect 23247 33096 23259 33099
rect 25406 33096 25412 33108
rect 23247 33068 25412 33096
rect 23247 33065 23259 33068
rect 23201 33059 23259 33065
rect 25406 33056 25412 33068
rect 25464 33056 25470 33108
rect 25685 33099 25743 33105
rect 25685 33065 25697 33099
rect 25731 33096 25743 33099
rect 25774 33096 25780 33108
rect 25731 33068 25780 33096
rect 25731 33065 25743 33068
rect 25685 33059 25743 33065
rect 25774 33056 25780 33068
rect 25832 33056 25838 33108
rect 28537 33099 28595 33105
rect 28537 33065 28549 33099
rect 28583 33096 28595 33099
rect 28626 33096 28632 33108
rect 28583 33068 28632 33096
rect 28583 33065 28595 33068
rect 28537 33059 28595 33065
rect 28626 33056 28632 33068
rect 28684 33056 28690 33108
rect 29086 33096 29092 33108
rect 28736 33068 29092 33096
rect 24394 33028 24400 33040
rect 22664 33000 24400 33028
rect 22005 32991 22063 32997
rect 24394 32988 24400 33000
rect 24452 32988 24458 33040
rect 27614 33028 27620 33040
rect 25240 33000 27620 33028
rect 11940 32932 12434 32960
rect 11940 32920 11946 32932
rect 13170 32920 13176 32972
rect 13228 32960 13234 32972
rect 15105 32963 15163 32969
rect 15105 32960 15117 32963
rect 13228 32932 15117 32960
rect 13228 32920 13234 32932
rect 15105 32929 15117 32932
rect 15151 32929 15163 32963
rect 15105 32923 15163 32929
rect 16132 32932 18736 32960
rect 10137 32895 10195 32901
rect 10137 32861 10149 32895
rect 10183 32892 10195 32895
rect 10226 32892 10232 32904
rect 10183 32864 10232 32892
rect 10183 32861 10195 32864
rect 10137 32855 10195 32861
rect 10226 32852 10232 32864
rect 10284 32852 10290 32904
rect 10873 32895 10931 32901
rect 10873 32861 10885 32895
rect 10919 32892 10931 32895
rect 12618 32892 12624 32904
rect 10919 32864 12624 32892
rect 10919 32861 10931 32864
rect 10873 32855 10931 32861
rect 12618 32852 12624 32864
rect 12676 32852 12682 32904
rect 12713 32895 12771 32901
rect 12713 32861 12725 32895
rect 12759 32892 12771 32895
rect 13078 32892 13084 32904
rect 12759 32864 13084 32892
rect 12759 32861 12771 32864
rect 12713 32855 12771 32861
rect 13078 32852 13084 32864
rect 13136 32852 13142 32904
rect 13357 32895 13415 32901
rect 13357 32861 13369 32895
rect 13403 32861 13415 32895
rect 13357 32855 13415 32861
rect 8938 32824 8944 32836
rect 8899 32796 8944 32824
rect 8938 32784 8944 32796
rect 8996 32784 9002 32836
rect 9157 32827 9215 32833
rect 9157 32793 9169 32827
rect 9203 32824 9215 32827
rect 9858 32824 9864 32836
rect 9203 32796 9864 32824
rect 9203 32793 9215 32796
rect 9157 32787 9215 32793
rect 9858 32784 9864 32796
rect 9916 32784 9922 32836
rect 9953 32827 10011 32833
rect 9953 32793 9965 32827
rect 9999 32824 10011 32827
rect 11118 32827 11176 32833
rect 11118 32824 11130 32827
rect 9999 32796 11130 32824
rect 9999 32793 10011 32796
rect 9953 32787 10011 32793
rect 11118 32793 11130 32796
rect 11164 32793 11176 32827
rect 11118 32787 11176 32793
rect 11698 32784 11704 32836
rect 11756 32824 11762 32836
rect 11882 32824 11888 32836
rect 11756 32796 11888 32824
rect 11756 32784 11762 32796
rect 11882 32784 11888 32796
rect 11940 32784 11946 32836
rect 13372 32824 13400 32855
rect 14182 32852 14188 32904
rect 14240 32892 14246 32904
rect 14277 32895 14335 32901
rect 14277 32892 14289 32895
rect 14240 32864 14289 32892
rect 14240 32852 14246 32864
rect 14277 32861 14289 32864
rect 14323 32861 14335 32895
rect 14277 32855 14335 32861
rect 14550 32852 14556 32904
rect 14608 32892 14614 32904
rect 14918 32892 14924 32904
rect 14608 32864 14924 32892
rect 14608 32852 14614 32864
rect 14918 32852 14924 32864
rect 14976 32852 14982 32904
rect 15378 32901 15384 32904
rect 15372 32892 15384 32901
rect 15339 32864 15384 32892
rect 15372 32855 15384 32864
rect 15378 32852 15384 32855
rect 15436 32852 15442 32904
rect 15746 32852 15752 32904
rect 15804 32892 15810 32904
rect 16132 32892 16160 32932
rect 15804 32864 16160 32892
rect 15804 32852 15810 32864
rect 16206 32852 16212 32904
rect 16264 32892 16270 32904
rect 18708 32901 18736 32932
rect 18782 32920 18788 32972
rect 18840 32960 18846 32972
rect 20346 32960 20352 32972
rect 18840 32932 20352 32960
rect 18840 32920 18846 32932
rect 20346 32920 20352 32932
rect 20404 32920 20410 32972
rect 20530 32920 20536 32972
rect 20588 32960 20594 32972
rect 20625 32963 20683 32969
rect 20625 32960 20637 32963
rect 20588 32932 20637 32960
rect 20588 32920 20594 32932
rect 20625 32929 20637 32932
rect 20671 32929 20683 32963
rect 20625 32923 20683 32929
rect 21818 32920 21824 32972
rect 21876 32920 21882 32972
rect 22465 32963 22523 32969
rect 22465 32929 22477 32963
rect 22511 32960 22523 32963
rect 23198 32960 23204 32972
rect 22511 32932 23204 32960
rect 22511 32929 22523 32932
rect 22465 32923 22523 32929
rect 23198 32920 23204 32932
rect 23256 32920 23262 32972
rect 23566 32960 23572 32972
rect 23527 32932 23572 32960
rect 23566 32920 23572 32932
rect 23624 32920 23630 32972
rect 23658 32920 23664 32972
rect 23716 32960 23722 32972
rect 25240 32969 25268 33000
rect 27614 32988 27620 33000
rect 27672 32988 27678 33040
rect 25225 32963 25283 32969
rect 23716 32932 23761 32960
rect 23716 32920 23722 32932
rect 25225 32929 25237 32963
rect 25271 32929 25283 32963
rect 26605 32963 26663 32969
rect 26605 32960 26617 32963
rect 25225 32923 25283 32929
rect 25884 32932 26617 32960
rect 18509 32895 18567 32901
rect 18509 32892 18521 32895
rect 16264 32864 18521 32892
rect 16264 32852 16270 32864
rect 18509 32861 18521 32864
rect 18555 32861 18567 32895
rect 18509 32855 18567 32861
rect 18693 32895 18751 32901
rect 18693 32861 18705 32895
rect 18739 32861 18751 32895
rect 18693 32855 18751 32861
rect 19337 32895 19395 32901
rect 19337 32861 19349 32895
rect 19383 32861 19395 32895
rect 19337 32855 19395 32861
rect 12406 32796 14228 32824
rect 9306 32756 9312 32768
rect 8159 32728 8340 32756
rect 9267 32728 9312 32756
rect 8159 32725 8171 32728
rect 8113 32719 8171 32725
rect 9306 32716 9312 32728
rect 9364 32716 9370 32768
rect 12250 32756 12256 32768
rect 12211 32728 12256 32756
rect 12250 32716 12256 32728
rect 12308 32756 12314 32768
rect 12406 32756 12434 32796
rect 12308 32728 12434 32756
rect 12805 32759 12863 32765
rect 12308 32716 12314 32728
rect 12805 32725 12817 32759
rect 12851 32756 12863 32759
rect 13170 32756 13176 32768
rect 12851 32728 13176 32756
rect 12851 32725 12863 32728
rect 12805 32719 12863 32725
rect 13170 32716 13176 32728
rect 13228 32716 13234 32768
rect 14090 32756 14096 32768
rect 14051 32728 14096 32756
rect 14090 32716 14096 32728
rect 14148 32716 14154 32768
rect 14200 32756 14228 32796
rect 16114 32784 16120 32836
rect 16172 32824 16178 32836
rect 17681 32827 17739 32833
rect 17681 32824 17693 32827
rect 16172 32796 17693 32824
rect 16172 32784 16178 32796
rect 17681 32793 17693 32796
rect 17727 32793 17739 32827
rect 17681 32787 17739 32793
rect 17957 32827 18015 32833
rect 17957 32793 17969 32827
rect 18003 32824 18015 32827
rect 18230 32824 18236 32836
rect 18003 32796 18236 32824
rect 18003 32793 18015 32796
rect 17957 32787 18015 32793
rect 18230 32784 18236 32796
rect 18288 32784 18294 32836
rect 19352 32824 19380 32855
rect 19610 32852 19616 32904
rect 19668 32892 19674 32904
rect 19981 32895 20039 32901
rect 19981 32892 19993 32895
rect 19668 32864 19993 32892
rect 19668 32852 19674 32864
rect 19981 32861 19993 32864
rect 20027 32892 20039 32895
rect 21726 32892 21732 32904
rect 20027 32864 21732 32892
rect 20027 32861 20039 32864
rect 19981 32855 20039 32861
rect 21726 32852 21732 32864
rect 21784 32852 21790 32904
rect 20438 32824 20444 32836
rect 19352 32796 20444 32824
rect 20438 32784 20444 32796
rect 20496 32784 20502 32836
rect 20892 32827 20950 32833
rect 20892 32793 20904 32827
rect 20938 32824 20950 32827
rect 21836 32824 21864 32920
rect 22649 32895 22707 32901
rect 22649 32861 22661 32895
rect 22695 32892 22707 32895
rect 22922 32892 22928 32904
rect 22695 32864 22928 32892
rect 22695 32861 22707 32864
rect 22649 32855 22707 32861
rect 22922 32852 22928 32864
rect 22980 32852 22986 32904
rect 23477 32895 23535 32901
rect 23477 32861 23489 32895
rect 23523 32861 23535 32895
rect 23477 32855 23535 32861
rect 23753 32895 23811 32901
rect 23753 32861 23765 32895
rect 23799 32892 23811 32895
rect 23842 32892 23848 32904
rect 23799 32864 23848 32892
rect 23799 32861 23811 32864
rect 23753 32855 23811 32861
rect 20938 32796 21864 32824
rect 20938 32793 20950 32796
rect 20892 32787 20950 32793
rect 21910 32784 21916 32836
rect 21968 32824 21974 32836
rect 23201 32827 23259 32833
rect 23201 32824 23213 32827
rect 21968 32796 23213 32824
rect 21968 32784 21974 32796
rect 23201 32793 23213 32796
rect 23247 32793 23259 32827
rect 23492 32824 23520 32855
rect 23842 32852 23848 32864
rect 23900 32852 23906 32904
rect 24946 32892 24952 32904
rect 24907 32864 24952 32892
rect 24946 32852 24952 32864
rect 25004 32852 25010 32904
rect 25884 32901 25912 32932
rect 26605 32929 26617 32932
rect 26651 32929 26663 32963
rect 27154 32960 27160 32972
rect 26605 32923 26663 32929
rect 26804 32932 27160 32960
rect 25133 32895 25191 32901
rect 25133 32861 25145 32895
rect 25179 32861 25191 32895
rect 25133 32855 25191 32861
rect 25869 32895 25927 32901
rect 25869 32861 25881 32895
rect 25915 32861 25927 32895
rect 26050 32892 26056 32904
rect 26011 32864 26056 32892
rect 25869 32855 25927 32861
rect 23934 32824 23940 32836
rect 23492 32796 23940 32824
rect 23201 32787 23259 32793
rect 23934 32784 23940 32796
rect 23992 32784 23998 32836
rect 25148 32824 25176 32855
rect 26050 32852 26056 32864
rect 26108 32852 26114 32904
rect 26145 32895 26203 32901
rect 26145 32861 26157 32895
rect 26191 32861 26203 32895
rect 26145 32855 26203 32861
rect 26068 32824 26096 32852
rect 25148 32796 26096 32824
rect 16390 32756 16396 32768
rect 14200 32728 16396 32756
rect 16390 32716 16396 32728
rect 16448 32716 16454 32768
rect 17218 32716 17224 32768
rect 17276 32756 17282 32768
rect 17865 32759 17923 32765
rect 17865 32756 17877 32759
rect 17276 32728 17877 32756
rect 17276 32716 17282 32728
rect 17865 32725 17877 32728
rect 17911 32725 17923 32759
rect 17865 32719 17923 32725
rect 19429 32759 19487 32765
rect 19429 32725 19441 32759
rect 19475 32756 19487 32759
rect 19702 32756 19708 32768
rect 19475 32728 19708 32756
rect 19475 32725 19487 32728
rect 19429 32719 19487 32725
rect 19702 32716 19708 32728
rect 19760 32716 19766 32768
rect 20073 32759 20131 32765
rect 20073 32725 20085 32759
rect 20119 32756 20131 32759
rect 21174 32756 21180 32768
rect 20119 32728 21180 32756
rect 20119 32725 20131 32728
rect 20073 32719 20131 32725
rect 21174 32716 21180 32728
rect 21232 32756 21238 32768
rect 22830 32756 22836 32768
rect 21232 32728 22836 32756
rect 21232 32716 21238 32728
rect 22830 32716 22836 32728
rect 22888 32716 22894 32768
rect 23293 32759 23351 32765
rect 23293 32725 23305 32759
rect 23339 32756 23351 32759
rect 23382 32756 23388 32768
rect 23339 32728 23388 32756
rect 23339 32725 23351 32728
rect 23293 32719 23351 32725
rect 23382 32716 23388 32728
rect 23440 32716 23446 32768
rect 24670 32716 24676 32768
rect 24728 32756 24734 32768
rect 24765 32759 24823 32765
rect 24765 32756 24777 32759
rect 24728 32728 24777 32756
rect 24728 32716 24734 32728
rect 24765 32725 24777 32728
rect 24811 32725 24823 32759
rect 26160 32756 26188 32855
rect 26694 32852 26700 32904
rect 26752 32892 26758 32904
rect 26804 32901 26832 32932
rect 27154 32920 27160 32932
rect 27212 32920 27218 32972
rect 27522 32920 27528 32972
rect 27580 32960 27586 32972
rect 28736 32960 28764 33068
rect 29086 33056 29092 33068
rect 29144 33056 29150 33108
rect 31294 33096 31300 33108
rect 31255 33068 31300 33096
rect 31294 33056 31300 33068
rect 31352 33056 31358 33108
rect 28902 33028 28908 33040
rect 28863 33000 28908 33028
rect 28902 32988 28908 33000
rect 28960 32988 28966 33040
rect 27580 32932 28764 32960
rect 27580 32920 27586 32932
rect 29270 32920 29276 32972
rect 29328 32960 29334 32972
rect 29917 32963 29975 32969
rect 29917 32960 29929 32963
rect 29328 32932 29929 32960
rect 29328 32920 29334 32932
rect 29917 32929 29929 32932
rect 29963 32929 29975 32963
rect 29917 32923 29975 32929
rect 26789 32895 26847 32901
rect 26789 32892 26801 32895
rect 26752 32864 26801 32892
rect 26752 32852 26758 32864
rect 26789 32861 26801 32864
rect 26835 32861 26847 32895
rect 27062 32892 27068 32904
rect 27023 32864 27068 32892
rect 26789 32855 26847 32861
rect 27062 32852 27068 32864
rect 27120 32852 27126 32904
rect 27249 32895 27307 32901
rect 27249 32861 27261 32895
rect 27295 32892 27307 32895
rect 27798 32892 27804 32904
rect 27295 32864 27804 32892
rect 27295 32861 27307 32864
rect 27249 32855 27307 32861
rect 27798 32852 27804 32864
rect 27856 32892 27862 32904
rect 28258 32892 28264 32904
rect 27856 32864 28264 32892
rect 27856 32852 27862 32864
rect 28258 32852 28264 32864
rect 28316 32892 28322 32904
rect 28626 32892 28632 32904
rect 28316 32864 28632 32892
rect 28316 32852 28322 32864
rect 28626 32852 28632 32864
rect 28684 32852 28690 32904
rect 30190 32901 30196 32904
rect 28721 32895 28779 32901
rect 28721 32861 28733 32895
rect 28767 32861 28779 32895
rect 28721 32855 28779 32861
rect 28997 32895 29055 32901
rect 28997 32861 29009 32895
rect 29043 32892 29055 32895
rect 30184 32892 30196 32901
rect 29043 32864 29684 32892
rect 30151 32864 30196 32892
rect 29043 32861 29055 32864
rect 28997 32855 29055 32861
rect 26326 32784 26332 32836
rect 26384 32824 26390 32836
rect 27080 32824 27108 32852
rect 26384 32796 27108 32824
rect 27893 32827 27951 32833
rect 26384 32784 26390 32796
rect 27893 32793 27905 32827
rect 27939 32824 27951 32827
rect 28074 32824 28080 32836
rect 27939 32796 28080 32824
rect 27939 32793 27951 32796
rect 27893 32787 27951 32793
rect 28074 32784 28080 32796
rect 28132 32784 28138 32836
rect 28736 32824 28764 32855
rect 29546 32824 29552 32836
rect 28736 32796 29552 32824
rect 29546 32784 29552 32796
rect 29604 32784 29610 32836
rect 29656 32824 29684 32864
rect 30184 32855 30196 32864
rect 30190 32852 30196 32855
rect 30248 32852 30254 32904
rect 30466 32824 30472 32836
rect 29656 32796 30472 32824
rect 30466 32784 30472 32796
rect 30524 32824 30530 32836
rect 30926 32824 30932 32836
rect 30524 32796 30932 32824
rect 30524 32784 30530 32796
rect 30926 32784 30932 32796
rect 30984 32784 30990 32836
rect 27522 32756 27528 32768
rect 26160 32728 27528 32756
rect 24765 32719 24823 32725
rect 27522 32716 27528 32728
rect 27580 32716 27586 32768
rect 27985 32759 28043 32765
rect 27985 32725 27997 32759
rect 28031 32756 28043 32759
rect 28902 32756 28908 32768
rect 28031 32728 28908 32756
rect 28031 32725 28043 32728
rect 27985 32719 28043 32725
rect 28902 32716 28908 32728
rect 28960 32716 28966 32768
rect 29638 32716 29644 32768
rect 29696 32756 29702 32768
rect 31110 32756 31116 32768
rect 29696 32728 31116 32756
rect 29696 32716 29702 32728
rect 31110 32716 31116 32728
rect 31168 32716 31174 32768
rect 1104 32666 32016 32688
rect 1104 32614 7288 32666
rect 7340 32614 17592 32666
rect 17644 32614 27896 32666
rect 27948 32614 32016 32666
rect 1104 32592 32016 32614
rect 5626 32512 5632 32564
rect 5684 32552 5690 32564
rect 5813 32555 5871 32561
rect 5813 32552 5825 32555
rect 5684 32524 5825 32552
rect 5684 32512 5690 32524
rect 5813 32521 5825 32524
rect 5859 32521 5871 32555
rect 5813 32515 5871 32521
rect 5902 32512 5908 32564
rect 5960 32552 5966 32564
rect 6365 32555 6423 32561
rect 6365 32552 6377 32555
rect 5960 32524 6377 32552
rect 5960 32512 5966 32524
rect 6365 32521 6377 32524
rect 6411 32521 6423 32555
rect 6365 32515 6423 32521
rect 8665 32555 8723 32561
rect 8665 32521 8677 32555
rect 8711 32552 8723 32555
rect 9306 32552 9312 32564
rect 8711 32524 9312 32552
rect 8711 32521 8723 32524
rect 8665 32515 8723 32521
rect 9306 32512 9312 32524
rect 9364 32512 9370 32564
rect 11885 32555 11943 32561
rect 11885 32521 11897 32555
rect 11931 32552 11943 32555
rect 12250 32552 12256 32564
rect 11931 32524 12256 32552
rect 11931 32521 11943 32524
rect 11885 32515 11943 32521
rect 12250 32512 12256 32524
rect 12308 32512 12314 32564
rect 13354 32552 13360 32564
rect 12406 32524 13360 32552
rect 3050 32444 3056 32496
rect 3108 32484 3114 32496
rect 4246 32484 4252 32496
rect 3108 32456 4252 32484
rect 3108 32444 3114 32456
rect 1394 32416 1400 32428
rect 1355 32388 1400 32416
rect 1394 32376 1400 32388
rect 1452 32376 1458 32428
rect 1664 32419 1722 32425
rect 1664 32385 1676 32419
rect 1710 32416 1722 32419
rect 2406 32416 2412 32428
rect 1710 32388 2412 32416
rect 1710 32385 1722 32388
rect 1664 32379 1722 32385
rect 2406 32376 2412 32388
rect 2464 32376 2470 32428
rect 3418 32416 3424 32428
rect 3379 32388 3424 32416
rect 3418 32376 3424 32388
rect 3476 32376 3482 32428
rect 3712 32425 3740 32456
rect 4246 32444 4252 32456
rect 4304 32484 4310 32496
rect 4522 32484 4528 32496
rect 4304 32456 4528 32484
rect 4304 32444 4310 32456
rect 4522 32444 4528 32456
rect 4580 32444 4586 32496
rect 4700 32487 4758 32493
rect 4700 32453 4712 32487
rect 4746 32484 4758 32487
rect 5718 32484 5724 32496
rect 4746 32456 5724 32484
rect 4746 32453 4758 32456
rect 4700 32447 4758 32453
rect 5718 32444 5724 32456
rect 5776 32444 5782 32496
rect 7653 32487 7711 32493
rect 7653 32484 7665 32487
rect 5828 32456 7665 32484
rect 3697 32419 3755 32425
rect 3697 32385 3709 32419
rect 3743 32385 3755 32419
rect 3697 32379 3755 32385
rect 3881 32419 3939 32425
rect 3881 32385 3893 32419
rect 3927 32416 3939 32419
rect 4430 32416 4436 32428
rect 3927 32388 4016 32416
rect 4391 32388 4436 32416
rect 3927 32385 3939 32388
rect 3881 32379 3939 32385
rect 2498 32240 2504 32292
rect 2556 32280 2562 32292
rect 2777 32283 2835 32289
rect 2777 32280 2789 32283
rect 2556 32252 2789 32280
rect 2556 32240 2562 32252
rect 2777 32249 2789 32252
rect 2823 32280 2835 32283
rect 3988 32280 4016 32388
rect 4430 32376 4436 32388
rect 4488 32376 4494 32428
rect 4982 32376 4988 32428
rect 5040 32416 5046 32428
rect 5828 32416 5856 32456
rect 7653 32453 7665 32456
rect 7699 32453 7711 32487
rect 7834 32484 7840 32496
rect 7795 32456 7840 32484
rect 7653 32447 7711 32453
rect 7834 32444 7840 32456
rect 7892 32444 7898 32496
rect 8202 32444 8208 32496
rect 8260 32484 8266 32496
rect 8757 32487 8815 32493
rect 8757 32484 8769 32487
rect 8260 32456 8769 32484
rect 8260 32444 8266 32456
rect 8757 32453 8769 32456
rect 8803 32453 8815 32487
rect 11514 32484 11520 32496
rect 8757 32447 8815 32453
rect 9508 32456 11520 32484
rect 5040 32388 5856 32416
rect 6549 32419 6607 32425
rect 5040 32376 5046 32388
rect 6549 32385 6561 32419
rect 6595 32385 6607 32419
rect 6549 32379 6607 32385
rect 5442 32308 5448 32360
rect 5500 32348 5506 32360
rect 6564 32348 6592 32379
rect 6638 32376 6644 32428
rect 6696 32416 6702 32428
rect 6825 32419 6883 32425
rect 6825 32416 6837 32419
rect 6696 32388 6837 32416
rect 6696 32376 6702 32388
rect 6825 32385 6837 32388
rect 6871 32385 6883 32419
rect 7009 32419 7067 32425
rect 7009 32416 7021 32419
rect 6825 32379 6883 32385
rect 6932 32388 7021 32416
rect 5500 32320 6592 32348
rect 5500 32308 5506 32320
rect 6546 32280 6552 32292
rect 2823 32252 4016 32280
rect 2823 32249 2835 32252
rect 2777 32243 2835 32249
rect 2682 32172 2688 32224
rect 2740 32212 2746 32224
rect 3237 32215 3295 32221
rect 3237 32212 3249 32215
rect 2740 32184 3249 32212
rect 2740 32172 2746 32184
rect 3237 32181 3249 32184
rect 3283 32181 3295 32215
rect 3988 32212 4016 32252
rect 5368 32252 6552 32280
rect 5368 32212 5396 32252
rect 6546 32240 6552 32252
rect 6604 32240 6610 32292
rect 3988 32184 5396 32212
rect 3237 32175 3295 32181
rect 5626 32172 5632 32224
rect 5684 32212 5690 32224
rect 6638 32212 6644 32224
rect 5684 32184 6644 32212
rect 5684 32172 5690 32184
rect 6638 32172 6644 32184
rect 6696 32212 6702 32224
rect 6932 32212 6960 32388
rect 7009 32385 7021 32388
rect 7055 32385 7067 32419
rect 7009 32379 7067 32385
rect 8573 32419 8631 32425
rect 8573 32385 8585 32419
rect 8619 32416 8631 32419
rect 9214 32416 9220 32428
rect 8619 32388 9220 32416
rect 8619 32385 8631 32388
rect 8573 32379 8631 32385
rect 9214 32376 9220 32388
rect 9272 32376 9278 32428
rect 9508 32425 9536 32456
rect 11514 32444 11520 32456
rect 11572 32444 11578 32496
rect 11606 32444 11612 32496
rect 11664 32484 11670 32496
rect 12406 32484 12434 32524
rect 13354 32512 13360 32524
rect 13412 32552 13418 32564
rect 14458 32552 14464 32564
rect 13412 32524 14228 32552
rect 14419 32524 14464 32552
rect 13412 32512 13418 32524
rect 11664 32456 12434 32484
rect 12529 32487 12587 32493
rect 11664 32444 11670 32456
rect 12529 32453 12541 32487
rect 12575 32484 12587 32487
rect 12710 32484 12716 32496
rect 12575 32456 12716 32484
rect 12575 32453 12587 32456
rect 12529 32447 12587 32453
rect 12710 32444 12716 32456
rect 12768 32444 12774 32496
rect 12888 32487 12946 32493
rect 12888 32453 12900 32487
rect 12934 32484 12946 32487
rect 14090 32484 14096 32496
rect 12934 32456 14096 32484
rect 12934 32453 12946 32456
rect 12888 32447 12946 32453
rect 14090 32444 14096 32456
rect 14148 32444 14154 32496
rect 14200 32484 14228 32524
rect 14458 32512 14464 32524
rect 14516 32512 14522 32564
rect 15378 32552 15384 32564
rect 14568 32524 15384 32552
rect 14568 32484 14596 32524
rect 15378 32512 15384 32524
rect 15436 32512 15442 32564
rect 16114 32552 16120 32564
rect 16075 32524 16120 32552
rect 16114 32512 16120 32524
rect 16172 32512 16178 32564
rect 16666 32552 16672 32564
rect 16627 32524 16672 32552
rect 16666 32512 16672 32524
rect 16724 32512 16730 32564
rect 17862 32552 17868 32564
rect 17823 32524 17868 32552
rect 17862 32512 17868 32524
rect 17920 32512 17926 32564
rect 19334 32512 19340 32564
rect 19392 32552 19398 32564
rect 19392 32524 19647 32552
rect 19392 32512 19398 32524
rect 15194 32484 15200 32496
rect 14200 32456 14596 32484
rect 14936 32456 15200 32484
rect 9493 32419 9551 32425
rect 9493 32385 9505 32419
rect 9539 32385 9551 32419
rect 9749 32419 9807 32425
rect 9749 32416 9761 32419
rect 9493 32379 9551 32385
rect 9600 32388 9761 32416
rect 9033 32351 9091 32357
rect 9033 32317 9045 32351
rect 9079 32348 9091 32351
rect 9398 32348 9404 32360
rect 9079 32320 9404 32348
rect 9079 32317 9091 32320
rect 9033 32311 9091 32317
rect 9398 32308 9404 32320
rect 9456 32308 9462 32360
rect 9600 32348 9628 32388
rect 9749 32385 9761 32388
rect 9795 32385 9807 32419
rect 9749 32379 9807 32385
rect 12250 32376 12256 32428
rect 12308 32416 12314 32428
rect 14936 32425 14964 32456
rect 15194 32444 15200 32456
rect 15252 32484 15258 32496
rect 15654 32484 15660 32496
rect 15252 32456 15660 32484
rect 15252 32444 15258 32456
rect 15654 32444 15660 32456
rect 15712 32444 15718 32496
rect 19518 32484 19524 32496
rect 18340 32456 19524 32484
rect 14645 32419 14703 32425
rect 12308 32388 14044 32416
rect 12308 32376 12314 32388
rect 12618 32348 12624 32360
rect 9508 32320 9628 32348
rect 12579 32320 12624 32348
rect 8297 32283 8355 32289
rect 8297 32249 8309 32283
rect 8343 32280 8355 32283
rect 9508 32280 9536 32320
rect 12618 32308 12624 32320
rect 12676 32308 12682 32360
rect 8343 32252 9536 32280
rect 8343 32249 8355 32252
rect 8297 32243 8355 32249
rect 10502 32240 10508 32292
rect 10560 32280 10566 32292
rect 11517 32283 11575 32289
rect 11517 32280 11529 32283
rect 10560 32252 11529 32280
rect 10560 32240 10566 32252
rect 11517 32249 11529 32252
rect 11563 32249 11575 32283
rect 11517 32243 11575 32249
rect 8938 32212 8944 32224
rect 6696 32184 6960 32212
rect 8899 32184 8944 32212
rect 6696 32172 6702 32184
rect 8938 32172 8944 32184
rect 8996 32172 9002 32224
rect 10873 32215 10931 32221
rect 10873 32181 10885 32215
rect 10919 32212 10931 32215
rect 11885 32215 11943 32221
rect 11885 32212 11897 32215
rect 10919 32184 11897 32212
rect 10919 32181 10931 32184
rect 10873 32175 10931 32181
rect 11885 32181 11897 32184
rect 11931 32181 11943 32215
rect 12066 32212 12072 32224
rect 12027 32184 12072 32212
rect 11885 32175 11943 32181
rect 12066 32172 12072 32184
rect 12124 32212 12130 32224
rect 12529 32215 12587 32221
rect 12529 32212 12541 32215
rect 12124 32184 12541 32212
rect 12124 32172 12130 32184
rect 12529 32181 12541 32184
rect 12575 32181 12587 32215
rect 12636 32212 12664 32308
rect 14016 32289 14044 32388
rect 14645 32385 14657 32419
rect 14691 32385 14703 32419
rect 14645 32379 14703 32385
rect 14921 32419 14979 32425
rect 14921 32385 14933 32419
rect 14967 32385 14979 32419
rect 14921 32379 14979 32385
rect 14366 32308 14372 32360
rect 14424 32348 14430 32360
rect 14660 32348 14688 32379
rect 15010 32376 15016 32428
rect 15068 32416 15074 32428
rect 15105 32419 15163 32425
rect 15105 32416 15117 32419
rect 15068 32388 15117 32416
rect 15068 32376 15074 32388
rect 15105 32385 15117 32388
rect 15151 32385 15163 32419
rect 15105 32379 15163 32385
rect 15562 32376 15568 32428
rect 15620 32416 15626 32428
rect 15933 32419 15991 32425
rect 15933 32416 15945 32419
rect 15620 32388 15945 32416
rect 15620 32376 15626 32388
rect 15933 32385 15945 32388
rect 15979 32385 15991 32419
rect 17034 32416 17040 32428
rect 16995 32388 17040 32416
rect 15933 32379 15991 32385
rect 17034 32376 17040 32388
rect 17092 32376 17098 32428
rect 17144 32388 17632 32416
rect 17144 32360 17172 32388
rect 15286 32348 15292 32360
rect 14424 32320 15292 32348
rect 14424 32308 14430 32320
rect 15286 32308 15292 32320
rect 15344 32348 15350 32360
rect 15470 32348 15476 32360
rect 15344 32320 15476 32348
rect 15344 32308 15350 32320
rect 15470 32308 15476 32320
rect 15528 32308 15534 32360
rect 15749 32351 15807 32357
rect 15749 32317 15761 32351
rect 15795 32348 15807 32351
rect 16942 32348 16948 32360
rect 15795 32320 16948 32348
rect 15795 32317 15807 32320
rect 15749 32311 15807 32317
rect 16942 32308 16948 32320
rect 17000 32308 17006 32360
rect 17126 32348 17132 32360
rect 17087 32320 17132 32348
rect 17126 32308 17132 32320
rect 17184 32308 17190 32360
rect 17221 32351 17279 32357
rect 17221 32317 17233 32351
rect 17267 32317 17279 32351
rect 17604 32348 17632 32388
rect 17678 32376 17684 32428
rect 17736 32416 17742 32428
rect 18049 32419 18107 32425
rect 18049 32416 18061 32419
rect 17736 32388 18061 32416
rect 17736 32376 17742 32388
rect 18049 32385 18061 32388
rect 18095 32385 18107 32419
rect 18049 32379 18107 32385
rect 18138 32376 18144 32428
rect 18196 32416 18202 32428
rect 18340 32425 18368 32456
rect 19518 32444 19524 32456
rect 19576 32444 19582 32496
rect 19619 32484 19647 32524
rect 19978 32512 19984 32564
rect 20036 32552 20042 32564
rect 20441 32555 20499 32561
rect 20441 32552 20453 32555
rect 20036 32524 20453 32552
rect 20036 32512 20042 32524
rect 20441 32521 20453 32524
rect 20487 32552 20499 32555
rect 27706 32552 27712 32564
rect 20487 32524 27712 32552
rect 20487 32521 20499 32524
rect 20441 32515 20499 32521
rect 27706 32512 27712 32524
rect 27764 32512 27770 32564
rect 28074 32512 28080 32564
rect 28132 32552 28138 32564
rect 28350 32552 28356 32564
rect 28132 32524 28356 32552
rect 28132 32512 28138 32524
rect 28350 32512 28356 32524
rect 28408 32512 28414 32564
rect 28442 32512 28448 32564
rect 28500 32552 28506 32564
rect 31297 32555 31355 32561
rect 31297 32552 31309 32555
rect 28500 32524 31309 32552
rect 28500 32512 28506 32524
rect 31297 32521 31309 32524
rect 31343 32521 31355 32555
rect 31297 32515 31355 32521
rect 19619 32456 21119 32484
rect 18325 32419 18383 32425
rect 18325 32416 18337 32419
rect 18196 32388 18337 32416
rect 18196 32376 18202 32388
rect 18325 32385 18337 32388
rect 18371 32385 18383 32419
rect 18325 32379 18383 32385
rect 18966 32376 18972 32428
rect 19024 32416 19030 32428
rect 19337 32419 19395 32425
rect 19337 32416 19349 32419
rect 19024 32388 19349 32416
rect 19024 32376 19030 32388
rect 19337 32385 19349 32388
rect 19383 32385 19395 32419
rect 19610 32416 19616 32428
rect 19571 32388 19616 32416
rect 19337 32379 19395 32385
rect 19610 32376 19616 32388
rect 19668 32376 19674 32428
rect 20346 32416 20352 32428
rect 20307 32388 20352 32416
rect 20346 32376 20352 32388
rect 20404 32376 20410 32428
rect 20993 32419 21051 32425
rect 20993 32385 21005 32419
rect 21039 32385 21051 32419
rect 21091 32416 21119 32456
rect 21174 32444 21180 32496
rect 21232 32484 21238 32496
rect 22005 32487 22063 32493
rect 21232 32456 21277 32484
rect 21376 32456 21947 32484
rect 21232 32444 21238 32456
rect 21269 32419 21327 32425
rect 21269 32416 21281 32419
rect 21091 32388 21281 32416
rect 20993 32379 21051 32385
rect 21269 32385 21281 32388
rect 21315 32416 21327 32419
rect 21376 32416 21404 32456
rect 21315 32388 21404 32416
rect 21637 32419 21695 32425
rect 21315 32385 21327 32388
rect 21269 32379 21327 32385
rect 21637 32385 21649 32419
rect 21683 32416 21695 32419
rect 21821 32419 21879 32425
rect 21821 32416 21833 32419
rect 21683 32388 21833 32416
rect 21683 32385 21695 32388
rect 21637 32379 21695 32385
rect 21821 32385 21833 32388
rect 21867 32385 21879 32419
rect 21919 32416 21947 32456
rect 22005 32453 22017 32487
rect 22051 32484 22063 32487
rect 22824 32487 22882 32493
rect 22051 32456 22775 32484
rect 22051 32453 22063 32456
rect 22005 32447 22063 32453
rect 21919 32388 22048 32416
rect 21821 32379 21879 32385
rect 20162 32348 20168 32360
rect 17604 32320 20168 32348
rect 17221 32311 17279 32317
rect 14001 32283 14059 32289
rect 14001 32249 14013 32283
rect 14047 32280 14059 32283
rect 14826 32280 14832 32292
rect 14047 32252 14832 32280
rect 14047 32249 14059 32252
rect 14001 32243 14059 32249
rect 14826 32240 14832 32252
rect 14884 32240 14890 32292
rect 16298 32240 16304 32292
rect 16356 32280 16362 32292
rect 17236 32280 17264 32311
rect 20162 32308 20168 32320
rect 20220 32308 20226 32360
rect 20622 32308 20628 32360
rect 20680 32348 20686 32360
rect 21008 32348 21036 32379
rect 21174 32348 21180 32360
rect 20680 32320 20946 32348
rect 21008 32320 21180 32348
rect 20680 32308 20686 32320
rect 16356 32252 17264 32280
rect 16356 32240 16362 32252
rect 17770 32240 17776 32292
rect 17828 32280 17834 32292
rect 18233 32283 18291 32289
rect 18233 32280 18245 32283
rect 17828 32252 18245 32280
rect 17828 32240 17834 32252
rect 18233 32249 18245 32252
rect 18279 32280 18291 32283
rect 19521 32283 19579 32289
rect 19521 32280 19533 32283
rect 18279 32252 19533 32280
rect 18279 32249 18291 32252
rect 18233 32243 18291 32249
rect 19521 32249 19533 32252
rect 19567 32249 19579 32283
rect 20918 32280 20946 32320
rect 21174 32308 21180 32320
rect 21232 32308 21238 32360
rect 21358 32308 21364 32360
rect 21416 32348 21422 32360
rect 21910 32348 21916 32360
rect 21416 32320 21916 32348
rect 21416 32308 21422 32320
rect 21910 32308 21916 32320
rect 21968 32308 21974 32360
rect 22020 32348 22048 32388
rect 22094 32376 22100 32428
rect 22152 32416 22158 32428
rect 22554 32416 22560 32428
rect 22152 32388 22197 32416
rect 22515 32388 22560 32416
rect 22152 32376 22158 32388
rect 22554 32376 22560 32388
rect 22612 32376 22618 32428
rect 22747 32416 22775 32456
rect 22824 32453 22836 32487
rect 22870 32484 22882 32487
rect 23290 32484 23296 32496
rect 22870 32456 23296 32484
rect 22870 32453 22882 32456
rect 22824 32447 22882 32453
rect 23290 32444 23296 32456
rect 23348 32444 23354 32496
rect 26510 32484 26516 32496
rect 24412 32456 26516 32484
rect 23566 32416 23572 32428
rect 22747 32388 23572 32416
rect 23566 32376 23572 32388
rect 23624 32376 23630 32428
rect 24412 32425 24440 32456
rect 26510 32444 26516 32456
rect 26568 32444 26574 32496
rect 24670 32425 24676 32428
rect 24397 32419 24455 32425
rect 24397 32385 24409 32419
rect 24443 32385 24455 32419
rect 24664 32416 24676 32425
rect 24631 32388 24676 32416
rect 24397 32379 24455 32385
rect 24664 32379 24676 32388
rect 24670 32376 24676 32379
rect 24728 32376 24734 32428
rect 26421 32419 26479 32425
rect 26421 32385 26433 32419
rect 26467 32416 26479 32419
rect 26786 32416 26792 32428
rect 26467 32388 26792 32416
rect 26467 32385 26479 32388
rect 26421 32379 26479 32385
rect 26786 32376 26792 32388
rect 26844 32376 26850 32428
rect 27157 32419 27215 32425
rect 27157 32385 27169 32419
rect 27203 32416 27215 32419
rect 27522 32416 27528 32428
rect 27203 32388 27528 32416
rect 27203 32385 27215 32388
rect 27157 32379 27215 32385
rect 27522 32376 27528 32388
rect 27580 32376 27586 32428
rect 28258 32425 28264 32428
rect 28215 32419 28264 32425
rect 28215 32385 28227 32419
rect 28261 32385 28264 32419
rect 28215 32379 28264 32385
rect 28258 32376 28264 32379
rect 28316 32376 28322 32428
rect 29454 32416 29460 32428
rect 29415 32388 29460 32416
rect 29454 32376 29460 32388
rect 29512 32376 29518 32428
rect 29564 32388 29868 32416
rect 22189 32351 22247 32357
rect 22189 32348 22201 32351
rect 22020 32320 22201 32348
rect 22189 32317 22201 32320
rect 22235 32317 22247 32351
rect 22189 32311 22247 32317
rect 27341 32351 27399 32357
rect 27341 32317 27353 32351
rect 27387 32317 27399 32351
rect 28077 32351 28135 32357
rect 28077 32348 28089 32351
rect 27341 32311 27399 32317
rect 27632 32320 28089 32348
rect 21821 32283 21879 32289
rect 20918 32252 21680 32280
rect 19521 32243 19579 32249
rect 12894 32212 12900 32224
rect 12636 32184 12900 32212
rect 12529 32175 12587 32181
rect 12894 32172 12900 32184
rect 12952 32172 12958 32224
rect 14458 32172 14464 32224
rect 14516 32212 14522 32224
rect 17954 32212 17960 32224
rect 14516 32184 17960 32212
rect 14516 32172 14522 32184
rect 17954 32172 17960 32184
rect 18012 32172 18018 32224
rect 19153 32215 19211 32221
rect 19153 32181 19165 32215
rect 19199 32212 19211 32215
rect 19426 32212 19432 32224
rect 19199 32184 19432 32212
rect 19199 32181 19211 32184
rect 19153 32175 19211 32181
rect 19426 32172 19432 32184
rect 19484 32172 19490 32224
rect 19702 32172 19708 32224
rect 19760 32212 19766 32224
rect 20714 32212 20720 32224
rect 19760 32184 20720 32212
rect 19760 32172 19766 32184
rect 20714 32172 20720 32184
rect 20772 32172 20778 32224
rect 20990 32212 20996 32224
rect 20951 32184 20996 32212
rect 20990 32172 20996 32184
rect 21048 32172 21054 32224
rect 21652 32221 21680 32252
rect 21821 32249 21833 32283
rect 21867 32280 21879 32283
rect 22462 32280 22468 32292
rect 21867 32252 22468 32280
rect 21867 32249 21879 32252
rect 21821 32243 21879 32249
rect 22462 32240 22468 32252
rect 22520 32240 22526 32292
rect 23934 32280 23940 32292
rect 23895 32252 23940 32280
rect 23934 32240 23940 32252
rect 23992 32240 23998 32292
rect 27356 32280 27384 32311
rect 27632 32292 27660 32320
rect 28077 32317 28089 32320
rect 28123 32317 28135 32351
rect 28077 32311 28135 32317
rect 28353 32351 28411 32357
rect 28353 32317 28365 32351
rect 28399 32348 28411 32351
rect 29564 32348 29592 32388
rect 28399 32320 29592 32348
rect 28399 32317 28411 32320
rect 28353 32311 28411 32317
rect 29638 32308 29644 32360
rect 29696 32348 29702 32360
rect 29840 32348 29868 32388
rect 30374 32348 30380 32360
rect 29696 32320 29741 32348
rect 29840 32320 30236 32348
rect 30335 32320 30380 32348
rect 29696 32308 29702 32320
rect 27522 32280 27528 32292
rect 27356 32252 27528 32280
rect 27522 32240 27528 32252
rect 27580 32240 27586 32292
rect 27614 32240 27620 32292
rect 27672 32240 27678 32292
rect 27801 32283 27859 32289
rect 27801 32249 27813 32283
rect 27847 32249 27859 32283
rect 29822 32280 29828 32292
rect 27801 32243 27859 32249
rect 28920 32252 29828 32280
rect 21637 32215 21695 32221
rect 21637 32181 21649 32215
rect 21683 32212 21695 32215
rect 21910 32212 21916 32224
rect 21683 32184 21916 32212
rect 21683 32181 21695 32184
rect 21637 32175 21695 32181
rect 21910 32172 21916 32184
rect 21968 32172 21974 32224
rect 22189 32215 22247 32221
rect 22189 32181 22201 32215
rect 22235 32212 22247 32215
rect 23474 32212 23480 32224
rect 22235 32184 23480 32212
rect 22235 32181 22247 32184
rect 22189 32175 22247 32181
rect 23474 32172 23480 32184
rect 23532 32172 23538 32224
rect 25777 32215 25835 32221
rect 25777 32181 25789 32215
rect 25823 32212 25835 32215
rect 25866 32212 25872 32224
rect 25823 32184 25872 32212
rect 25823 32181 25835 32184
rect 25777 32175 25835 32181
rect 25866 32172 25872 32184
rect 25924 32172 25930 32224
rect 26234 32212 26240 32224
rect 26195 32184 26240 32212
rect 26234 32172 26240 32184
rect 26292 32172 26298 32224
rect 27816 32212 27844 32243
rect 28920 32212 28948 32252
rect 29822 32240 29828 32252
rect 29880 32280 29886 32292
rect 30101 32283 30159 32289
rect 30101 32280 30113 32283
rect 29880 32252 30113 32280
rect 29880 32240 29886 32252
rect 30101 32249 30113 32252
rect 30147 32249 30159 32283
rect 30101 32243 30159 32249
rect 27816 32184 28948 32212
rect 28997 32215 29055 32221
rect 28997 32181 29009 32215
rect 29043 32212 29055 32215
rect 29086 32212 29092 32224
rect 29043 32184 29092 32212
rect 29043 32181 29055 32184
rect 28997 32175 29055 32181
rect 29086 32172 29092 32184
rect 29144 32172 29150 32224
rect 30208 32212 30236 32320
rect 30374 32308 30380 32320
rect 30432 32308 30438 32360
rect 30466 32308 30472 32360
rect 30524 32357 30530 32360
rect 30524 32351 30552 32357
rect 30540 32317 30552 32351
rect 30524 32311 30552 32317
rect 30524 32308 30530 32311
rect 30650 32308 30656 32360
rect 30708 32348 30714 32360
rect 30708 32320 30753 32348
rect 30708 32308 30714 32320
rect 30374 32212 30380 32224
rect 30208 32184 30380 32212
rect 30374 32172 30380 32184
rect 30432 32212 30438 32224
rect 30650 32212 30656 32224
rect 30432 32184 30656 32212
rect 30432 32172 30438 32184
rect 30650 32172 30656 32184
rect 30708 32172 30714 32224
rect 1104 32122 32016 32144
rect 1104 32070 2136 32122
rect 2188 32070 12440 32122
rect 12492 32070 22744 32122
rect 22796 32070 32016 32122
rect 1104 32048 32016 32070
rect 2406 32008 2412 32020
rect 2367 31980 2412 32008
rect 2406 31968 2412 31980
rect 2464 31968 2470 32020
rect 2958 31968 2964 32020
rect 3016 32008 3022 32020
rect 3789 32011 3847 32017
rect 3789 32008 3801 32011
rect 3016 31980 3801 32008
rect 3016 31968 3022 31980
rect 3789 31977 3801 31980
rect 3835 31977 3847 32011
rect 3789 31971 3847 31977
rect 7561 32011 7619 32017
rect 7561 31977 7573 32011
rect 7607 32008 7619 32011
rect 8938 32008 8944 32020
rect 7607 31980 8944 32008
rect 7607 31977 7619 31980
rect 7561 31971 7619 31977
rect 8938 31968 8944 31980
rect 8996 32008 9002 32020
rect 9585 32011 9643 32017
rect 9585 32008 9597 32011
rect 8996 31980 9597 32008
rect 8996 31968 9002 31980
rect 9585 31977 9597 31980
rect 9631 31977 9643 32011
rect 9585 31971 9643 31977
rect 10873 32011 10931 32017
rect 10873 31977 10885 32011
rect 10919 32008 10931 32011
rect 11698 32008 11704 32020
rect 10919 31980 11704 32008
rect 10919 31977 10931 31980
rect 10873 31971 10931 31977
rect 11698 31968 11704 31980
rect 11756 31968 11762 32020
rect 11974 31968 11980 32020
rect 12032 32008 12038 32020
rect 13449 32011 13507 32017
rect 13449 32008 13461 32011
rect 12032 31980 13461 32008
rect 12032 31968 12038 31980
rect 13449 31977 13461 31980
rect 13495 32008 13507 32011
rect 20346 32008 20352 32020
rect 13495 31980 20352 32008
rect 13495 31977 13507 31980
rect 13449 31971 13507 31977
rect 20346 31968 20352 31980
rect 20404 31968 20410 32020
rect 20993 32011 21051 32017
rect 20993 31977 21005 32011
rect 21039 32008 21051 32011
rect 21174 32008 21180 32020
rect 21039 31980 21180 32008
rect 21039 31977 21051 31980
rect 20993 31971 21051 31977
rect 21174 31968 21180 31980
rect 21232 32008 21238 32020
rect 21232 31980 22497 32008
rect 21232 31968 21238 31980
rect 2774 31900 2780 31952
rect 2832 31940 2838 31952
rect 2832 31912 3924 31940
rect 2832 31900 2838 31912
rect 1949 31807 2007 31813
rect 1949 31773 1961 31807
rect 1995 31804 2007 31807
rect 2038 31804 2044 31816
rect 1995 31776 2044 31804
rect 1995 31773 2007 31776
rect 1949 31767 2007 31773
rect 2038 31764 2044 31776
rect 2096 31764 2102 31816
rect 2593 31807 2651 31813
rect 2593 31773 2605 31807
rect 2639 31804 2651 31807
rect 2682 31804 2688 31816
rect 2639 31776 2688 31804
rect 2639 31773 2651 31776
rect 2593 31767 2651 31773
rect 2682 31764 2688 31776
rect 2740 31764 2746 31816
rect 2866 31764 2872 31816
rect 2924 31804 2930 31816
rect 2924 31776 2969 31804
rect 2924 31764 2930 31776
rect 0 31736 800 31750
rect 1765 31739 1823 31745
rect 1765 31736 1777 31739
rect 0 31708 1777 31736
rect 0 31694 800 31708
rect 1765 31705 1777 31708
rect 1811 31705 1823 31739
rect 3896 31736 3924 31912
rect 4062 31900 4068 31952
rect 4120 31940 4126 31952
rect 6822 31940 6828 31952
rect 4120 31912 6828 31940
rect 4120 31900 4126 31912
rect 6822 31900 6828 31912
rect 6880 31900 6886 31952
rect 7101 31943 7159 31949
rect 7101 31909 7113 31943
rect 7147 31940 7159 31943
rect 9033 31943 9091 31949
rect 7147 31912 8248 31940
rect 7147 31909 7159 31912
rect 7101 31903 7159 31909
rect 4982 31872 4988 31884
rect 4943 31844 4988 31872
rect 4982 31832 4988 31844
rect 5040 31832 5046 31884
rect 5261 31875 5319 31881
rect 5261 31872 5273 31875
rect 5184 31844 5273 31872
rect 3973 31807 4031 31813
rect 3973 31773 3985 31807
rect 4019 31804 4031 31807
rect 4154 31804 4160 31816
rect 4019 31776 4160 31804
rect 4019 31773 4031 31776
rect 3973 31767 4031 31773
rect 4154 31764 4160 31776
rect 4212 31764 4218 31816
rect 4246 31764 4252 31816
rect 4304 31804 4310 31816
rect 4433 31807 4491 31813
rect 4304 31776 4349 31804
rect 4304 31764 4310 31776
rect 4433 31773 4445 31807
rect 4479 31804 4491 31807
rect 4614 31804 4620 31816
rect 4479 31776 4620 31804
rect 4479 31773 4491 31776
rect 4433 31767 4491 31773
rect 4614 31764 4620 31776
rect 4672 31764 4678 31816
rect 5184 31736 5212 31844
rect 5261 31841 5273 31844
rect 5307 31872 5319 31875
rect 6086 31872 6092 31884
rect 5307 31844 6092 31872
rect 5307 31841 5319 31844
rect 5261 31835 5319 31841
rect 6086 31832 6092 31844
rect 6144 31832 6150 31884
rect 6362 31832 6368 31884
rect 6420 31872 6426 31884
rect 6420 31844 7604 31872
rect 6420 31832 6426 31844
rect 6454 31804 6460 31816
rect 6415 31776 6460 31804
rect 6454 31764 6460 31776
rect 6512 31764 6518 31816
rect 6546 31764 6552 31816
rect 6604 31804 6610 31816
rect 6748 31813 6776 31844
rect 6733 31807 6791 31813
rect 6604 31776 6649 31804
rect 6604 31764 6610 31776
rect 6733 31773 6745 31807
rect 6779 31773 6791 31807
rect 6733 31767 6791 31773
rect 6822 31764 6828 31816
rect 6880 31804 6886 31816
rect 6963 31807 7021 31813
rect 6880 31776 6925 31804
rect 6880 31764 6886 31776
rect 6963 31773 6975 31807
rect 7009 31804 7021 31807
rect 7009 31776 7236 31804
rect 7009 31773 7021 31776
rect 6963 31767 7021 31773
rect 3896 31708 5212 31736
rect 7208 31736 7236 31776
rect 7466 31736 7472 31748
rect 7208 31708 7472 31736
rect 1765 31699 1823 31705
rect 7466 31696 7472 31708
rect 7524 31696 7530 31748
rect 7576 31736 7604 31844
rect 7650 31832 7656 31884
rect 7708 31872 7714 31884
rect 7837 31875 7895 31881
rect 7837 31872 7849 31875
rect 7708 31844 7849 31872
rect 7708 31832 7714 31844
rect 7837 31841 7849 31844
rect 7883 31841 7895 31875
rect 8018 31872 8024 31884
rect 7979 31844 8024 31872
rect 7837 31835 7895 31841
rect 8018 31832 8024 31844
rect 8076 31832 8082 31884
rect 7742 31804 7748 31816
rect 7703 31776 7748 31804
rect 7742 31764 7748 31776
rect 7800 31764 7806 31816
rect 7926 31764 7932 31816
rect 7984 31804 7990 31816
rect 8220 31813 8248 31912
rect 9033 31909 9045 31943
rect 9079 31940 9091 31943
rect 12437 31943 12495 31949
rect 12437 31940 12449 31943
rect 9079 31912 12449 31940
rect 9079 31909 9091 31912
rect 9033 31903 9091 31909
rect 9217 31875 9275 31881
rect 9217 31841 9229 31875
rect 9263 31872 9275 31875
rect 10689 31875 10747 31881
rect 10689 31872 10701 31875
rect 9263 31844 10701 31872
rect 9263 31841 9275 31844
rect 9217 31835 9275 31841
rect 10689 31841 10701 31844
rect 10735 31841 10747 31875
rect 10689 31835 10747 31841
rect 8205 31807 8263 31813
rect 7984 31776 8029 31804
rect 7984 31764 7990 31776
rect 8205 31773 8217 31807
rect 8251 31773 8263 31807
rect 8205 31767 8263 31773
rect 8294 31764 8300 31816
rect 8352 31804 8358 31816
rect 9493 31807 9551 31813
rect 9493 31804 9505 31807
rect 8352 31776 9505 31804
rect 8352 31764 8358 31776
rect 9493 31773 9505 31776
rect 9539 31773 9551 31807
rect 9769 31807 9827 31813
rect 9769 31804 9781 31807
rect 9493 31767 9551 31773
rect 9692 31776 9781 31804
rect 8018 31736 8024 31748
rect 7576 31708 8024 31736
rect 8018 31696 8024 31708
rect 8076 31696 8082 31748
rect 9306 31736 9312 31748
rect 9267 31708 9312 31736
rect 9306 31696 9312 31708
rect 9364 31696 9370 31748
rect 9398 31696 9404 31748
rect 9456 31736 9462 31748
rect 9692 31736 9720 31776
rect 9769 31773 9781 31776
rect 9815 31773 9827 31807
rect 9769 31767 9827 31773
rect 10321 31807 10379 31813
rect 10321 31773 10333 31807
rect 10367 31804 10379 31807
rect 10502 31804 10508 31816
rect 10367 31776 10401 31804
rect 10463 31776 10508 31804
rect 10367 31773 10379 31776
rect 10321 31767 10379 31773
rect 9456 31708 9720 31736
rect 10336 31736 10364 31767
rect 10502 31764 10508 31776
rect 10560 31764 10566 31816
rect 11348 31813 11376 31912
rect 12437 31909 12449 31912
rect 12483 31909 12495 31943
rect 12437 31903 12495 31909
rect 12529 31943 12587 31949
rect 12529 31909 12541 31943
rect 12575 31940 12587 31943
rect 12710 31940 12716 31952
rect 12575 31912 12716 31940
rect 12575 31909 12587 31912
rect 12529 31903 12587 31909
rect 12710 31900 12716 31912
rect 12768 31900 12774 31952
rect 12802 31900 12808 31952
rect 12860 31940 12866 31952
rect 14182 31940 14188 31952
rect 12860 31912 12931 31940
rect 14143 31912 14188 31940
rect 12860 31900 12866 31912
rect 12158 31872 12164 31884
rect 12119 31844 12164 31872
rect 12158 31832 12164 31844
rect 12216 31832 12222 31884
rect 10873 31807 10931 31813
rect 10873 31804 10885 31807
rect 10612 31776 10885 31804
rect 10612 31736 10640 31776
rect 10873 31773 10885 31776
rect 10919 31773 10931 31807
rect 10873 31767 10931 31773
rect 11333 31807 11391 31813
rect 11333 31773 11345 31807
rect 11379 31773 11391 31807
rect 11333 31767 11391 31773
rect 11609 31807 11667 31813
rect 11609 31773 11621 31807
rect 11655 31804 11667 31807
rect 12066 31804 12072 31816
rect 11655 31776 12072 31804
rect 11655 31773 11667 31776
rect 11609 31767 11667 31773
rect 12066 31764 12072 31776
rect 12124 31764 12130 31816
rect 12345 31807 12403 31813
rect 12345 31804 12357 31807
rect 12268 31776 12357 31804
rect 10336 31708 10640 31736
rect 9456 31696 9462 31708
rect 11882 31696 11888 31748
rect 11940 31736 11946 31748
rect 12268 31736 12296 31776
rect 12345 31773 12357 31776
rect 12391 31773 12403 31807
rect 12345 31767 12403 31773
rect 12620 31807 12678 31813
rect 12620 31773 12632 31807
rect 12666 31782 12678 31807
rect 12710 31782 12716 31816
rect 12666 31773 12716 31782
rect 12620 31767 12716 31773
rect 12636 31764 12716 31767
rect 12768 31764 12774 31816
rect 12817 31807 12875 31813
rect 12817 31773 12829 31807
rect 12863 31804 12875 31807
rect 12903 31804 12931 31912
rect 14182 31900 14188 31912
rect 14240 31900 14246 31952
rect 15194 31940 15200 31952
rect 14660 31912 15200 31940
rect 13354 31804 13360 31816
rect 12863 31776 12931 31804
rect 13315 31776 13360 31804
rect 12863 31773 12875 31776
rect 12817 31767 12875 31773
rect 13354 31764 13360 31776
rect 13412 31764 13418 31816
rect 14366 31804 14372 31816
rect 14327 31776 14372 31804
rect 14366 31764 14372 31776
rect 14424 31764 14430 31816
rect 14660 31813 14688 31912
rect 15194 31900 15200 31912
rect 15252 31900 15258 31952
rect 17218 31940 17224 31952
rect 17179 31912 17224 31940
rect 17218 31900 17224 31912
rect 17276 31900 17282 31952
rect 17862 31900 17868 31952
rect 17920 31940 17926 31952
rect 18417 31943 18475 31949
rect 18417 31940 18429 31943
rect 17920 31912 18429 31940
rect 17920 31900 17926 31912
rect 18417 31909 18429 31912
rect 18463 31909 18475 31943
rect 18417 31903 18475 31909
rect 21542 31900 21548 31952
rect 21600 31940 21606 31952
rect 22189 31943 22247 31949
rect 22189 31940 22201 31943
rect 21600 31912 22201 31940
rect 21600 31900 21606 31912
rect 22189 31909 22201 31912
rect 22235 31909 22247 31943
rect 22189 31903 22247 31909
rect 22370 31900 22376 31952
rect 22428 31900 22434 31952
rect 22469 31940 22497 31980
rect 22922 31968 22928 32020
rect 22980 32008 22986 32020
rect 23201 32011 23259 32017
rect 23201 32008 23213 32011
rect 22980 31980 23213 32008
rect 22980 31968 22986 31980
rect 23201 31977 23213 31980
rect 23247 31977 23259 32011
rect 23201 31971 23259 31977
rect 24946 31968 24952 32020
rect 25004 32008 25010 32020
rect 25409 32011 25467 32017
rect 25409 32008 25421 32011
rect 25004 31980 25421 32008
rect 25004 31968 25010 31980
rect 25409 31977 25421 31980
rect 25455 31977 25467 32011
rect 25409 31971 25467 31977
rect 26234 31968 26240 32020
rect 26292 32008 26298 32020
rect 26292 31980 27568 32008
rect 26292 31968 26298 31980
rect 24857 31943 24915 31949
rect 22469 31912 23244 31940
rect 15102 31832 15108 31884
rect 15160 31872 15166 31884
rect 15841 31875 15899 31881
rect 15841 31872 15853 31875
rect 15160 31844 15853 31872
rect 15160 31832 15166 31844
rect 15841 31841 15853 31844
rect 15887 31841 15899 31875
rect 15841 31835 15899 31841
rect 16022 31832 16028 31884
rect 16080 31872 16086 31884
rect 16761 31875 16819 31881
rect 16761 31872 16773 31875
rect 16080 31844 16773 31872
rect 16080 31832 16086 31844
rect 16761 31841 16773 31844
rect 16807 31841 16819 31875
rect 16761 31835 16819 31841
rect 16942 31832 16948 31884
rect 17000 31872 17006 31884
rect 17773 31875 17831 31881
rect 17773 31872 17785 31875
rect 17000 31844 17785 31872
rect 17000 31832 17006 31844
rect 17773 31841 17785 31844
rect 17819 31872 17831 31875
rect 18138 31872 18144 31884
rect 17819 31844 18144 31872
rect 17819 31841 17831 31844
rect 17773 31835 17831 31841
rect 18138 31832 18144 31844
rect 18196 31832 18202 31884
rect 21085 31875 21143 31881
rect 18432 31844 19380 31872
rect 14645 31807 14703 31813
rect 14645 31773 14657 31807
rect 14691 31773 14703 31807
rect 14826 31804 14832 31816
rect 14787 31776 14832 31804
rect 14645 31767 14703 31773
rect 14826 31764 14832 31776
rect 14884 31764 14890 31816
rect 15654 31804 15660 31816
rect 15615 31776 15660 31804
rect 15654 31764 15660 31776
rect 15712 31764 15718 31816
rect 15933 31807 15991 31813
rect 15933 31773 15945 31807
rect 15979 31804 15991 31807
rect 16574 31804 16580 31816
rect 15979 31776 16436 31804
rect 16535 31776 16580 31804
rect 15979 31773 15991 31776
rect 15933 31767 15991 31773
rect 12636 31754 12756 31764
rect 16114 31736 16120 31748
rect 11940 31708 12296 31736
rect 15304 31708 16120 31736
rect 11940 31696 11946 31708
rect 7558 31628 7564 31680
rect 7616 31668 7622 31680
rect 9030 31668 9036 31680
rect 7616 31640 9036 31668
rect 7616 31628 7622 31640
rect 9030 31628 9036 31640
rect 9088 31628 9094 31680
rect 11422 31668 11428 31680
rect 11383 31640 11428 31668
rect 11422 31628 11428 31640
rect 11480 31668 11486 31680
rect 15304 31668 15332 31708
rect 16114 31696 16120 31708
rect 16172 31696 16178 31748
rect 15470 31668 15476 31680
rect 11480 31640 15332 31668
rect 15431 31640 15476 31668
rect 11480 31628 11486 31640
rect 15470 31628 15476 31640
rect 15528 31628 15534 31680
rect 16408 31668 16436 31776
rect 16574 31764 16580 31776
rect 16632 31764 16638 31816
rect 18322 31804 18328 31816
rect 16868 31776 18328 31804
rect 16868 31668 16896 31776
rect 18322 31764 18328 31776
rect 18380 31764 18386 31816
rect 18432 31813 18460 31844
rect 18417 31807 18475 31813
rect 18417 31773 18429 31807
rect 18463 31773 18475 31807
rect 18417 31767 18475 31773
rect 18693 31807 18751 31813
rect 18693 31773 18705 31807
rect 18739 31804 18751 31807
rect 19242 31804 19248 31816
rect 18739 31776 19012 31804
rect 19203 31776 19248 31804
rect 18739 31773 18751 31776
rect 18693 31767 18751 31773
rect 17770 31736 17776 31748
rect 17144 31708 17776 31736
rect 16408 31640 16896 31668
rect 17034 31628 17040 31680
rect 17092 31668 17098 31680
rect 17144 31668 17172 31708
rect 17770 31696 17776 31708
rect 17828 31696 17834 31748
rect 18984 31736 19012 31776
rect 19242 31764 19248 31776
rect 19300 31764 19306 31816
rect 19352 31804 19380 31844
rect 21085 31841 21097 31875
rect 21131 31872 21143 31875
rect 22388 31872 22416 31900
rect 21131 31844 22416 31872
rect 22465 31875 22523 31881
rect 21131 31841 21143 31844
rect 21085 31835 21143 31841
rect 22465 31841 22477 31875
rect 22511 31841 22523 31875
rect 22465 31835 22523 31841
rect 19518 31813 19524 31816
rect 19352 31776 19472 31804
rect 19334 31736 19340 31748
rect 18984 31708 19340 31736
rect 19334 31696 19340 31708
rect 19392 31696 19398 31748
rect 19444 31736 19472 31776
rect 19512 31767 19524 31813
rect 19576 31804 19582 31816
rect 19576 31776 19612 31804
rect 19518 31764 19524 31767
rect 19576 31764 19582 31776
rect 20714 31764 20720 31816
rect 20772 31804 20778 31816
rect 21361 31807 21419 31813
rect 21361 31804 21373 31807
rect 20772 31776 21373 31804
rect 20772 31764 20778 31776
rect 21361 31773 21373 31776
rect 21407 31773 21419 31807
rect 21361 31767 21419 31773
rect 21453 31807 21511 31813
rect 21453 31773 21465 31807
rect 21499 31773 21511 31807
rect 21453 31767 21511 31773
rect 19444 31708 21036 31736
rect 17092 31640 17172 31668
rect 17092 31628 17098 31640
rect 17402 31628 17408 31680
rect 17460 31668 17466 31680
rect 17589 31671 17647 31677
rect 17589 31668 17601 31671
rect 17460 31640 17601 31668
rect 17460 31628 17466 31640
rect 17589 31637 17601 31640
rect 17635 31637 17647 31671
rect 17589 31631 17647 31637
rect 17681 31671 17739 31677
rect 17681 31637 17693 31671
rect 17727 31668 17739 31671
rect 17954 31668 17960 31680
rect 17727 31640 17960 31668
rect 17727 31637 17739 31640
rect 17681 31631 17739 31637
rect 17954 31628 17960 31640
rect 18012 31668 18018 31680
rect 18506 31668 18512 31680
rect 18012 31640 18512 31668
rect 18012 31628 18018 31640
rect 18506 31628 18512 31640
rect 18564 31628 18570 31680
rect 18601 31671 18659 31677
rect 18601 31637 18613 31671
rect 18647 31668 18659 31671
rect 19058 31668 19064 31680
rect 18647 31640 19064 31668
rect 18647 31637 18659 31640
rect 18601 31631 18659 31637
rect 19058 31628 19064 31640
rect 19116 31628 19122 31680
rect 20254 31628 20260 31680
rect 20312 31668 20318 31680
rect 21008 31677 21036 31708
rect 20625 31671 20683 31677
rect 20625 31668 20637 31671
rect 20312 31640 20637 31668
rect 20312 31628 20318 31640
rect 20625 31637 20637 31640
rect 20671 31637 20683 31671
rect 20625 31631 20683 31637
rect 20993 31671 21051 31677
rect 20993 31637 21005 31671
rect 21039 31668 21051 31671
rect 21082 31668 21088 31680
rect 21039 31640 21088 31668
rect 21039 31637 21051 31640
rect 20993 31631 21051 31637
rect 21082 31628 21088 31640
rect 21140 31628 21146 31680
rect 21358 31628 21364 31680
rect 21416 31668 21422 31680
rect 21468 31668 21496 31767
rect 21542 31764 21548 31816
rect 21600 31804 21606 31816
rect 21600 31776 21645 31804
rect 21600 31764 21606 31776
rect 21726 31764 21732 31816
rect 21784 31804 21790 31816
rect 22370 31804 22376 31816
rect 21784 31776 21829 31804
rect 22331 31776 22376 31804
rect 21784 31764 21790 31776
rect 22370 31764 22376 31776
rect 22428 31764 22434 31816
rect 22469 31748 22497 31835
rect 22646 31832 22652 31884
rect 22704 31872 22710 31884
rect 22704 31844 22749 31872
rect 22704 31832 22710 31844
rect 22548 31807 22606 31813
rect 22548 31773 22560 31807
rect 22594 31798 22606 31807
rect 22830 31804 22836 31816
rect 22747 31798 22836 31804
rect 22594 31776 22836 31798
rect 22594 31773 22775 31776
rect 22548 31770 22775 31773
rect 22548 31767 22606 31770
rect 22830 31764 22836 31776
rect 22888 31764 22894 31816
rect 23216 31813 23244 31912
rect 24857 31909 24869 31943
rect 24903 31940 24915 31943
rect 25682 31940 25688 31952
rect 24903 31912 25688 31940
rect 24903 31909 24915 31912
rect 24857 31903 24915 31909
rect 25682 31900 25688 31912
rect 25740 31900 25746 31952
rect 27540 31940 27568 31980
rect 27614 31968 27620 32020
rect 27672 32008 27678 32020
rect 27893 32011 27951 32017
rect 27893 32008 27905 32011
rect 27672 31980 27905 32008
rect 27672 31968 27678 31980
rect 27893 31977 27905 31980
rect 27939 31977 27951 32011
rect 28534 32008 28540 32020
rect 28495 31980 28540 32008
rect 27893 31971 27951 31977
rect 28534 31968 28540 31980
rect 28592 31968 28598 32020
rect 29730 32008 29736 32020
rect 28828 31980 29736 32008
rect 28828 31940 28856 31980
rect 29730 31968 29736 31980
rect 29788 31968 29794 32020
rect 27540 31912 28856 31940
rect 28902 31900 28908 31952
rect 28960 31940 28966 31952
rect 30469 31943 30527 31949
rect 30469 31940 30481 31943
rect 28960 31912 30481 31940
rect 28960 31900 28966 31912
rect 30469 31909 30481 31912
rect 30515 31909 30527 31943
rect 30469 31903 30527 31909
rect 25498 31872 25504 31884
rect 24780 31844 25504 31872
rect 23201 31807 23259 31813
rect 23201 31773 23213 31807
rect 23247 31773 23259 31807
rect 23474 31804 23480 31816
rect 23435 31776 23480 31804
rect 23201 31767 23259 31773
rect 23474 31764 23480 31776
rect 23532 31764 23538 31816
rect 24780 31813 24808 31844
rect 25498 31832 25504 31844
rect 25556 31832 25562 31884
rect 26326 31872 26332 31884
rect 25884 31844 26332 31872
rect 25884 31813 25912 31844
rect 26326 31832 26332 31844
rect 26384 31832 26390 31884
rect 26510 31872 26516 31884
rect 26471 31844 26516 31872
rect 26510 31832 26516 31844
rect 26568 31832 26574 31884
rect 27522 31832 27528 31884
rect 27580 31872 27586 31884
rect 28997 31875 29055 31881
rect 28997 31872 29009 31875
rect 27580 31844 29009 31872
rect 27580 31832 27586 31844
rect 28997 31841 29009 31844
rect 29043 31872 29055 31875
rect 29178 31872 29184 31884
rect 29043 31844 29184 31872
rect 29043 31841 29055 31844
rect 28997 31835 29055 31841
rect 29178 31832 29184 31844
rect 29236 31832 29242 31884
rect 30098 31832 30104 31884
rect 30156 31872 30162 31884
rect 30561 31875 30619 31881
rect 30561 31872 30573 31875
rect 30156 31844 30573 31872
rect 30156 31832 30162 31844
rect 30561 31841 30573 31844
rect 30607 31841 30619 31875
rect 30561 31835 30619 31841
rect 24765 31807 24823 31813
rect 24765 31773 24777 31807
rect 24811 31773 24823 31807
rect 24765 31767 24823 31773
rect 25593 31807 25651 31813
rect 25593 31773 25605 31807
rect 25639 31804 25651 31807
rect 25869 31807 25927 31813
rect 25639 31776 25820 31804
rect 25639 31773 25651 31776
rect 25593 31767 25651 31773
rect 22462 31696 22468 31748
rect 22520 31696 22526 31748
rect 25792 31736 25820 31776
rect 25869 31773 25881 31807
rect 25915 31773 25927 31807
rect 25869 31767 25927 31773
rect 25958 31764 25964 31816
rect 26016 31804 26022 31816
rect 26053 31807 26111 31813
rect 26053 31804 26065 31807
rect 26016 31776 26065 31804
rect 26016 31764 26022 31776
rect 26053 31773 26065 31776
rect 26099 31773 26111 31807
rect 26053 31767 26111 31773
rect 26780 31807 26838 31813
rect 26780 31773 26792 31807
rect 26826 31804 26838 31807
rect 28350 31804 28356 31816
rect 26826 31776 28356 31804
rect 26826 31773 26838 31776
rect 26780 31767 26838 31773
rect 28350 31764 28356 31776
rect 28408 31764 28414 31816
rect 28718 31804 28724 31816
rect 28679 31776 28724 31804
rect 28718 31764 28724 31776
rect 28776 31764 28782 31816
rect 28810 31764 28816 31816
rect 28868 31804 28874 31816
rect 28905 31807 28963 31813
rect 28905 31804 28917 31807
rect 28868 31776 28917 31804
rect 28868 31764 28874 31776
rect 28905 31773 28917 31776
rect 28951 31773 28963 31807
rect 30282 31804 30288 31816
rect 30243 31776 30288 31804
rect 28905 31767 28963 31773
rect 30282 31764 30288 31776
rect 30340 31764 30346 31816
rect 30742 31764 30748 31816
rect 30800 31804 30806 31816
rect 31113 31807 31171 31813
rect 31113 31804 31125 31807
rect 30800 31776 31125 31804
rect 30800 31764 30806 31776
rect 31113 31773 31125 31776
rect 31159 31773 31171 31807
rect 31113 31767 31171 31773
rect 26418 31736 26424 31748
rect 25792 31708 26424 31736
rect 26418 31696 26424 31708
rect 26476 31736 26482 31748
rect 26694 31736 26700 31748
rect 26476 31708 26700 31736
rect 26476 31696 26482 31708
rect 26694 31696 26700 31708
rect 26752 31696 26758 31748
rect 32320 31736 33120 31750
rect 32232 31708 33120 31736
rect 21416 31640 21496 31668
rect 21416 31628 21422 31640
rect 23014 31628 23020 31680
rect 23072 31668 23078 31680
rect 23385 31671 23443 31677
rect 23385 31668 23397 31671
rect 23072 31640 23397 31668
rect 23072 31628 23078 31640
rect 23385 31637 23397 31640
rect 23431 31637 23443 31671
rect 23385 31631 23443 31637
rect 24026 31628 24032 31680
rect 24084 31668 24090 31680
rect 24486 31668 24492 31680
rect 24084 31640 24492 31668
rect 24084 31628 24090 31640
rect 24486 31628 24492 31640
rect 24544 31628 24550 31680
rect 30101 31671 30159 31677
rect 30101 31637 30113 31671
rect 30147 31668 30159 31671
rect 30190 31668 30196 31680
rect 30147 31640 30196 31668
rect 30147 31637 30159 31640
rect 30101 31631 30159 31637
rect 30190 31628 30196 31640
rect 30248 31628 30254 31680
rect 31202 31668 31208 31680
rect 31163 31640 31208 31668
rect 31202 31628 31208 31640
rect 31260 31628 31266 31680
rect 32232 31600 32260 31708
rect 32320 31694 33120 31708
rect 1104 31578 32016 31600
rect 1104 31526 7288 31578
rect 7340 31526 17592 31578
rect 17644 31526 27896 31578
rect 27948 31526 32016 31578
rect 32232 31572 32352 31600
rect 1104 31504 32016 31526
rect 3878 31424 3884 31476
rect 3936 31464 3942 31476
rect 7285 31467 7343 31473
rect 3936 31436 5856 31464
rect 3936 31424 3942 31436
rect 2038 31356 2044 31408
rect 2096 31396 2102 31408
rect 2498 31396 2504 31408
rect 2096 31368 2504 31396
rect 2096 31356 2102 31368
rect 2498 31356 2504 31368
rect 2556 31356 2562 31408
rect 2590 31328 2596 31340
rect 2551 31300 2596 31328
rect 2590 31288 2596 31300
rect 2648 31288 2654 31340
rect 3881 31331 3939 31337
rect 3881 31297 3893 31331
rect 3927 31328 3939 31331
rect 3970 31328 3976 31340
rect 3927 31300 3976 31328
rect 3927 31297 3939 31300
rect 3881 31291 3939 31297
rect 3970 31288 3976 31300
rect 4028 31288 4034 31340
rect 4246 31288 4252 31340
rect 4304 31328 4310 31340
rect 5828 31337 5856 31436
rect 7285 31433 7297 31467
rect 7331 31464 7343 31467
rect 7926 31464 7932 31476
rect 7331 31436 7932 31464
rect 7331 31433 7343 31436
rect 7285 31427 7343 31433
rect 7926 31424 7932 31436
rect 7984 31424 7990 31476
rect 8018 31424 8024 31476
rect 8076 31464 8082 31476
rect 8297 31467 8355 31473
rect 8297 31464 8309 31467
rect 8076 31436 8309 31464
rect 8076 31424 8082 31436
rect 8297 31433 8309 31436
rect 8343 31433 8355 31467
rect 8297 31427 8355 31433
rect 8404 31436 9812 31464
rect 6638 31356 6644 31408
rect 6696 31396 6702 31408
rect 6733 31399 6791 31405
rect 6733 31396 6745 31399
rect 6696 31368 6745 31396
rect 6696 31356 6702 31368
rect 6733 31365 6745 31368
rect 6779 31365 6791 31399
rect 6733 31359 6791 31365
rect 7101 31399 7159 31405
rect 7101 31365 7113 31399
rect 7147 31396 7159 31399
rect 8113 31399 8171 31405
rect 8113 31396 8125 31399
rect 7147 31368 8125 31396
rect 7147 31365 7159 31368
rect 7101 31359 7159 31365
rect 8113 31365 8125 31368
rect 8159 31365 8171 31399
rect 8404 31396 8432 31436
rect 9309 31399 9367 31405
rect 8113 31359 8171 31365
rect 8312 31368 8432 31396
rect 8496 31368 8892 31396
rect 4525 31331 4583 31337
rect 4525 31328 4537 31331
rect 4304 31300 4537 31328
rect 4304 31288 4310 31300
rect 4525 31297 4537 31300
rect 4571 31297 4583 31331
rect 4525 31291 4583 31297
rect 5813 31331 5871 31337
rect 5813 31297 5825 31331
rect 5859 31297 5871 31331
rect 5813 31291 5871 31297
rect 6917 31331 6975 31337
rect 6917 31297 6929 31331
rect 6963 31297 6975 31331
rect 6917 31291 6975 31297
rect 1762 31220 1768 31272
rect 1820 31260 1826 31272
rect 2038 31260 2044 31272
rect 1820 31232 2044 31260
rect 1820 31220 1826 31232
rect 2038 31220 2044 31232
rect 2096 31220 2102 31272
rect 2869 31263 2927 31269
rect 2869 31229 2881 31263
rect 2915 31260 2927 31263
rect 3602 31260 3608 31272
rect 2915 31232 3608 31260
rect 2915 31229 2927 31232
rect 2869 31223 2927 31229
rect 3602 31220 3608 31232
rect 3660 31260 3666 31272
rect 4062 31260 4068 31272
rect 3660 31232 4068 31260
rect 3660 31220 3666 31232
rect 4062 31220 4068 31232
rect 4120 31220 4126 31272
rect 4798 31260 4804 31272
rect 4759 31232 4804 31260
rect 4798 31220 4804 31232
rect 4856 31220 4862 31272
rect 6932 31260 6960 31291
rect 7006 31288 7012 31340
rect 7064 31328 7070 31340
rect 8312 31337 8340 31368
rect 8297 31331 8355 31337
rect 7064 31300 7109 31328
rect 7064 31288 7070 31300
rect 8297 31297 8309 31331
rect 8343 31297 8355 31331
rect 8297 31291 8355 31297
rect 7374 31260 7380 31272
rect 6932 31232 7380 31260
rect 7374 31220 7380 31232
rect 7432 31220 7438 31272
rect 7650 31220 7656 31272
rect 7708 31260 7714 31272
rect 8110 31260 8116 31272
rect 7708 31232 8116 31260
rect 7708 31220 7714 31232
rect 8110 31220 8116 31232
rect 8168 31260 8174 31272
rect 8496 31260 8524 31368
rect 8573 31331 8631 31337
rect 8573 31297 8585 31331
rect 8619 31297 8631 31331
rect 8573 31291 8631 31297
rect 8168 31232 8524 31260
rect 8168 31220 8174 31232
rect 2777 31195 2835 31201
rect 2777 31161 2789 31195
rect 2823 31192 2835 31195
rect 4709 31195 4767 31201
rect 4709 31192 4721 31195
rect 2823 31164 4721 31192
rect 2823 31161 2835 31164
rect 2777 31155 2835 31161
rect 4709 31161 4721 31164
rect 4755 31192 4767 31195
rect 5166 31192 5172 31204
rect 4755 31164 5172 31192
rect 4755 31161 4767 31164
rect 4709 31155 4767 31161
rect 5166 31152 5172 31164
rect 5224 31152 5230 31204
rect 7006 31152 7012 31204
rect 7064 31192 7070 31204
rect 8588 31192 8616 31291
rect 8662 31220 8668 31272
rect 8720 31260 8726 31272
rect 8864 31260 8892 31368
rect 9309 31365 9321 31399
rect 9355 31396 9367 31399
rect 9582 31396 9588 31408
rect 9355 31368 9588 31396
rect 9355 31365 9367 31368
rect 9309 31359 9367 31365
rect 9582 31356 9588 31368
rect 9640 31356 9646 31408
rect 9784 31396 9812 31436
rect 9858 31424 9864 31476
rect 9916 31464 9922 31476
rect 9953 31467 10011 31473
rect 9953 31464 9965 31467
rect 9916 31436 9965 31464
rect 9916 31424 9922 31436
rect 9953 31433 9965 31436
rect 9999 31433 10011 31467
rect 9953 31427 10011 31433
rect 11882 31424 11888 31476
rect 11940 31464 11946 31476
rect 13262 31464 13268 31476
rect 11940 31436 13032 31464
rect 13223 31436 13268 31464
rect 11940 31424 11946 31436
rect 11698 31396 11704 31408
rect 9784 31368 11704 31396
rect 11698 31356 11704 31368
rect 11756 31356 11762 31408
rect 11974 31396 11980 31408
rect 11935 31368 11980 31396
rect 11974 31356 11980 31368
rect 12032 31356 12038 31408
rect 12636 31368 12940 31396
rect 9769 31331 9827 31337
rect 9769 31297 9781 31331
rect 9815 31297 9827 31331
rect 9769 31291 9827 31297
rect 9677 31263 9735 31269
rect 9677 31260 9689 31263
rect 8720 31232 8765 31260
rect 8864 31232 9689 31260
rect 8720 31220 8726 31232
rect 9677 31229 9689 31232
rect 9723 31229 9735 31263
rect 9784 31260 9812 31291
rect 10042 31288 10048 31340
rect 10100 31328 10106 31340
rect 10597 31331 10655 31337
rect 10597 31328 10609 31331
rect 10100 31300 10609 31328
rect 10100 31288 10106 31300
rect 10597 31297 10609 31300
rect 10643 31297 10655 31331
rect 10597 31291 10655 31297
rect 10873 31331 10931 31337
rect 10873 31297 10885 31331
rect 10919 31328 10931 31331
rect 11054 31328 11060 31340
rect 10919 31300 11060 31328
rect 10919 31297 10931 31300
rect 10873 31291 10931 31297
rect 11054 31288 11060 31300
rect 11112 31288 11118 31340
rect 11146 31260 11152 31272
rect 9784 31232 11152 31260
rect 9677 31223 9735 31229
rect 11146 31220 11152 31232
rect 11204 31220 11210 31272
rect 11790 31220 11796 31272
rect 11848 31260 11854 31272
rect 12636 31260 12664 31368
rect 12802 31260 12808 31272
rect 11848 31232 12664 31260
rect 12728 31232 12808 31260
rect 11848 31220 11854 31232
rect 7064 31164 8616 31192
rect 7064 31152 7070 31164
rect 10594 31152 10600 31204
rect 10652 31192 10658 31204
rect 10652 31164 11008 31192
rect 10652 31152 10658 31164
rect 10980 31136 11008 31164
rect 11882 31152 11888 31204
rect 11940 31192 11946 31204
rect 12728 31201 12756 31232
rect 12802 31220 12808 31232
rect 12860 31220 12866 31272
rect 12912 31260 12940 31368
rect 13004 31328 13032 31436
rect 13262 31424 13268 31436
rect 13320 31424 13326 31476
rect 14277 31467 14335 31473
rect 14277 31433 14289 31467
rect 14323 31464 14335 31467
rect 14642 31464 14648 31476
rect 14323 31436 14648 31464
rect 14323 31433 14335 31436
rect 14277 31427 14335 31433
rect 14642 31424 14648 31436
rect 14700 31424 14706 31476
rect 15289 31467 15347 31473
rect 15289 31433 15301 31467
rect 15335 31464 15347 31467
rect 15654 31464 15660 31476
rect 15335 31436 15660 31464
rect 15335 31433 15347 31436
rect 15289 31427 15347 31433
rect 15654 31424 15660 31436
rect 15712 31424 15718 31476
rect 16114 31424 16120 31476
rect 16172 31464 16178 31476
rect 17221 31467 17279 31473
rect 17221 31464 17233 31467
rect 16172 31436 17233 31464
rect 16172 31424 16178 31436
rect 17221 31433 17233 31436
rect 17267 31433 17279 31467
rect 18417 31467 18475 31473
rect 18417 31464 18429 31467
rect 17221 31427 17279 31433
rect 17788 31436 18429 31464
rect 13081 31399 13139 31405
rect 13081 31365 13093 31399
rect 13127 31396 13139 31399
rect 13127 31368 13308 31396
rect 13127 31365 13139 31368
rect 13081 31359 13139 31365
rect 13280 31340 13308 31368
rect 15194 31356 15200 31408
rect 15252 31396 15258 31408
rect 15252 31368 15792 31396
rect 15252 31356 15258 31368
rect 13170 31328 13176 31340
rect 13004 31300 13176 31328
rect 13170 31288 13176 31300
rect 13228 31288 13234 31340
rect 13262 31288 13268 31340
rect 13320 31288 13326 31340
rect 14274 31288 14280 31340
rect 14332 31328 14338 31340
rect 14461 31331 14519 31337
rect 14461 31328 14473 31331
rect 14332 31300 14473 31328
rect 14332 31288 14338 31300
rect 14461 31297 14473 31300
rect 14507 31297 14519 31331
rect 14461 31291 14519 31297
rect 15286 31288 15292 31340
rect 15344 31328 15350 31340
rect 15473 31331 15531 31337
rect 15473 31328 15485 31331
rect 15344 31300 15485 31328
rect 15344 31288 15350 31300
rect 15473 31297 15485 31300
rect 15519 31297 15531 31331
rect 15473 31291 15531 31297
rect 15654 31288 15660 31340
rect 15712 31328 15718 31340
rect 15764 31337 15792 31368
rect 15749 31331 15807 31337
rect 15749 31328 15761 31331
rect 15712 31300 15761 31328
rect 15712 31288 15718 31300
rect 15749 31297 15761 31300
rect 15795 31297 15807 31331
rect 15930 31328 15936 31340
rect 15891 31300 15936 31328
rect 15749 31291 15807 31297
rect 15930 31288 15936 31300
rect 15988 31328 15994 31340
rect 16298 31328 16304 31340
rect 15988 31300 16304 31328
rect 15988 31288 15994 31300
rect 16298 31288 16304 31300
rect 16356 31288 16362 31340
rect 16850 31328 16856 31340
rect 16811 31300 16856 31328
rect 16850 31288 16856 31300
rect 16908 31288 16914 31340
rect 17310 31288 17316 31340
rect 17368 31328 17374 31340
rect 17788 31337 17816 31436
rect 18417 31433 18429 31436
rect 18463 31433 18475 31467
rect 18966 31464 18972 31476
rect 18927 31436 18972 31464
rect 18417 31427 18475 31433
rect 18966 31424 18972 31436
rect 19024 31424 19030 31476
rect 19058 31424 19064 31476
rect 19116 31464 19122 31476
rect 19334 31464 19340 31476
rect 19116 31436 19340 31464
rect 19116 31424 19122 31436
rect 19334 31424 19340 31436
rect 19392 31424 19398 31476
rect 20901 31467 20959 31473
rect 20901 31433 20913 31467
rect 20947 31464 20959 31467
rect 21542 31464 21548 31476
rect 20947 31436 21548 31464
rect 20947 31433 20959 31436
rect 20901 31427 20959 31433
rect 21542 31424 21548 31436
rect 21600 31424 21606 31476
rect 21818 31464 21824 31476
rect 21779 31436 21824 31464
rect 21818 31424 21824 31436
rect 21876 31424 21882 31476
rect 22094 31424 22100 31476
rect 22152 31464 22158 31476
rect 23842 31464 23848 31476
rect 22152 31436 23848 31464
rect 22152 31424 22158 31436
rect 23842 31424 23848 31436
rect 23900 31464 23906 31476
rect 24305 31467 24363 31473
rect 24305 31464 24317 31467
rect 23900 31436 24317 31464
rect 23900 31424 23906 31436
rect 24305 31433 24317 31436
rect 24351 31433 24363 31467
rect 28350 31464 28356 31476
rect 28311 31436 28356 31464
rect 24305 31427 24363 31433
rect 28350 31424 28356 31436
rect 28408 31424 28414 31476
rect 31110 31424 31116 31476
rect 31168 31464 31174 31476
rect 31294 31464 31300 31476
rect 31168 31436 31300 31464
rect 31168 31424 31174 31436
rect 31294 31424 31300 31436
rect 31352 31424 31358 31476
rect 18064 31368 19472 31396
rect 17589 31331 17647 31337
rect 17589 31328 17601 31331
rect 17368 31300 17601 31328
rect 17368 31288 17374 31300
rect 17589 31297 17601 31300
rect 17635 31297 17647 31331
rect 17589 31291 17647 31297
rect 17773 31331 17831 31337
rect 17773 31297 17785 31331
rect 17819 31297 17831 31331
rect 17773 31291 17831 31297
rect 17954 31288 17960 31340
rect 18012 31328 18018 31340
rect 18064 31337 18092 31368
rect 18049 31331 18107 31337
rect 18049 31328 18061 31331
rect 18012 31300 18061 31328
rect 18012 31288 18018 31300
rect 18049 31297 18061 31300
rect 18095 31297 18107 31331
rect 18049 31291 18107 31297
rect 18230 31288 18236 31340
rect 18288 31328 18294 31340
rect 18417 31331 18475 31337
rect 18288 31300 18381 31328
rect 18288 31288 18294 31300
rect 18417 31297 18429 31331
rect 18463 31328 18475 31331
rect 19150 31328 19156 31340
rect 18463 31300 19156 31328
rect 18463 31297 18475 31300
rect 18417 31291 18475 31297
rect 19150 31288 19156 31300
rect 19208 31288 19214 31340
rect 19444 31337 19472 31368
rect 20438 31356 20444 31408
rect 20496 31396 20502 31408
rect 20717 31399 20775 31405
rect 20717 31396 20729 31399
rect 20496 31368 20729 31396
rect 20496 31356 20502 31368
rect 20717 31365 20729 31368
rect 20763 31396 20775 31399
rect 21726 31396 21732 31408
rect 20763 31368 21732 31396
rect 20763 31365 20775 31368
rect 20717 31359 20775 31365
rect 21726 31356 21732 31368
rect 21784 31396 21790 31408
rect 22462 31396 22468 31408
rect 21784 31368 22468 31396
rect 21784 31356 21790 31368
rect 19429 31331 19487 31337
rect 19429 31297 19441 31331
rect 19475 31297 19487 31331
rect 19610 31328 19616 31340
rect 19571 31300 19616 31328
rect 19429 31291 19487 31297
rect 19610 31288 19616 31300
rect 19668 31328 19674 31340
rect 20254 31328 20260 31340
rect 19668 31300 20260 31328
rect 19668 31288 19674 31300
rect 20254 31288 20260 31300
rect 20312 31288 20318 31340
rect 20530 31328 20536 31340
rect 20491 31300 20536 31328
rect 20530 31288 20536 31300
rect 20588 31288 20594 31340
rect 20990 31288 20996 31340
rect 21048 31328 21054 31340
rect 22296 31337 22324 31368
rect 22462 31356 22468 31368
rect 22520 31356 22526 31408
rect 32324 31396 32352 31572
rect 23216 31368 32352 31396
rect 22005 31331 22063 31337
rect 22005 31328 22017 31331
rect 21048 31300 22017 31328
rect 21048 31288 21054 31300
rect 22005 31297 22017 31300
rect 22051 31297 22063 31331
rect 22005 31291 22063 31297
rect 22281 31331 22339 31337
rect 22281 31297 22293 31331
rect 22327 31297 22339 31331
rect 22281 31291 22339 31297
rect 14090 31260 14096 31272
rect 12912 31232 13952 31260
rect 14051 31232 14096 31260
rect 12713 31195 12771 31201
rect 12713 31192 12725 31195
rect 11940 31164 12725 31192
rect 11940 31152 11946 31164
rect 12713 31161 12725 31164
rect 12759 31161 12771 31195
rect 13630 31192 13636 31204
rect 12713 31155 12771 31161
rect 12820 31164 13636 31192
rect 1762 31084 1768 31136
rect 1820 31124 1826 31136
rect 2409 31127 2467 31133
rect 2409 31124 2421 31127
rect 1820 31096 2421 31124
rect 1820 31084 1826 31096
rect 2409 31093 2421 31096
rect 2455 31093 2467 31127
rect 3694 31124 3700 31136
rect 3655 31096 3700 31124
rect 2409 31087 2467 31093
rect 3694 31084 3700 31096
rect 3752 31084 3758 31136
rect 4338 31124 4344 31136
rect 4299 31096 4344 31124
rect 4338 31084 4344 31096
rect 4396 31084 4402 31136
rect 5629 31127 5687 31133
rect 5629 31093 5641 31127
rect 5675 31124 5687 31127
rect 5810 31124 5816 31136
rect 5675 31096 5816 31124
rect 5675 31093 5687 31096
rect 5629 31087 5687 31093
rect 5810 31084 5816 31096
rect 5868 31084 5874 31136
rect 8113 31127 8171 31133
rect 8113 31093 8125 31127
rect 8159 31124 8171 31127
rect 8662 31124 8668 31136
rect 8159 31096 8668 31124
rect 8159 31093 8171 31096
rect 8113 31087 8171 31093
rect 8662 31084 8668 31096
rect 8720 31084 8726 31136
rect 8846 31084 8852 31136
rect 8904 31124 8910 31136
rect 9401 31127 9459 31133
rect 9401 31124 9413 31127
rect 8904 31096 9413 31124
rect 8904 31084 8910 31096
rect 9401 31093 9413 31096
rect 9447 31093 9459 31127
rect 10410 31124 10416 31136
rect 10371 31096 10416 31124
rect 9401 31087 9459 31093
rect 10410 31084 10416 31096
rect 10468 31084 10474 31136
rect 10502 31084 10508 31136
rect 10560 31124 10566 31136
rect 10781 31127 10839 31133
rect 10781 31124 10793 31127
rect 10560 31096 10793 31124
rect 10560 31084 10566 31096
rect 10781 31093 10793 31096
rect 10827 31093 10839 31127
rect 10781 31087 10839 31093
rect 10962 31084 10968 31136
rect 11020 31124 11026 31136
rect 12069 31127 12127 31133
rect 12069 31124 12081 31127
rect 11020 31096 12081 31124
rect 11020 31084 11026 31096
rect 12069 31093 12081 31096
rect 12115 31124 12127 31127
rect 12250 31124 12256 31136
rect 12115 31096 12256 31124
rect 12115 31093 12127 31096
rect 12069 31087 12127 31093
rect 12250 31084 12256 31096
rect 12308 31084 12314 31136
rect 12526 31084 12532 31136
rect 12584 31124 12590 31136
rect 12820 31124 12848 31164
rect 13630 31152 13636 31164
rect 13688 31152 13694 31204
rect 13924 31192 13952 31232
rect 14090 31220 14096 31232
rect 14148 31220 14154 31272
rect 17129 31263 17187 31269
rect 17129 31229 17141 31263
rect 17175 31260 17187 31263
rect 18248 31260 18276 31288
rect 17175 31232 18276 31260
rect 17175 31229 17187 31232
rect 17129 31223 17187 31229
rect 19794 31220 19800 31272
rect 19852 31260 19858 31272
rect 23216 31260 23244 31368
rect 23382 31288 23388 31340
rect 23440 31328 23446 31340
rect 23477 31331 23535 31337
rect 23477 31328 23489 31331
rect 23440 31300 23489 31328
rect 23440 31288 23446 31300
rect 23477 31297 23489 31300
rect 23523 31297 23535 31331
rect 23477 31291 23535 31297
rect 23934 31288 23940 31340
rect 23992 31328 23998 31340
rect 24121 31331 24179 31337
rect 24121 31328 24133 31331
rect 23992 31300 24133 31328
rect 23992 31288 23998 31300
rect 24121 31297 24133 31300
rect 24167 31328 24179 31331
rect 25130 31328 25136 31340
rect 24167 31300 25136 31328
rect 24167 31297 24179 31300
rect 24121 31291 24179 31297
rect 25130 31288 25136 31300
rect 25188 31288 25194 31340
rect 25225 31331 25283 31337
rect 25225 31297 25237 31331
rect 25271 31328 25283 31331
rect 25958 31328 25964 31340
rect 25271 31300 25964 31328
rect 25271 31297 25283 31300
rect 25225 31291 25283 31297
rect 25958 31288 25964 31300
rect 26016 31288 26022 31340
rect 26053 31331 26111 31337
rect 26053 31297 26065 31331
rect 26099 31328 26111 31331
rect 26142 31328 26148 31340
rect 26099 31300 26148 31328
rect 26099 31297 26111 31300
rect 26053 31291 26111 31297
rect 26142 31288 26148 31300
rect 26200 31288 26206 31340
rect 26973 31331 27031 31337
rect 26973 31297 26985 31331
rect 27019 31328 27031 31331
rect 27982 31328 27988 31340
rect 27019 31300 27988 31328
rect 27019 31297 27031 31300
rect 26973 31291 27031 31297
rect 27982 31288 27988 31300
rect 28040 31288 28046 31340
rect 28166 31288 28172 31340
rect 28224 31328 28230 31340
rect 28537 31331 28595 31337
rect 28537 31328 28549 31331
rect 28224 31300 28549 31328
rect 28224 31288 28230 31300
rect 28537 31297 28549 31300
rect 28583 31297 28595 31331
rect 28537 31291 28595 31297
rect 28626 31288 28632 31340
rect 28684 31328 28690 31340
rect 30190 31337 30196 31340
rect 28813 31331 28871 31337
rect 28813 31328 28825 31331
rect 28684 31300 28825 31328
rect 28684 31288 28690 31300
rect 28813 31297 28825 31300
rect 28859 31297 28871 31331
rect 29457 31331 29515 31337
rect 29457 31328 29469 31331
rect 28813 31291 28871 31297
rect 28920 31300 29469 31328
rect 19852 31232 23244 31260
rect 23293 31263 23351 31269
rect 19852 31220 19858 31232
rect 23293 31229 23305 31263
rect 23339 31260 23351 31263
rect 24026 31260 24032 31272
rect 23339 31232 24032 31260
rect 23339 31229 23351 31232
rect 23293 31223 23351 31229
rect 24026 31220 24032 31232
rect 24084 31220 24090 31272
rect 25501 31263 25559 31269
rect 25501 31229 25513 31263
rect 25547 31260 25559 31263
rect 25866 31260 25872 31272
rect 25547 31232 25872 31260
rect 25547 31229 25559 31232
rect 25501 31223 25559 31229
rect 25866 31220 25872 31232
rect 25924 31220 25930 31272
rect 27249 31263 27307 31269
rect 27249 31260 27261 31263
rect 26160 31232 27261 31260
rect 17221 31195 17279 31201
rect 13924 31164 17172 31192
rect 13078 31124 13084 31136
rect 12584 31096 12848 31124
rect 13039 31096 13084 31124
rect 12584 31084 12590 31096
rect 13078 31084 13084 31096
rect 13136 31084 13142 31136
rect 14458 31124 14464 31136
rect 14419 31096 14464 31124
rect 14458 31084 14464 31096
rect 14516 31084 14522 31136
rect 16666 31124 16672 31136
rect 16627 31096 16672 31124
rect 16666 31084 16672 31096
rect 16724 31084 16730 31136
rect 17034 31124 17040 31136
rect 16995 31096 17040 31124
rect 17034 31084 17040 31096
rect 17092 31084 17098 31136
rect 17144 31124 17172 31164
rect 17221 31161 17233 31195
rect 17267 31192 17279 31195
rect 25130 31192 25136 31204
rect 17267 31164 25136 31192
rect 17267 31161 17279 31164
rect 17221 31155 17279 31161
rect 25130 31152 25136 31164
rect 25188 31152 25194 31204
rect 25222 31152 25228 31204
rect 25280 31192 25286 31204
rect 25409 31195 25467 31201
rect 25409 31192 25421 31195
rect 25280 31164 25421 31192
rect 25280 31152 25286 31164
rect 25409 31161 25421 31164
rect 25455 31192 25467 31195
rect 26050 31192 26056 31204
rect 25455 31164 26056 31192
rect 25455 31161 25467 31164
rect 25409 31155 25467 31161
rect 26050 31152 26056 31164
rect 26108 31192 26114 31204
rect 26160 31192 26188 31232
rect 27249 31229 27261 31232
rect 27295 31260 27307 31263
rect 28721 31263 28779 31269
rect 28721 31260 28733 31263
rect 27295 31232 28733 31260
rect 27295 31229 27307 31232
rect 27249 31223 27307 31229
rect 28721 31229 28733 31232
rect 28767 31229 28779 31263
rect 28721 31223 28779 31229
rect 26108 31164 26188 31192
rect 26237 31195 26295 31201
rect 26108 31152 26114 31164
rect 26237 31161 26249 31195
rect 26283 31192 26295 31195
rect 26786 31192 26792 31204
rect 26283 31164 26792 31192
rect 26283 31161 26295 31164
rect 26237 31155 26295 31161
rect 26786 31152 26792 31164
rect 26844 31152 26850 31204
rect 22094 31124 22100 31136
rect 17144 31096 22100 31124
rect 22094 31084 22100 31096
rect 22152 31084 22158 31136
rect 22189 31127 22247 31133
rect 22189 31093 22201 31127
rect 22235 31124 22247 31127
rect 22462 31124 22468 31136
rect 22235 31096 22468 31124
rect 22235 31093 22247 31096
rect 22189 31087 22247 31093
rect 22462 31084 22468 31096
rect 22520 31084 22526 31136
rect 23658 31124 23664 31136
rect 23619 31096 23664 31124
rect 23658 31084 23664 31096
rect 23716 31084 23722 31136
rect 25038 31124 25044 31136
rect 24999 31096 25044 31124
rect 25038 31084 25044 31096
rect 25096 31084 25102 31136
rect 26602 31084 26608 31136
rect 26660 31124 26666 31136
rect 28920 31124 28948 31300
rect 29457 31297 29469 31300
rect 29503 31297 29515 31331
rect 30184 31328 30196 31337
rect 30151 31300 30196 31328
rect 29457 31291 29515 31297
rect 30184 31291 30196 31300
rect 30190 31288 30196 31291
rect 30248 31288 30254 31340
rect 29914 31260 29920 31272
rect 29875 31232 29920 31260
rect 29914 31220 29920 31232
rect 29972 31220 29978 31272
rect 26660 31096 28948 31124
rect 29273 31127 29331 31133
rect 26660 31084 26666 31096
rect 29273 31093 29285 31127
rect 29319 31124 29331 31127
rect 30650 31124 30656 31136
rect 29319 31096 30656 31124
rect 29319 31093 29331 31096
rect 29273 31087 29331 31093
rect 30650 31084 30656 31096
rect 30708 31084 30714 31136
rect 1104 31034 32016 31056
rect 1104 30982 2136 31034
rect 2188 30982 12440 31034
rect 12492 30982 22744 31034
rect 22796 30982 32016 31034
rect 1104 30960 32016 30982
rect 4246 30920 4252 30932
rect 4207 30892 4252 30920
rect 4246 30880 4252 30892
rect 4304 30880 4310 30932
rect 6454 30880 6460 30932
rect 6512 30920 6518 30932
rect 6733 30923 6791 30929
rect 6733 30920 6745 30923
rect 6512 30892 6745 30920
rect 6512 30880 6518 30892
rect 6733 30889 6745 30892
rect 6779 30889 6791 30923
rect 6733 30883 6791 30889
rect 7837 30923 7895 30929
rect 7837 30889 7849 30923
rect 7883 30920 7895 30923
rect 8202 30920 8208 30932
rect 7883 30892 8208 30920
rect 7883 30889 7895 30892
rect 7837 30883 7895 30889
rect 8202 30880 8208 30892
rect 8260 30880 8266 30932
rect 9217 30923 9275 30929
rect 9217 30889 9229 30923
rect 9263 30920 9275 30923
rect 9398 30920 9404 30932
rect 9263 30892 9404 30920
rect 9263 30889 9275 30892
rect 9217 30883 9275 30889
rect 9398 30880 9404 30892
rect 9456 30880 9462 30932
rect 10962 30920 10968 30932
rect 9784 30892 10968 30920
rect 2866 30852 2872 30864
rect 2779 30824 2872 30852
rect 2866 30812 2872 30824
rect 2924 30852 2930 30864
rect 6181 30855 6239 30861
rect 6181 30852 6193 30855
rect 2924 30824 6193 30852
rect 2924 30812 2930 30824
rect 6181 30821 6193 30824
rect 6227 30821 6239 30855
rect 6181 30815 6239 30821
rect 7742 30812 7748 30864
rect 7800 30852 7806 30864
rect 9784 30852 9812 30892
rect 10962 30880 10968 30892
rect 11020 30880 11026 30932
rect 11146 30920 11152 30932
rect 11107 30892 11152 30920
rect 11146 30880 11152 30892
rect 11204 30880 11210 30932
rect 11698 30880 11704 30932
rect 11756 30920 11762 30932
rect 11756 30892 12572 30920
rect 11756 30880 11762 30892
rect 12437 30855 12495 30861
rect 12437 30852 12449 30855
rect 7800 30824 9812 30852
rect 11900 30824 12449 30852
rect 7800 30812 7806 30824
rect 7926 30744 7932 30796
rect 7984 30784 7990 30796
rect 7984 30756 9904 30784
rect 7984 30744 7990 30756
rect 9876 30728 9904 30756
rect 1394 30676 1400 30728
rect 1452 30716 1458 30728
rect 1762 30725 1768 30728
rect 1489 30719 1547 30725
rect 1489 30716 1501 30719
rect 1452 30688 1501 30716
rect 1452 30676 1458 30688
rect 1489 30685 1501 30688
rect 1535 30685 1547 30719
rect 1756 30716 1768 30725
rect 1723 30688 1768 30716
rect 1489 30679 1547 30685
rect 1756 30679 1768 30688
rect 1762 30676 1768 30679
rect 1820 30676 1826 30728
rect 3694 30676 3700 30728
rect 3752 30716 3758 30728
rect 4433 30719 4491 30725
rect 4433 30716 4445 30719
rect 3752 30688 4445 30716
rect 3752 30676 3758 30688
rect 4433 30685 4445 30688
rect 4479 30685 4491 30719
rect 4433 30679 4491 30685
rect 4709 30719 4767 30725
rect 4709 30685 4721 30719
rect 4755 30685 4767 30719
rect 4890 30716 4896 30728
rect 4851 30688 4896 30716
rect 4709 30679 4767 30685
rect 4154 30608 4160 30660
rect 4212 30648 4218 30660
rect 4724 30648 4752 30679
rect 4890 30676 4896 30688
rect 4948 30676 4954 30728
rect 5721 30719 5779 30725
rect 5721 30685 5733 30719
rect 5767 30716 5779 30719
rect 5902 30716 5908 30728
rect 5767 30688 5908 30716
rect 5767 30685 5779 30688
rect 5721 30679 5779 30685
rect 5902 30676 5908 30688
rect 5960 30676 5966 30728
rect 7377 30719 7435 30725
rect 7377 30685 7389 30719
rect 7423 30716 7435 30719
rect 7558 30716 7564 30728
rect 7423 30688 7564 30716
rect 7423 30685 7435 30688
rect 7377 30679 7435 30685
rect 7558 30676 7564 30688
rect 7616 30676 7622 30728
rect 8021 30719 8079 30725
rect 8021 30685 8033 30719
rect 8067 30685 8079 30719
rect 8021 30679 8079 30685
rect 4212 30620 4752 30648
rect 6457 30651 6515 30657
rect 4212 30608 4218 30620
rect 6457 30617 6469 30651
rect 6503 30648 6515 30651
rect 7006 30648 7012 30660
rect 6503 30620 7012 30648
rect 6503 30617 6515 30620
rect 6457 30611 6515 30617
rect 7006 30608 7012 30620
rect 7064 30608 7070 30660
rect 8036 30648 8064 30679
rect 8110 30676 8116 30728
rect 8168 30716 8174 30728
rect 8294 30716 8300 30728
rect 8168 30688 8213 30716
rect 8255 30688 8300 30716
rect 8168 30676 8174 30688
rect 8294 30676 8300 30688
rect 8352 30676 8358 30728
rect 8389 30719 8447 30725
rect 8389 30685 8401 30719
rect 8435 30716 8447 30719
rect 8846 30716 8852 30728
rect 8435 30688 8852 30716
rect 8435 30685 8447 30688
rect 8389 30679 8447 30685
rect 8846 30676 8852 30688
rect 8904 30716 8910 30728
rect 9125 30719 9183 30725
rect 9125 30716 9137 30719
rect 8904 30688 9137 30716
rect 8904 30676 8910 30688
rect 9125 30685 9137 30688
rect 9171 30685 9183 30719
rect 9766 30716 9772 30728
rect 9727 30688 9772 30716
rect 9125 30679 9183 30685
rect 9766 30676 9772 30688
rect 9824 30676 9830 30728
rect 9858 30676 9864 30728
rect 9916 30676 9922 30728
rect 10036 30719 10094 30725
rect 10036 30685 10048 30719
rect 10082 30716 10094 30719
rect 10410 30716 10416 30728
rect 10082 30688 10416 30716
rect 10082 30685 10094 30688
rect 10036 30679 10094 30685
rect 10410 30676 10416 30688
rect 10468 30676 10474 30728
rect 11900 30725 11928 30824
rect 12437 30821 12449 30824
rect 12483 30821 12495 30855
rect 12544 30852 12572 30892
rect 12710 30880 12716 30932
rect 12768 30920 12774 30932
rect 12897 30923 12955 30929
rect 12897 30920 12909 30923
rect 12768 30892 12909 30920
rect 12768 30880 12774 30892
rect 12897 30889 12909 30892
rect 12943 30889 12955 30923
rect 14090 30920 14096 30932
rect 14051 30892 14096 30920
rect 12897 30883 12955 30889
rect 14090 30880 14096 30892
rect 14148 30880 14154 30932
rect 15930 30880 15936 30932
rect 15988 30920 15994 30932
rect 16577 30923 16635 30929
rect 16577 30920 16589 30923
rect 15988 30892 16589 30920
rect 15988 30880 15994 30892
rect 16577 30889 16589 30892
rect 16623 30889 16635 30923
rect 16577 30883 16635 30889
rect 17310 30880 17316 30932
rect 17368 30920 17374 30932
rect 17770 30920 17776 30932
rect 17368 30892 17776 30920
rect 17368 30880 17374 30892
rect 17770 30880 17776 30892
rect 17828 30880 17834 30932
rect 19245 30923 19303 30929
rect 19245 30889 19257 30923
rect 19291 30920 19303 30923
rect 22094 30920 22100 30932
rect 19291 30892 22100 30920
rect 19291 30889 19303 30892
rect 19245 30883 19303 30889
rect 22094 30880 22100 30892
rect 22152 30880 22158 30932
rect 23566 30920 23572 30932
rect 22204 30892 23572 30920
rect 13449 30855 13507 30861
rect 13449 30852 13461 30855
rect 12544 30824 13461 30852
rect 12437 30815 12495 30821
rect 13449 30821 13461 30824
rect 13495 30852 13507 30855
rect 14274 30852 14280 30864
rect 13495 30824 14280 30852
rect 13495 30821 13507 30824
rect 13449 30815 13507 30821
rect 14274 30812 14280 30824
rect 14332 30812 14338 30864
rect 14553 30855 14611 30861
rect 14553 30821 14565 30855
rect 14599 30852 14611 30855
rect 15102 30852 15108 30864
rect 14599 30824 15108 30852
rect 14599 30821 14611 30824
rect 14553 30815 14611 30821
rect 15102 30812 15108 30824
rect 15160 30812 15166 30864
rect 19426 30812 19432 30864
rect 19484 30852 19490 30864
rect 19978 30852 19984 30864
rect 19484 30824 19984 30852
rect 19484 30812 19490 30824
rect 19978 30812 19984 30824
rect 20036 30812 20042 30864
rect 21726 30852 21732 30864
rect 21687 30824 21732 30852
rect 21726 30812 21732 30824
rect 21784 30812 21790 30864
rect 22204 30852 22232 30892
rect 23566 30880 23572 30892
rect 23624 30880 23630 30932
rect 25958 30880 25964 30932
rect 26016 30920 26022 30932
rect 26237 30923 26295 30929
rect 26237 30920 26249 30923
rect 26016 30892 26249 30920
rect 26016 30880 26022 30892
rect 26237 30889 26249 30892
rect 26283 30889 26295 30923
rect 26237 30883 26295 30889
rect 30282 30880 30288 30932
rect 30340 30920 30346 30932
rect 30653 30923 30711 30929
rect 30653 30920 30665 30923
rect 30340 30892 30665 30920
rect 30340 30880 30346 30892
rect 30653 30889 30665 30892
rect 30699 30889 30711 30923
rect 30653 30883 30711 30889
rect 21928 30824 22232 30852
rect 11977 30787 12035 30793
rect 11977 30753 11989 30787
rect 12023 30784 12035 30787
rect 14737 30787 14795 30793
rect 14737 30784 14749 30787
rect 12023 30756 14320 30784
rect 14647 30756 14749 30784
rect 12023 30753 12035 30756
rect 11977 30747 12035 30753
rect 11885 30719 11943 30725
rect 11885 30685 11897 30719
rect 11931 30685 11943 30719
rect 11885 30679 11943 30685
rect 12069 30719 12127 30725
rect 12069 30685 12081 30719
rect 12115 30716 12127 30719
rect 12158 30716 12164 30728
rect 12115 30688 12164 30716
rect 12115 30685 12127 30688
rect 12069 30679 12127 30685
rect 12158 30676 12164 30688
rect 12216 30676 12222 30728
rect 12713 30719 12771 30725
rect 12713 30685 12725 30719
rect 12759 30716 12771 30719
rect 13078 30716 13084 30728
rect 12759 30688 13084 30716
rect 12759 30685 12771 30688
rect 12713 30679 12771 30685
rect 13078 30676 13084 30688
rect 13136 30676 13142 30728
rect 14292 30725 14320 30756
rect 13357 30719 13415 30725
rect 13357 30685 13369 30719
rect 13403 30685 13415 30719
rect 13357 30679 13415 30685
rect 14277 30719 14335 30725
rect 14277 30685 14289 30719
rect 14323 30685 14335 30719
rect 14277 30679 14335 30685
rect 8938 30648 8944 30660
rect 8036 30620 8944 30648
rect 8938 30608 8944 30620
rect 8996 30608 9002 30660
rect 12526 30648 12532 30660
rect 12487 30620 12532 30648
rect 12526 30608 12532 30620
rect 12584 30608 12590 30660
rect 12618 30608 12624 30660
rect 12676 30648 12682 30660
rect 13372 30648 13400 30679
rect 14366 30676 14372 30728
rect 14424 30716 14430 30728
rect 14660 30725 14688 30756
rect 14737 30753 14749 30756
rect 14783 30784 14795 30787
rect 14918 30784 14924 30796
rect 14783 30756 14924 30784
rect 14783 30753 14795 30756
rect 14737 30747 14795 30753
rect 14918 30744 14924 30756
rect 14976 30744 14982 30796
rect 19242 30784 19248 30796
rect 18064 30756 19248 30784
rect 18064 30728 18092 30756
rect 19242 30744 19248 30756
rect 19300 30784 19306 30796
rect 20349 30787 20407 30793
rect 20349 30784 20361 30787
rect 19300 30756 20361 30784
rect 19300 30744 19306 30756
rect 20349 30753 20361 30756
rect 20395 30753 20407 30787
rect 20349 30747 20407 30753
rect 14645 30719 14703 30725
rect 14424 30688 14469 30716
rect 14424 30676 14430 30688
rect 14645 30685 14657 30719
rect 14691 30685 14703 30719
rect 15194 30716 15200 30728
rect 15155 30688 15200 30716
rect 14645 30679 14703 30685
rect 15194 30676 15200 30688
rect 15252 30676 15258 30728
rect 15470 30725 15476 30728
rect 15464 30716 15476 30725
rect 15431 30688 15476 30716
rect 15464 30679 15476 30688
rect 15470 30676 15476 30679
rect 15528 30676 15534 30728
rect 17037 30719 17095 30725
rect 17037 30685 17049 30719
rect 17083 30716 17095 30719
rect 18046 30716 18052 30728
rect 17083 30688 18052 30716
rect 17083 30685 17095 30688
rect 17037 30679 17095 30685
rect 18046 30676 18052 30688
rect 18104 30676 18110 30728
rect 19150 30676 19156 30728
rect 19208 30716 19214 30728
rect 19429 30719 19487 30725
rect 19429 30716 19441 30719
rect 19208 30688 19441 30716
rect 19208 30676 19214 30688
rect 19429 30685 19441 30688
rect 19475 30685 19487 30719
rect 19429 30679 19487 30685
rect 19705 30719 19763 30725
rect 19705 30685 19717 30719
rect 19751 30685 19763 30719
rect 19705 30679 19763 30685
rect 19889 30719 19947 30725
rect 19889 30685 19901 30719
rect 19935 30716 19947 30719
rect 21928 30716 21956 30824
rect 22186 30784 22192 30796
rect 22147 30756 22192 30784
rect 22186 30744 22192 30756
rect 22244 30744 22250 30796
rect 26326 30744 26332 30796
rect 26384 30784 26390 30796
rect 29549 30787 29607 30793
rect 29549 30784 29561 30787
rect 26384 30756 26740 30784
rect 26384 30744 26390 30756
rect 24397 30719 24455 30725
rect 24397 30716 24409 30719
rect 19935 30688 21956 30716
rect 22066 30688 24409 30716
rect 19935 30685 19947 30688
rect 19889 30679 19947 30685
rect 12676 30620 13400 30648
rect 12676 30608 12682 30620
rect 16666 30608 16672 30660
rect 16724 30648 16730 30660
rect 17282 30651 17340 30657
rect 17282 30648 17294 30651
rect 16724 30620 17294 30648
rect 16724 30608 16730 30620
rect 17282 30617 17294 30620
rect 17328 30617 17340 30651
rect 17282 30611 17340 30617
rect 19242 30608 19248 30660
rect 19300 30648 19306 30660
rect 19720 30648 19748 30679
rect 20622 30657 20628 30660
rect 19300 30620 19748 30648
rect 19300 30608 19306 30620
rect 20616 30611 20628 30657
rect 20680 30648 20686 30660
rect 22066 30648 22094 30688
rect 24397 30685 24409 30688
rect 24443 30685 24455 30719
rect 24397 30679 24455 30685
rect 24664 30719 24722 30725
rect 24664 30685 24676 30719
rect 24710 30716 24722 30719
rect 25038 30716 25044 30728
rect 24710 30688 25044 30716
rect 24710 30685 24722 30688
rect 24664 30679 24722 30685
rect 25038 30676 25044 30688
rect 25096 30676 25102 30728
rect 25130 30676 25136 30728
rect 25188 30716 25194 30728
rect 26234 30716 26240 30728
rect 25188 30688 26240 30716
rect 25188 30676 25194 30688
rect 26234 30676 26240 30688
rect 26292 30676 26298 30728
rect 26418 30716 26424 30728
rect 26379 30688 26424 30716
rect 26418 30676 26424 30688
rect 26476 30676 26482 30728
rect 26712 30725 26740 30756
rect 28736 30756 29561 30784
rect 26697 30719 26755 30725
rect 26697 30685 26709 30719
rect 26743 30685 26755 30719
rect 26697 30679 26755 30685
rect 26881 30719 26939 30725
rect 26881 30685 26893 30719
rect 26927 30685 26939 30719
rect 26881 30679 26939 30685
rect 27893 30719 27951 30725
rect 27893 30685 27905 30719
rect 27939 30716 27951 30719
rect 27982 30716 27988 30728
rect 27939 30688 27988 30716
rect 27939 30685 27951 30688
rect 27893 30679 27951 30685
rect 20680 30620 20716 30648
rect 21836 30620 22094 30648
rect 20622 30608 20628 30611
rect 20680 30608 20686 30620
rect 21836 30592 21864 30620
rect 22186 30608 22192 30660
rect 22244 30648 22250 30660
rect 22434 30651 22492 30657
rect 22434 30648 22446 30651
rect 22244 30620 22446 30648
rect 22244 30608 22250 30620
rect 22434 30617 22446 30620
rect 22480 30617 22492 30651
rect 22434 30611 22492 30617
rect 5537 30583 5595 30589
rect 5537 30549 5549 30583
rect 5583 30580 5595 30583
rect 6086 30580 6092 30592
rect 5583 30552 6092 30580
rect 5583 30549 5595 30552
rect 5537 30543 5595 30549
rect 6086 30540 6092 30552
rect 6144 30540 6150 30592
rect 6362 30580 6368 30592
rect 6323 30552 6368 30580
rect 6362 30540 6368 30552
rect 6420 30540 6426 30592
rect 6549 30583 6607 30589
rect 6549 30549 6561 30583
rect 6595 30580 6607 30583
rect 6730 30580 6736 30592
rect 6595 30552 6736 30580
rect 6595 30549 6607 30552
rect 6549 30543 6607 30549
rect 6730 30540 6736 30552
rect 6788 30540 6794 30592
rect 7190 30580 7196 30592
rect 7151 30552 7196 30580
rect 7190 30540 7196 30552
rect 7248 30540 7254 30592
rect 7374 30540 7380 30592
rect 7432 30580 7438 30592
rect 12066 30580 12072 30592
rect 7432 30552 12072 30580
rect 7432 30540 7438 30552
rect 12066 30540 12072 30552
rect 12124 30540 12130 30592
rect 12437 30583 12495 30589
rect 12437 30549 12449 30583
rect 12483 30580 12495 30583
rect 13906 30580 13912 30592
rect 12483 30552 13912 30580
rect 12483 30549 12495 30552
rect 12437 30543 12495 30549
rect 13906 30540 13912 30552
rect 13964 30580 13970 30592
rect 14737 30583 14795 30589
rect 14737 30580 14749 30583
rect 13964 30552 14749 30580
rect 13964 30540 13970 30552
rect 14737 30549 14749 30552
rect 14783 30549 14795 30583
rect 14737 30543 14795 30549
rect 16942 30540 16948 30592
rect 17000 30580 17006 30592
rect 17402 30580 17408 30592
rect 17000 30552 17408 30580
rect 17000 30540 17006 30552
rect 17402 30540 17408 30552
rect 17460 30540 17466 30592
rect 18138 30540 18144 30592
rect 18196 30580 18202 30592
rect 18417 30583 18475 30589
rect 18417 30580 18429 30583
rect 18196 30552 18429 30580
rect 18196 30540 18202 30552
rect 18417 30549 18429 30552
rect 18463 30549 18475 30583
rect 18417 30543 18475 30549
rect 21818 30540 21824 30592
rect 21876 30540 21882 30592
rect 25314 30540 25320 30592
rect 25372 30580 25378 30592
rect 25777 30583 25835 30589
rect 25777 30580 25789 30583
rect 25372 30552 25789 30580
rect 25372 30540 25378 30552
rect 25777 30549 25789 30552
rect 25823 30580 25835 30583
rect 26896 30580 26924 30679
rect 27982 30676 27988 30688
rect 28040 30676 28046 30728
rect 28736 30725 28764 30756
rect 29549 30753 29561 30756
rect 29595 30753 29607 30787
rect 30742 30784 30748 30796
rect 29549 30747 29607 30753
rect 30024 30756 30748 30784
rect 28721 30719 28779 30725
rect 28721 30685 28733 30719
rect 28767 30685 28779 30719
rect 28902 30716 28908 30728
rect 28863 30688 28908 30716
rect 28721 30679 28779 30685
rect 28902 30676 28908 30688
rect 28960 30676 28966 30728
rect 28994 30676 29000 30728
rect 29052 30716 29058 30728
rect 30024 30725 30052 30756
rect 30742 30744 30748 30756
rect 30800 30784 30806 30796
rect 31202 30784 31208 30796
rect 30800 30756 31208 30784
rect 30800 30744 30806 30756
rect 29733 30719 29791 30725
rect 29052 30688 29097 30716
rect 29052 30676 29058 30688
rect 29733 30685 29745 30719
rect 29779 30685 29791 30719
rect 29733 30679 29791 30685
rect 30009 30719 30067 30725
rect 30009 30685 30021 30719
rect 30055 30685 30067 30719
rect 30009 30679 30067 30685
rect 28077 30651 28135 30657
rect 28077 30617 28089 30651
rect 28123 30648 28135 30651
rect 28920 30648 28948 30676
rect 28123 30620 28948 30648
rect 29748 30648 29776 30679
rect 30098 30676 30104 30728
rect 30156 30716 30162 30728
rect 31128 30725 31156 30756
rect 31202 30744 31208 30756
rect 31260 30744 31266 30796
rect 30193 30719 30251 30725
rect 30193 30716 30205 30719
rect 30156 30688 30205 30716
rect 30156 30676 30162 30688
rect 30193 30685 30205 30688
rect 30239 30685 30251 30719
rect 30837 30719 30895 30725
rect 30837 30716 30849 30719
rect 30193 30679 30251 30685
rect 30668 30688 30849 30716
rect 30668 30660 30696 30688
rect 30837 30685 30849 30688
rect 30883 30685 30895 30719
rect 30837 30679 30895 30685
rect 31113 30719 31171 30725
rect 31113 30685 31125 30719
rect 31159 30685 31171 30719
rect 31294 30716 31300 30728
rect 31255 30688 31300 30716
rect 31113 30679 31171 30685
rect 31294 30676 31300 30688
rect 31352 30676 31358 30728
rect 30650 30648 30656 30660
rect 29748 30620 30656 30648
rect 28123 30617 28135 30620
rect 28077 30611 28135 30617
rect 30650 30608 30656 30620
rect 30708 30608 30714 30660
rect 25823 30552 26924 30580
rect 28537 30583 28595 30589
rect 25823 30549 25835 30552
rect 25777 30543 25835 30549
rect 28537 30549 28549 30583
rect 28583 30580 28595 30583
rect 30006 30580 30012 30592
rect 28583 30552 30012 30580
rect 28583 30549 28595 30552
rect 28537 30543 28595 30549
rect 30006 30540 30012 30552
rect 30064 30540 30070 30592
rect 1104 30490 32016 30512
rect 1104 30438 7288 30490
rect 7340 30438 17592 30490
rect 17644 30438 27896 30490
rect 27948 30438 32016 30490
rect 1104 30416 32016 30438
rect 1857 30379 1915 30385
rect 1857 30345 1869 30379
rect 1903 30376 1915 30379
rect 2590 30376 2596 30388
rect 1903 30348 2596 30376
rect 1903 30345 1915 30348
rect 1857 30339 1915 30345
rect 2590 30336 2596 30348
rect 2648 30336 2654 30388
rect 8478 30376 8484 30388
rect 8220 30348 8484 30376
rect 3694 30308 3700 30320
rect 2056 30280 3700 30308
rect 2056 30249 2084 30280
rect 2041 30243 2099 30249
rect 2041 30209 2053 30243
rect 2087 30209 2099 30243
rect 2041 30203 2099 30209
rect 2317 30243 2375 30249
rect 2317 30209 2329 30243
rect 2363 30209 2375 30243
rect 2317 30203 2375 30209
rect 2501 30243 2559 30249
rect 2501 30209 2513 30243
rect 2547 30240 2559 30243
rect 2866 30240 2872 30252
rect 2547 30212 2872 30240
rect 2547 30209 2559 30212
rect 2501 30203 2559 30209
rect 2332 30172 2360 30203
rect 2866 30200 2872 30212
rect 2924 30200 2930 30252
rect 3160 30249 3188 30280
rect 3694 30268 3700 30280
rect 3752 30268 3758 30320
rect 4338 30268 4344 30320
rect 4396 30308 4402 30320
rect 4494 30311 4552 30317
rect 4494 30308 4506 30311
rect 4396 30280 4506 30308
rect 4396 30268 4402 30280
rect 4494 30277 4506 30280
rect 4540 30277 4552 30311
rect 4494 30271 4552 30277
rect 6638 30268 6644 30320
rect 6696 30308 6702 30320
rect 8220 30308 8248 30348
rect 8478 30336 8484 30348
rect 8536 30336 8542 30388
rect 8573 30379 8631 30385
rect 8573 30345 8585 30379
rect 8619 30376 8631 30379
rect 8662 30376 8668 30388
rect 8619 30348 8668 30376
rect 8619 30345 8631 30348
rect 8573 30339 8631 30345
rect 8662 30336 8668 30348
rect 8720 30336 8726 30388
rect 9309 30379 9367 30385
rect 9309 30345 9321 30379
rect 9355 30376 9367 30379
rect 9674 30376 9680 30388
rect 9355 30348 9680 30376
rect 9355 30345 9367 30348
rect 9309 30339 9367 30345
rect 9674 30336 9680 30348
rect 9732 30336 9738 30388
rect 12526 30336 12532 30388
rect 12584 30376 12590 30388
rect 12802 30376 12808 30388
rect 12584 30348 12808 30376
rect 12584 30336 12590 30348
rect 12802 30336 12808 30348
rect 12860 30336 12866 30388
rect 12894 30336 12900 30388
rect 12952 30376 12958 30388
rect 14550 30376 14556 30388
rect 12952 30348 14556 30376
rect 12952 30336 12958 30348
rect 14550 30336 14556 30348
rect 14608 30376 14614 30388
rect 14829 30379 14887 30385
rect 14829 30376 14841 30379
rect 14608 30348 14841 30376
rect 14608 30336 14614 30348
rect 14829 30345 14841 30348
rect 14875 30376 14887 30379
rect 15194 30376 15200 30388
rect 14875 30348 15200 30376
rect 14875 30345 14887 30348
rect 14829 30339 14887 30345
rect 15194 30336 15200 30348
rect 15252 30336 15258 30388
rect 16850 30336 16856 30388
rect 16908 30376 16914 30388
rect 17497 30379 17555 30385
rect 17497 30376 17509 30379
rect 16908 30348 17509 30376
rect 16908 30336 16914 30348
rect 17497 30345 17509 30348
rect 17543 30345 17555 30379
rect 18230 30376 18236 30388
rect 17497 30339 17555 30345
rect 17696 30348 18236 30376
rect 6696 30280 8248 30308
rect 6696 30268 6702 30280
rect 3145 30243 3203 30249
rect 3145 30209 3157 30243
rect 3191 30209 3203 30243
rect 3145 30203 3203 30209
rect 3421 30243 3479 30249
rect 3421 30209 3433 30243
rect 3467 30209 3479 30243
rect 3602 30240 3608 30252
rect 3563 30212 3608 30240
rect 3421 30203 3479 30209
rect 3436 30172 3464 30203
rect 3602 30200 3608 30212
rect 3660 30200 3666 30252
rect 6730 30200 6736 30252
rect 6788 30240 6794 30252
rect 7208 30249 7236 30280
rect 8294 30268 8300 30320
rect 8352 30308 8358 30320
rect 11517 30311 11575 30317
rect 11517 30308 11529 30311
rect 8352 30280 11529 30308
rect 8352 30268 8358 30280
rect 11517 30277 11529 30280
rect 11563 30277 11575 30311
rect 11517 30271 11575 30277
rect 12250 30268 12256 30320
rect 12308 30308 12314 30320
rect 13541 30311 13599 30317
rect 13541 30308 13553 30311
rect 12308 30280 13553 30308
rect 12308 30268 12314 30280
rect 13541 30277 13553 30280
rect 13587 30277 13599 30311
rect 13541 30271 13599 30277
rect 14918 30268 14924 30320
rect 14976 30308 14982 30320
rect 16761 30311 16819 30317
rect 16761 30308 16773 30311
rect 14976 30280 16773 30308
rect 14976 30268 14982 30280
rect 16761 30277 16773 30280
rect 16807 30308 16819 30311
rect 17405 30311 17463 30317
rect 17405 30308 17417 30311
rect 16807 30280 17417 30308
rect 16807 30277 16819 30280
rect 16761 30271 16819 30277
rect 17405 30277 17417 30280
rect 17451 30277 17463 30311
rect 17405 30271 17463 30277
rect 7009 30243 7067 30249
rect 7009 30240 7021 30243
rect 6788 30212 7021 30240
rect 6788 30200 6794 30212
rect 7009 30209 7021 30212
rect 7055 30209 7067 30243
rect 7009 30203 7067 30209
rect 7193 30243 7251 30249
rect 7193 30209 7205 30243
rect 7239 30209 7251 30243
rect 7374 30240 7380 30252
rect 7335 30212 7380 30240
rect 7193 30203 7251 30209
rect 7374 30200 7380 30212
rect 7432 30200 7438 30252
rect 8202 30200 8208 30252
rect 8260 30240 8266 30252
rect 8389 30243 8447 30249
rect 8389 30240 8401 30243
rect 8260 30212 8401 30240
rect 8260 30200 8266 30212
rect 8389 30209 8401 30212
rect 8435 30209 8447 30243
rect 8389 30203 8447 30209
rect 8478 30200 8484 30252
rect 8536 30240 8542 30252
rect 9490 30240 9496 30252
rect 8536 30212 8581 30240
rect 9451 30212 9496 30240
rect 8536 30200 8542 30212
rect 9490 30200 9496 30212
rect 9548 30200 9554 30252
rect 9582 30200 9588 30252
rect 9640 30240 9646 30252
rect 11701 30243 11759 30249
rect 11701 30240 11713 30243
rect 9640 30212 11713 30240
rect 9640 30200 9646 30212
rect 11701 30209 11713 30212
rect 11747 30209 11759 30243
rect 12526 30240 12532 30252
rect 12487 30212 12532 30240
rect 11701 30203 11759 30209
rect 12526 30200 12532 30212
rect 12584 30200 12590 30252
rect 12713 30243 12771 30249
rect 12713 30209 12725 30243
rect 12759 30240 12771 30243
rect 12986 30240 12992 30252
rect 12759 30212 12992 30240
rect 12759 30209 12771 30212
rect 12713 30203 12771 30209
rect 4246 30172 4252 30184
rect 2332 30144 3556 30172
rect 4207 30144 4252 30172
rect 3528 30104 3556 30144
rect 4246 30132 4252 30144
rect 4304 30132 4310 30184
rect 7285 30175 7343 30181
rect 7285 30141 7297 30175
rect 7331 30172 7343 30175
rect 7466 30172 7472 30184
rect 7331 30144 7472 30172
rect 7331 30141 7343 30144
rect 7285 30135 7343 30141
rect 7466 30132 7472 30144
rect 7524 30172 7530 30184
rect 9600 30172 9628 30200
rect 7524 30144 9628 30172
rect 7524 30132 7530 30144
rect 9858 30132 9864 30184
rect 9916 30172 9922 30184
rect 9953 30175 10011 30181
rect 9953 30172 9965 30175
rect 9916 30144 9965 30172
rect 9916 30132 9922 30144
rect 9953 30141 9965 30144
rect 9999 30141 10011 30175
rect 9953 30135 10011 30141
rect 10229 30175 10287 30181
rect 10229 30141 10241 30175
rect 10275 30172 10287 30175
rect 10502 30172 10508 30184
rect 10275 30144 10508 30172
rect 10275 30141 10287 30144
rect 10229 30135 10287 30141
rect 10502 30132 10508 30144
rect 10560 30132 10566 30184
rect 11974 30172 11980 30184
rect 11935 30144 11980 30172
rect 11974 30132 11980 30144
rect 12032 30132 12038 30184
rect 12066 30132 12072 30184
rect 12124 30172 12130 30184
rect 12728 30172 12756 30203
rect 12986 30200 12992 30212
rect 13044 30200 13050 30252
rect 15470 30240 15476 30252
rect 13648 30212 15476 30240
rect 12124 30144 12756 30172
rect 12124 30132 12130 30144
rect 4154 30104 4160 30116
rect 3528 30076 4160 30104
rect 4154 30064 4160 30076
rect 4212 30064 4218 30116
rect 8205 30107 8263 30113
rect 8205 30073 8217 30107
rect 8251 30104 8263 30107
rect 8251 30076 8423 30104
rect 8251 30073 8263 30076
rect 8205 30067 8263 30073
rect 8395 30048 8423 30076
rect 9490 30064 9496 30116
rect 9548 30104 9554 30116
rect 13648 30104 13676 30212
rect 15470 30200 15476 30212
rect 15528 30240 15534 30252
rect 15841 30243 15899 30249
rect 15841 30240 15853 30243
rect 15528 30212 15853 30240
rect 15528 30200 15534 30212
rect 15841 30209 15853 30212
rect 15887 30209 15899 30243
rect 15841 30203 15899 30209
rect 16574 30200 16580 30252
rect 16632 30240 16638 30252
rect 17494 30240 17500 30252
rect 16632 30212 17500 30240
rect 16632 30200 16638 30212
rect 17494 30200 17500 30212
rect 17552 30200 17558 30252
rect 17696 30249 17724 30348
rect 18230 30336 18236 30348
rect 18288 30376 18294 30388
rect 19150 30376 19156 30388
rect 18288 30348 19156 30376
rect 18288 30336 18294 30348
rect 19150 30336 19156 30348
rect 19208 30336 19214 30388
rect 19518 30336 19524 30388
rect 19576 30376 19582 30388
rect 20073 30379 20131 30385
rect 20073 30376 20085 30379
rect 19576 30348 20085 30376
rect 19576 30336 19582 30348
rect 20073 30345 20085 30348
rect 20119 30376 20131 30379
rect 20438 30376 20444 30388
rect 20119 30348 20444 30376
rect 20119 30345 20131 30348
rect 20073 30339 20131 30345
rect 20438 30336 20444 30348
rect 20496 30336 20502 30388
rect 20622 30376 20628 30388
rect 20583 30348 20628 30376
rect 20622 30336 20628 30348
rect 20680 30336 20686 30388
rect 22097 30379 22155 30385
rect 22097 30345 22109 30379
rect 22143 30376 22155 30379
rect 22186 30376 22192 30388
rect 22143 30348 22192 30376
rect 22143 30345 22155 30348
rect 22097 30339 22155 30345
rect 22186 30336 22192 30348
rect 22244 30336 22250 30388
rect 26418 30376 26424 30388
rect 26252 30348 26424 30376
rect 19242 30308 19248 30320
rect 17972 30280 19248 30308
rect 17972 30252 18000 30280
rect 17681 30243 17739 30249
rect 17681 30209 17693 30243
rect 17727 30209 17739 30243
rect 17954 30240 17960 30252
rect 17915 30212 17960 30240
rect 17681 30203 17739 30209
rect 17954 30200 17960 30212
rect 18012 30200 18018 30252
rect 18138 30240 18144 30252
rect 18099 30212 18144 30240
rect 18138 30200 18144 30212
rect 18196 30200 18202 30252
rect 18506 30200 18512 30252
rect 18564 30240 18570 30252
rect 18892 30249 18920 30280
rect 19242 30268 19248 30280
rect 19300 30268 19306 30320
rect 19334 30268 19340 30320
rect 19392 30308 19398 30320
rect 23109 30311 23167 30317
rect 23109 30308 23121 30311
rect 19392 30280 23121 30308
rect 19392 30268 19398 30280
rect 23109 30277 23121 30280
rect 23155 30277 23167 30311
rect 26252 30308 26280 30348
rect 26418 30336 26424 30348
rect 26476 30336 26482 30388
rect 23109 30271 23167 30277
rect 25976 30280 26280 30308
rect 26344 30280 27292 30308
rect 18877 30243 18935 30249
rect 18564 30212 18736 30240
rect 18564 30200 18570 30212
rect 16114 30132 16120 30184
rect 16172 30172 16178 30184
rect 17512 30172 17540 30200
rect 18233 30175 18291 30181
rect 18233 30172 18245 30175
rect 16172 30144 17448 30172
rect 17512 30144 18245 30172
rect 16172 30132 16178 30144
rect 9548 30076 13676 30104
rect 9548 30064 9554 30076
rect 14366 30064 14372 30116
rect 14424 30104 14430 30116
rect 15010 30104 15016 30116
rect 14424 30076 15016 30104
rect 14424 30064 14430 30076
rect 15010 30064 15016 30076
rect 15068 30104 15074 30116
rect 16945 30107 17003 30113
rect 16945 30104 16957 30107
rect 15068 30076 16957 30104
rect 15068 30064 15074 30076
rect 16945 30073 16957 30076
rect 16991 30073 17003 30107
rect 17420 30104 17448 30144
rect 18233 30141 18245 30144
rect 18279 30141 18291 30175
rect 18598 30172 18604 30184
rect 18233 30135 18291 30141
rect 18340 30144 18604 30172
rect 18340 30104 18368 30144
rect 18598 30132 18604 30144
rect 18656 30132 18662 30184
rect 18708 30172 18736 30212
rect 18877 30209 18889 30243
rect 18923 30209 18935 30243
rect 18877 30203 18935 30209
rect 19797 30243 19855 30249
rect 19797 30209 19809 30243
rect 19843 30240 19855 30243
rect 19889 30243 19947 30249
rect 19889 30240 19901 30243
rect 19843 30212 19901 30240
rect 19843 30209 19855 30212
rect 19797 30203 19855 30209
rect 19889 30209 19901 30212
rect 19935 30209 19947 30243
rect 20806 30240 20812 30252
rect 20767 30212 20812 30240
rect 19889 30203 19947 30209
rect 20806 30200 20812 30212
rect 20864 30200 20870 30252
rect 22094 30200 22100 30252
rect 22152 30240 22158 30252
rect 22281 30243 22339 30249
rect 22281 30240 22293 30243
rect 22152 30212 22293 30240
rect 22152 30200 22158 30212
rect 22281 30209 22293 30212
rect 22327 30209 22339 30243
rect 22462 30240 22468 30252
rect 22423 30212 22468 30240
rect 22281 30203 22339 30209
rect 22462 30200 22468 30212
rect 22520 30200 22526 30252
rect 23017 30243 23075 30249
rect 23017 30209 23029 30243
rect 23063 30209 23075 30243
rect 23658 30240 23664 30252
rect 23619 30212 23664 30240
rect 23017 30203 23075 30209
rect 20990 30172 20996 30184
rect 18708 30144 20996 30172
rect 20990 30132 20996 30144
rect 21048 30132 21054 30184
rect 21085 30175 21143 30181
rect 21085 30141 21097 30175
rect 21131 30172 21143 30175
rect 22557 30175 22615 30181
rect 21131 30144 22140 30172
rect 21131 30141 21143 30144
rect 21085 30135 21143 30141
rect 22112 30116 22140 30144
rect 22557 30141 22569 30175
rect 22603 30172 22615 30175
rect 22830 30172 22836 30184
rect 22603 30144 22836 30172
rect 22603 30141 22615 30144
rect 22557 30135 22615 30141
rect 22830 30132 22836 30144
rect 22888 30132 22894 30184
rect 17420 30076 18368 30104
rect 18417 30107 18475 30113
rect 16945 30067 17003 30073
rect 18417 30073 18429 30107
rect 18463 30104 18475 30107
rect 19794 30104 19800 30116
rect 18463 30076 19800 30104
rect 18463 30073 18475 30076
rect 18417 30067 18475 30073
rect 19794 30064 19800 30076
rect 19852 30064 19858 30116
rect 20070 30064 20076 30116
rect 20128 30104 20134 30116
rect 20128 30076 21119 30104
rect 20128 30064 20134 30076
rect 2774 29996 2780 30048
rect 2832 30036 2838 30048
rect 2961 30039 3019 30045
rect 2961 30036 2973 30039
rect 2832 30008 2973 30036
rect 2832 29996 2838 30008
rect 2961 30005 2973 30008
rect 3007 30005 3019 30039
rect 2961 29999 3019 30005
rect 4890 29996 4896 30048
rect 4948 30036 4954 30048
rect 5629 30039 5687 30045
rect 5629 30036 5641 30039
rect 4948 30008 5641 30036
rect 4948 29996 4954 30008
rect 5629 30005 5641 30008
rect 5675 30005 5687 30039
rect 5629 29999 5687 30005
rect 8386 29996 8392 30048
rect 8444 29996 8450 30048
rect 8754 30036 8760 30048
rect 8715 30008 8760 30036
rect 8754 29996 8760 30008
rect 8812 29996 8818 30048
rect 11698 29996 11704 30048
rect 11756 30036 11762 30048
rect 11885 30039 11943 30045
rect 11885 30036 11897 30039
rect 11756 30008 11897 30036
rect 11756 29996 11762 30008
rect 11885 30005 11897 30008
rect 11931 30005 11943 30039
rect 11885 29999 11943 30005
rect 15933 30039 15991 30045
rect 15933 30005 15945 30039
rect 15979 30036 15991 30039
rect 16298 30036 16304 30048
rect 15979 30008 16304 30036
rect 15979 30005 15991 30008
rect 15933 29999 15991 30005
rect 16298 29996 16304 30008
rect 16356 29996 16362 30048
rect 17405 30039 17463 30045
rect 17405 30005 17417 30039
rect 17451 30036 17463 30039
rect 18690 30036 18696 30048
rect 17451 30008 18696 30036
rect 17451 30005 17463 30008
rect 17405 29999 17463 30005
rect 18690 29996 18696 30008
rect 18748 29996 18754 30048
rect 20622 29996 20628 30048
rect 20680 30036 20686 30048
rect 20993 30039 21051 30045
rect 20993 30036 21005 30039
rect 20680 30008 21005 30036
rect 20680 29996 20686 30008
rect 20993 30005 21005 30008
rect 21039 30005 21051 30039
rect 21091 30036 21119 30076
rect 22094 30064 22100 30116
rect 22152 30064 22158 30116
rect 23032 30036 23060 30203
rect 23658 30200 23664 30212
rect 23716 30200 23722 30252
rect 25976 30249 26004 30280
rect 26344 30252 26372 30280
rect 25041 30243 25099 30249
rect 25041 30209 25053 30243
rect 25087 30240 25099 30243
rect 25777 30243 25835 30249
rect 25777 30240 25789 30243
rect 25087 30212 25789 30240
rect 25087 30209 25099 30212
rect 25041 30203 25099 30209
rect 25777 30209 25789 30212
rect 25823 30209 25835 30243
rect 25777 30203 25835 30209
rect 25961 30243 26019 30249
rect 25961 30209 25973 30243
rect 26007 30209 26019 30243
rect 25961 30203 26019 30209
rect 26237 30243 26295 30249
rect 26237 30209 26249 30243
rect 26283 30240 26295 30243
rect 26326 30240 26332 30252
rect 26283 30212 26332 30240
rect 26283 30209 26295 30212
rect 26237 30203 26295 30209
rect 26326 30200 26332 30212
rect 26384 30200 26390 30252
rect 26418 30200 26424 30252
rect 26476 30240 26482 30252
rect 27264 30249 27292 30280
rect 27706 30268 27712 30320
rect 27764 30308 27770 30320
rect 28258 30308 28264 30320
rect 27764 30280 28264 30308
rect 27764 30268 27770 30280
rect 28258 30268 28264 30280
rect 28316 30268 28322 30320
rect 27249 30243 27307 30249
rect 26476 30212 26521 30240
rect 26476 30200 26482 30212
rect 27249 30209 27261 30243
rect 27295 30209 27307 30243
rect 30650 30240 30656 30252
rect 30611 30212 30656 30240
rect 27249 30203 27307 30209
rect 30650 30200 30656 30212
rect 30708 30200 30714 30252
rect 30742 30200 30748 30252
rect 30800 30240 30806 30252
rect 30929 30243 30987 30249
rect 30929 30240 30941 30243
rect 30800 30212 30941 30240
rect 30800 30200 30806 30212
rect 30929 30209 30941 30212
rect 30975 30209 30987 30243
rect 31110 30240 31116 30252
rect 31071 30212 31116 30240
rect 30929 30203 30987 30209
rect 31110 30200 31116 30212
rect 31168 30200 31174 30252
rect 23845 30175 23903 30181
rect 23845 30141 23857 30175
rect 23891 30141 23903 30175
rect 25314 30172 25320 30184
rect 25275 30144 25320 30172
rect 23845 30135 23903 30141
rect 23658 30064 23664 30116
rect 23716 30104 23722 30116
rect 23860 30104 23888 30135
rect 25314 30132 25320 30144
rect 25372 30132 25378 30184
rect 26973 30175 27031 30181
rect 26973 30141 26985 30175
rect 27019 30172 27031 30175
rect 27338 30172 27344 30184
rect 27019 30144 27344 30172
rect 27019 30141 27031 30144
rect 26973 30135 27031 30141
rect 27338 30132 27344 30144
rect 27396 30132 27402 30184
rect 29822 30172 29828 30184
rect 27448 30144 29828 30172
rect 23716 30076 23888 30104
rect 24857 30107 24915 30113
rect 23716 30064 23722 30076
rect 24857 30073 24869 30107
rect 24903 30104 24915 30107
rect 26602 30104 26608 30116
rect 24903 30076 26608 30104
rect 24903 30073 24915 30076
rect 24857 30067 24915 30073
rect 26602 30064 26608 30076
rect 26660 30064 26666 30116
rect 25222 30036 25228 30048
rect 21091 30008 23060 30036
rect 25183 30008 25228 30036
rect 20993 29999 21051 30005
rect 25222 29996 25228 30008
rect 25280 29996 25286 30048
rect 25774 29996 25780 30048
rect 25832 30036 25838 30048
rect 27448 30036 27476 30144
rect 29822 30132 29828 30144
rect 29880 30132 29886 30184
rect 28718 30064 28724 30116
rect 28776 30104 28782 30116
rect 30469 30107 30527 30113
rect 30469 30104 30481 30107
rect 28776 30076 30481 30104
rect 28776 30064 28782 30076
rect 30469 30073 30481 30076
rect 30515 30073 30527 30107
rect 30469 30067 30527 30073
rect 25832 30008 27476 30036
rect 25832 29996 25838 30008
rect 27522 29996 27528 30048
rect 27580 30036 27586 30048
rect 29549 30039 29607 30045
rect 29549 30036 29561 30039
rect 27580 30008 29561 30036
rect 27580 29996 27586 30008
rect 29549 30005 29561 30008
rect 29595 30036 29607 30039
rect 29914 30036 29920 30048
rect 29595 30008 29920 30036
rect 29595 30005 29607 30008
rect 29549 29999 29607 30005
rect 29914 29996 29920 30008
rect 29972 29996 29978 30048
rect 1104 29946 32016 29968
rect 0 29900 800 29914
rect 0 29872 888 29900
rect 1104 29894 2136 29946
rect 2188 29894 12440 29946
rect 12492 29894 22744 29946
rect 22796 29894 32016 29946
rect 32320 29900 33120 29914
rect 1104 29872 32016 29894
rect 32232 29872 33120 29900
rect 0 29858 800 29872
rect 860 29696 888 29872
rect 2777 29835 2835 29841
rect 2777 29801 2789 29835
rect 2823 29832 2835 29835
rect 3602 29832 3608 29844
rect 2823 29804 3608 29832
rect 2823 29801 2835 29804
rect 2777 29795 2835 29801
rect 3602 29792 3608 29804
rect 3660 29792 3666 29844
rect 6457 29835 6515 29841
rect 6457 29801 6469 29835
rect 6503 29832 6515 29835
rect 6546 29832 6552 29844
rect 6503 29804 6552 29832
rect 6503 29801 6515 29804
rect 6457 29795 6515 29801
rect 6546 29792 6552 29804
rect 6604 29792 6610 29844
rect 6641 29835 6699 29841
rect 6641 29801 6653 29835
rect 6687 29832 6699 29835
rect 7098 29832 7104 29844
rect 6687 29804 7104 29832
rect 6687 29801 6699 29804
rect 6641 29795 6699 29801
rect 7098 29792 7104 29804
rect 7156 29792 7162 29844
rect 7190 29792 7196 29844
rect 7248 29832 7254 29844
rect 12894 29832 12900 29844
rect 7248 29804 12900 29832
rect 7248 29792 7254 29804
rect 12894 29792 12900 29804
rect 12952 29792 12958 29844
rect 13078 29792 13084 29844
rect 13136 29832 13142 29844
rect 13446 29832 13452 29844
rect 13136 29804 13452 29832
rect 13136 29792 13142 29804
rect 13446 29792 13452 29804
rect 13504 29832 13510 29844
rect 13541 29835 13599 29841
rect 13541 29832 13553 29835
rect 13504 29804 13553 29832
rect 13504 29792 13510 29804
rect 13541 29801 13553 29804
rect 13587 29801 13599 29835
rect 13541 29795 13599 29801
rect 16574 29792 16580 29844
rect 16632 29832 16638 29844
rect 16632 29804 16804 29832
rect 16632 29792 16638 29804
rect 4246 29764 4252 29776
rect 768 29668 888 29696
rect 2746 29736 4252 29764
rect 768 29220 796 29668
rect 1394 29628 1400 29640
rect 1355 29600 1400 29628
rect 1394 29588 1400 29600
rect 1452 29628 1458 29640
rect 2746 29628 2774 29736
rect 4246 29724 4252 29736
rect 4304 29724 4310 29776
rect 5994 29764 6000 29776
rect 5000 29736 6000 29764
rect 3142 29656 3148 29708
rect 3200 29696 3206 29708
rect 5000 29696 5028 29736
rect 5994 29724 6000 29736
rect 6052 29724 6058 29776
rect 6362 29724 6368 29776
rect 6420 29764 6426 29776
rect 8202 29764 8208 29776
rect 6420 29736 8208 29764
rect 6420 29724 6426 29736
rect 8202 29724 8208 29736
rect 8260 29724 8266 29776
rect 8294 29724 8300 29776
rect 8352 29764 8358 29776
rect 8478 29764 8484 29776
rect 8352 29736 8484 29764
rect 8352 29724 8358 29736
rect 8478 29724 8484 29736
rect 8536 29724 8542 29776
rect 8662 29724 8668 29776
rect 8720 29764 8726 29776
rect 11701 29767 11759 29773
rect 8720 29736 9626 29764
rect 8720 29724 8726 29736
rect 5166 29696 5172 29708
rect 3200 29668 5028 29696
rect 5127 29668 5172 29696
rect 3200 29656 3206 29668
rect 5166 29656 5172 29668
rect 5224 29656 5230 29708
rect 6178 29656 6184 29708
rect 6236 29696 6242 29708
rect 6730 29696 6736 29708
rect 6236 29668 6736 29696
rect 6236 29656 6242 29668
rect 6730 29656 6736 29668
rect 6788 29696 6794 29708
rect 7374 29696 7380 29708
rect 6788 29668 7144 29696
rect 7287 29668 7380 29696
rect 6788 29656 6794 29668
rect 1452 29600 2774 29628
rect 1452 29588 1458 29600
rect 3694 29588 3700 29640
rect 3752 29628 3758 29640
rect 3973 29631 4031 29637
rect 3973 29628 3985 29631
rect 3752 29600 3985 29628
rect 3752 29588 3758 29600
rect 3973 29597 3985 29600
rect 4019 29597 4031 29631
rect 3973 29591 4031 29597
rect 4249 29631 4307 29637
rect 4249 29597 4261 29631
rect 4295 29597 4307 29631
rect 4249 29591 4307 29597
rect 4433 29631 4491 29637
rect 4433 29597 4445 29631
rect 4479 29628 4491 29631
rect 4798 29628 4804 29640
rect 4479 29600 4804 29628
rect 4479 29597 4491 29600
rect 4433 29591 4491 29597
rect 1664 29563 1722 29569
rect 1664 29529 1676 29563
rect 1710 29560 1722 29563
rect 2590 29560 2596 29572
rect 1710 29532 2596 29560
rect 1710 29529 1722 29532
rect 1664 29523 1722 29529
rect 2590 29520 2596 29532
rect 2648 29520 2654 29572
rect 4154 29520 4160 29572
rect 4212 29560 4218 29572
rect 4264 29560 4292 29591
rect 4798 29588 4804 29600
rect 4856 29588 4862 29640
rect 4893 29631 4951 29637
rect 4893 29597 4905 29631
rect 4939 29628 4951 29631
rect 4982 29628 4988 29640
rect 4939 29600 4988 29628
rect 4939 29597 4951 29600
rect 4893 29591 4951 29597
rect 4982 29588 4988 29600
rect 5040 29628 5046 29640
rect 7116 29637 7144 29668
rect 7374 29656 7380 29668
rect 7432 29696 7438 29708
rect 8680 29696 8708 29724
rect 9598 29705 9626 29736
rect 11701 29733 11713 29767
rect 11747 29764 11759 29767
rect 11882 29764 11888 29776
rect 11747 29736 11888 29764
rect 11747 29733 11759 29736
rect 11701 29727 11759 29733
rect 11882 29724 11888 29736
rect 11940 29724 11946 29776
rect 14182 29724 14188 29776
rect 14240 29764 14246 29776
rect 14553 29767 14611 29773
rect 14553 29764 14565 29767
rect 14240 29736 14565 29764
rect 14240 29724 14246 29736
rect 14553 29733 14565 29736
rect 14599 29733 14611 29767
rect 14553 29727 14611 29733
rect 16669 29767 16727 29773
rect 16669 29733 16681 29767
rect 16715 29733 16727 29767
rect 16776 29764 16804 29804
rect 17034 29792 17040 29844
rect 17092 29832 17098 29844
rect 19981 29835 20039 29841
rect 19981 29832 19993 29835
rect 17092 29804 19993 29832
rect 17092 29792 17098 29804
rect 19981 29801 19993 29804
rect 20027 29832 20039 29835
rect 20622 29832 20628 29844
rect 20027 29804 20628 29832
rect 20027 29801 20039 29804
rect 19981 29795 20039 29801
rect 20622 29792 20628 29804
rect 20680 29792 20686 29844
rect 20806 29832 20812 29844
rect 20767 29804 20812 29832
rect 20806 29792 20812 29804
rect 20864 29792 20870 29844
rect 20990 29792 20996 29844
rect 21048 29832 21054 29844
rect 23658 29832 23664 29844
rect 21048 29804 23664 29832
rect 21048 29792 21054 29804
rect 23658 29792 23664 29804
rect 23716 29792 23722 29844
rect 24949 29835 25007 29841
rect 24949 29801 24961 29835
rect 24995 29832 25007 29835
rect 26694 29832 26700 29844
rect 24995 29804 26700 29832
rect 24995 29801 25007 29804
rect 24949 29795 25007 29801
rect 26694 29792 26700 29804
rect 26752 29792 26758 29844
rect 30098 29792 30104 29844
rect 30156 29832 30162 29844
rect 31297 29835 31355 29841
rect 31297 29832 31309 29835
rect 30156 29804 31309 29832
rect 30156 29792 30162 29804
rect 31297 29801 31309 29804
rect 31343 29801 31355 29835
rect 31297 29795 31355 29801
rect 17129 29767 17187 29773
rect 17129 29764 17141 29767
rect 16776 29736 17141 29764
rect 16669 29727 16727 29733
rect 17129 29733 17141 29736
rect 17175 29733 17187 29767
rect 17129 29727 17187 29733
rect 7432 29668 8708 29696
rect 9217 29699 9275 29705
rect 7432 29656 7438 29668
rect 9217 29665 9229 29699
rect 9263 29696 9275 29699
rect 9585 29699 9643 29705
rect 9263 29668 9444 29696
rect 9263 29665 9275 29668
rect 9217 29659 9275 29665
rect 7101 29631 7159 29637
rect 5040 29600 6776 29628
rect 5040 29588 5046 29600
rect 5350 29560 5356 29572
rect 4212 29532 5356 29560
rect 4212 29520 4218 29532
rect 5350 29520 5356 29532
rect 5408 29520 5414 29572
rect 6273 29563 6331 29569
rect 6273 29529 6285 29563
rect 6319 29560 6331 29563
rect 6362 29560 6368 29572
rect 6319 29532 6368 29560
rect 6319 29529 6331 29532
rect 6273 29523 6331 29529
rect 6362 29520 6368 29532
rect 6420 29520 6426 29572
rect 3789 29495 3847 29501
rect 3789 29461 3801 29495
rect 3835 29492 3847 29495
rect 4338 29492 4344 29504
rect 3835 29464 4344 29492
rect 3835 29461 3847 29464
rect 3789 29455 3847 29461
rect 4338 29452 4344 29464
rect 4396 29452 4402 29504
rect 6178 29452 6184 29504
rect 6236 29492 6242 29504
rect 6473 29495 6531 29501
rect 6473 29492 6485 29495
rect 6236 29464 6485 29492
rect 6236 29452 6242 29464
rect 6473 29461 6485 29464
rect 6519 29461 6531 29495
rect 6748 29492 6776 29600
rect 7101 29597 7113 29631
rect 7147 29597 7159 29631
rect 7101 29591 7159 29597
rect 7650 29588 7656 29640
rect 7708 29628 7714 29640
rect 9113 29631 9171 29637
rect 9113 29628 9125 29631
rect 7708 29600 9125 29628
rect 7708 29588 7714 29600
rect 9113 29597 9125 29600
rect 9159 29597 9171 29631
rect 9416 29628 9444 29668
rect 9585 29665 9597 29699
rect 9631 29665 9643 29699
rect 16684 29696 16712 29727
rect 18598 29724 18604 29776
rect 18656 29764 18662 29776
rect 19518 29764 19524 29776
rect 18656 29736 19524 29764
rect 18656 29724 18662 29736
rect 19518 29724 19524 29736
rect 19576 29724 19582 29776
rect 20898 29724 20904 29776
rect 20956 29764 20962 29776
rect 21358 29764 21364 29776
rect 20956 29736 21364 29764
rect 20956 29724 20962 29736
rect 21358 29724 21364 29736
rect 21416 29724 21422 29776
rect 22830 29724 22836 29776
rect 22888 29764 22894 29776
rect 23201 29767 23259 29773
rect 23201 29764 23213 29767
rect 22888 29736 23213 29764
rect 22888 29724 22894 29736
rect 23201 29733 23213 29736
rect 23247 29733 23259 29767
rect 23201 29727 23259 29733
rect 25314 29724 25320 29776
rect 25372 29764 25378 29776
rect 32232 29764 32260 29872
rect 32320 29858 33120 29872
rect 25372 29736 25912 29764
rect 32232 29736 32352 29764
rect 25372 29724 25378 29736
rect 18230 29696 18236 29708
rect 9585 29659 9643 29665
rect 14384 29668 16712 29696
rect 17696 29668 18236 29696
rect 10226 29628 10232 29640
rect 9113 29591 9171 29597
rect 6822 29520 6828 29572
rect 6880 29560 6886 29572
rect 8662 29560 8668 29572
rect 6880 29532 8668 29560
rect 6880 29520 6886 29532
rect 8662 29520 8668 29532
rect 8720 29520 8726 29572
rect 8941 29563 8999 29569
rect 8941 29529 8953 29563
rect 8987 29560 8999 29563
rect 9214 29560 9220 29606
rect 8987 29554 9220 29560
rect 9272 29554 9278 29606
rect 9416 29600 10232 29628
rect 10226 29588 10232 29600
rect 10284 29588 10290 29640
rect 10321 29631 10379 29637
rect 10321 29597 10333 29631
rect 10367 29628 10379 29631
rect 12161 29631 12219 29637
rect 12161 29628 12173 29631
rect 10367 29600 12173 29628
rect 10367 29597 10379 29600
rect 10321 29591 10379 29597
rect 12161 29597 12173 29600
rect 12207 29628 12219 29631
rect 12986 29628 12992 29640
rect 12207 29600 12992 29628
rect 12207 29597 12219 29600
rect 12161 29591 12219 29597
rect 12986 29588 12992 29600
rect 13044 29588 13050 29640
rect 14090 29588 14096 29640
rect 14148 29628 14154 29640
rect 14384 29637 14412 29668
rect 14369 29631 14427 29637
rect 14148 29600 14320 29628
rect 14148 29588 14154 29600
rect 10588 29563 10646 29569
rect 8987 29532 9260 29554
rect 8987 29529 8999 29532
rect 8941 29523 8999 29529
rect 10588 29529 10600 29563
rect 10634 29560 10646 29563
rect 11514 29560 11520 29572
rect 10634 29532 11520 29560
rect 10634 29529 10646 29532
rect 10588 29523 10646 29529
rect 11514 29520 11520 29532
rect 11572 29520 11578 29572
rect 12428 29563 12486 29569
rect 12428 29529 12440 29563
rect 12474 29560 12486 29563
rect 14185 29563 14243 29569
rect 14185 29560 14197 29563
rect 12474 29532 14197 29560
rect 12474 29529 12486 29532
rect 12428 29523 12486 29529
rect 14185 29529 14197 29532
rect 14231 29529 14243 29563
rect 14292 29560 14320 29600
rect 14369 29597 14381 29631
rect 14415 29597 14427 29631
rect 14369 29591 14427 29597
rect 14645 29631 14703 29637
rect 14645 29597 14657 29631
rect 14691 29628 14703 29631
rect 15194 29628 15200 29640
rect 14691 29600 15200 29628
rect 14691 29597 14703 29600
rect 14645 29591 14703 29597
rect 15194 29588 15200 29600
rect 15252 29588 15258 29640
rect 15381 29631 15439 29637
rect 15381 29597 15393 29631
rect 15427 29597 15439 29631
rect 15654 29628 15660 29640
rect 15615 29600 15660 29628
rect 15381 29591 15439 29597
rect 15396 29560 15424 29591
rect 15654 29588 15660 29600
rect 15712 29588 15718 29640
rect 17696 29637 17724 29668
rect 18230 29656 18236 29668
rect 18288 29656 18294 29708
rect 19242 29656 19248 29708
rect 19300 29696 19306 29708
rect 21821 29699 21879 29705
rect 21821 29696 21833 29699
rect 19300 29668 21833 29696
rect 19300 29656 19306 29668
rect 21821 29665 21833 29668
rect 21867 29665 21879 29699
rect 21821 29659 21879 29665
rect 24578 29656 24584 29708
rect 24636 29696 24642 29708
rect 25501 29699 25559 29705
rect 25501 29696 25513 29699
rect 24636 29668 25513 29696
rect 24636 29656 24642 29668
rect 25501 29665 25513 29668
rect 25547 29665 25559 29699
rect 25682 29696 25688 29708
rect 25643 29668 25688 29696
rect 25501 29659 25559 29665
rect 25682 29656 25688 29668
rect 25740 29656 25746 29708
rect 25884 29705 25912 29736
rect 25869 29699 25927 29705
rect 25869 29665 25881 29699
rect 25915 29665 25927 29699
rect 26510 29696 26516 29708
rect 26471 29668 26516 29696
rect 25869 29659 25927 29665
rect 26510 29656 26516 29668
rect 26568 29656 26574 29708
rect 29914 29696 29920 29708
rect 29875 29668 29920 29696
rect 29914 29656 29920 29668
rect 29972 29656 29978 29708
rect 16945 29631 17003 29637
rect 16945 29597 16957 29631
rect 16991 29628 17003 29631
rect 17129 29631 17187 29637
rect 17129 29628 17141 29631
rect 16991 29600 17141 29628
rect 16991 29597 17003 29600
rect 16945 29591 17003 29597
rect 17129 29597 17141 29600
rect 17175 29597 17187 29631
rect 17129 29591 17187 29597
rect 17681 29631 17739 29637
rect 17681 29597 17693 29631
rect 17727 29597 17739 29631
rect 17954 29628 17960 29640
rect 17915 29600 17960 29628
rect 17681 29591 17739 29597
rect 17954 29588 17960 29600
rect 18012 29588 18018 29640
rect 18141 29631 18199 29637
rect 18141 29597 18153 29631
rect 18187 29628 18199 29631
rect 18322 29628 18328 29640
rect 18187 29600 18328 29628
rect 18187 29597 18199 29600
rect 18141 29591 18199 29597
rect 18322 29588 18328 29600
rect 18380 29588 18386 29640
rect 18616 29600 20024 29628
rect 16114 29560 16120 29572
rect 14292 29532 16120 29560
rect 14185 29523 14243 29529
rect 16114 29520 16120 29532
rect 16172 29520 16178 29572
rect 16298 29520 16304 29572
rect 16356 29560 16362 29572
rect 16669 29563 16727 29569
rect 16669 29560 16681 29563
rect 16356 29532 16681 29560
rect 16356 29520 16362 29532
rect 16669 29529 16681 29532
rect 16715 29560 16727 29563
rect 18616 29560 18644 29600
rect 16715 29532 18644 29560
rect 16715 29529 16727 29532
rect 16669 29523 16727 29529
rect 18690 29520 18696 29572
rect 18748 29560 18754 29572
rect 19889 29563 19947 29569
rect 19889 29560 19901 29563
rect 18748 29532 19901 29560
rect 18748 29520 18754 29532
rect 19889 29529 19901 29532
rect 19935 29529 19947 29563
rect 19996 29560 20024 29600
rect 20714 29588 20720 29640
rect 20772 29628 20778 29640
rect 20993 29631 21051 29637
rect 20993 29628 21005 29631
rect 20772 29600 21005 29628
rect 20772 29588 20778 29600
rect 20993 29597 21005 29600
rect 21039 29597 21051 29631
rect 20993 29591 21051 29597
rect 21085 29631 21143 29637
rect 21085 29597 21097 29631
rect 21131 29597 21143 29631
rect 21085 29591 21143 29597
rect 20809 29563 20867 29569
rect 20809 29560 20821 29563
rect 19996 29532 20821 29560
rect 19889 29523 19947 29529
rect 20809 29529 20821 29532
rect 20855 29560 20867 29563
rect 20898 29560 20904 29572
rect 20855 29532 20904 29560
rect 20855 29529 20867 29532
rect 20809 29523 20867 29529
rect 20898 29520 20904 29532
rect 20956 29520 20962 29572
rect 21100 29560 21128 29591
rect 21542 29588 21548 29640
rect 21600 29628 21606 29640
rect 23661 29631 23719 29637
rect 23661 29628 23673 29631
rect 21600 29600 23673 29628
rect 21600 29588 21606 29600
rect 23661 29597 23673 29600
rect 23707 29597 23719 29631
rect 25774 29628 25780 29640
rect 25735 29600 25780 29628
rect 23661 29591 23719 29597
rect 25774 29588 25780 29600
rect 25832 29588 25838 29640
rect 25958 29628 25964 29640
rect 25919 29600 25964 29628
rect 25958 29588 25964 29600
rect 26016 29588 26022 29640
rect 26528 29628 26556 29656
rect 27522 29628 27528 29640
rect 26528 29600 27528 29628
rect 27522 29588 27528 29600
rect 27580 29588 27586 29640
rect 28718 29628 28724 29640
rect 28679 29600 28724 29628
rect 28718 29588 28724 29600
rect 28776 29588 28782 29640
rect 28902 29628 28908 29640
rect 28863 29600 28908 29628
rect 28902 29588 28908 29600
rect 28960 29588 28966 29640
rect 28997 29631 29055 29637
rect 28997 29597 29009 29631
rect 29043 29628 29055 29631
rect 29270 29628 29276 29640
rect 29043 29600 29276 29628
rect 29043 29597 29055 29600
rect 28997 29591 29055 29597
rect 29270 29588 29276 29600
rect 29328 29588 29334 29640
rect 30006 29588 30012 29640
rect 30064 29628 30070 29640
rect 30173 29631 30231 29637
rect 30173 29628 30185 29631
rect 30064 29600 30185 29628
rect 30064 29588 30070 29600
rect 30173 29597 30185 29600
rect 30219 29597 30231 29631
rect 30173 29591 30231 29597
rect 21008 29532 21128 29560
rect 7926 29492 7932 29504
rect 6748 29464 7932 29492
rect 6473 29455 6531 29461
rect 7926 29452 7932 29464
rect 7984 29452 7990 29504
rect 8202 29452 8208 29504
rect 8260 29492 8266 29504
rect 9214 29492 9220 29504
rect 8260 29464 9220 29492
rect 8260 29452 8266 29464
rect 9214 29452 9220 29464
rect 9272 29492 9278 29504
rect 9309 29495 9367 29501
rect 9309 29492 9321 29495
rect 9272 29464 9321 29492
rect 9272 29452 9278 29464
rect 9309 29461 9321 29464
rect 9355 29461 9367 29495
rect 9490 29492 9496 29504
rect 9451 29464 9496 29492
rect 9309 29455 9367 29461
rect 9490 29452 9496 29464
rect 9548 29452 9554 29504
rect 9858 29452 9864 29504
rect 9916 29492 9922 29504
rect 12250 29492 12256 29504
rect 9916 29464 12256 29492
rect 9916 29452 9922 29464
rect 12250 29452 12256 29464
rect 12308 29452 12314 29504
rect 13170 29452 13176 29504
rect 13228 29492 13234 29504
rect 16853 29495 16911 29501
rect 16853 29492 16865 29495
rect 13228 29464 16865 29492
rect 13228 29452 13234 29464
rect 16853 29461 16865 29464
rect 16899 29461 16911 29495
rect 16853 29455 16911 29461
rect 17310 29452 17316 29504
rect 17368 29492 17374 29504
rect 17497 29495 17555 29501
rect 17497 29492 17509 29495
rect 17368 29464 17509 29492
rect 17368 29452 17374 29464
rect 17497 29461 17509 29464
rect 17543 29461 17555 29495
rect 17497 29455 17555 29461
rect 17678 29452 17684 29504
rect 17736 29492 17742 29504
rect 20438 29492 20444 29504
rect 17736 29464 20444 29492
rect 17736 29452 17742 29464
rect 20438 29452 20444 29464
rect 20496 29492 20502 29504
rect 21008 29492 21036 29532
rect 21910 29520 21916 29572
rect 21968 29560 21974 29572
rect 22066 29563 22124 29569
rect 22066 29560 22078 29563
rect 21968 29532 22078 29560
rect 21968 29520 21974 29532
rect 22066 29529 22078 29532
rect 22112 29529 22124 29563
rect 22066 29523 22124 29529
rect 23106 29520 23112 29572
rect 23164 29560 23170 29572
rect 23474 29560 23480 29572
rect 23164 29532 23480 29560
rect 23164 29520 23170 29532
rect 23474 29520 23480 29532
rect 23532 29520 23538 29572
rect 24857 29563 24915 29569
rect 24857 29529 24869 29563
rect 24903 29560 24915 29563
rect 26050 29560 26056 29572
rect 24903 29532 26056 29560
rect 24903 29529 24915 29532
rect 24857 29523 24915 29529
rect 26050 29520 26056 29532
rect 26108 29520 26114 29572
rect 26602 29520 26608 29572
rect 26660 29560 26666 29572
rect 26758 29563 26816 29569
rect 26758 29560 26770 29563
rect 26660 29532 26770 29560
rect 26660 29520 26666 29532
rect 26758 29529 26770 29532
rect 26804 29529 26816 29563
rect 26758 29523 26816 29529
rect 29730 29520 29736 29572
rect 29788 29560 29794 29572
rect 30374 29560 30380 29572
rect 29788 29532 30380 29560
rect 29788 29520 29794 29532
rect 30374 29520 30380 29532
rect 30432 29520 30438 29572
rect 20496 29464 21036 29492
rect 20496 29452 20502 29464
rect 22186 29452 22192 29504
rect 22244 29492 22250 29504
rect 22922 29492 22928 29504
rect 22244 29464 22928 29492
rect 22244 29452 22250 29464
rect 22922 29452 22928 29464
rect 22980 29452 22986 29504
rect 23750 29492 23756 29504
rect 23711 29464 23756 29492
rect 23750 29452 23756 29464
rect 23808 29452 23814 29504
rect 24394 29452 24400 29504
rect 24452 29492 24458 29504
rect 24670 29492 24676 29504
rect 24452 29464 24676 29492
rect 24452 29452 24458 29464
rect 24670 29452 24676 29464
rect 24728 29452 24734 29504
rect 26418 29452 26424 29504
rect 26476 29492 26482 29504
rect 27893 29495 27951 29501
rect 27893 29492 27905 29495
rect 26476 29464 27905 29492
rect 26476 29452 26482 29464
rect 27893 29461 27905 29464
rect 27939 29461 27951 29495
rect 27893 29455 27951 29461
rect 28537 29495 28595 29501
rect 28537 29461 28549 29495
rect 28583 29492 28595 29495
rect 30006 29492 30012 29504
rect 28583 29464 30012 29492
rect 28583 29461 28595 29464
rect 28537 29455 28595 29461
rect 30006 29452 30012 29464
rect 30064 29452 30070 29504
rect 1104 29402 32016 29424
rect 1104 29350 7288 29402
rect 7340 29350 17592 29402
rect 17644 29350 27896 29402
rect 27948 29350 32016 29402
rect 1104 29328 32016 29350
rect 1673 29291 1731 29297
rect 1673 29257 1685 29291
rect 1719 29288 1731 29291
rect 3142 29288 3148 29300
rect 1719 29260 3148 29288
rect 1719 29257 1731 29260
rect 1673 29251 1731 29257
rect 3142 29248 3148 29260
rect 3200 29248 3206 29300
rect 3252 29260 4752 29288
rect 1581 29223 1639 29229
rect 1581 29220 1593 29223
rect 768 29192 1593 29220
rect 1581 29189 1593 29192
rect 1627 29189 1639 29223
rect 1581 29183 1639 29189
rect 2409 29155 2467 29161
rect 2409 29121 2421 29155
rect 2455 29152 2467 29155
rect 3145 29155 3203 29161
rect 3145 29152 3157 29155
rect 2455 29124 3157 29152
rect 2455 29121 2467 29124
rect 2409 29115 2467 29121
rect 3145 29121 3157 29124
rect 3191 29121 3203 29155
rect 3145 29115 3203 29121
rect 2685 29087 2743 29093
rect 2685 29053 2697 29087
rect 2731 29084 2743 29087
rect 3252 29084 3280 29260
rect 3694 29220 3700 29232
rect 3344 29192 3700 29220
rect 3344 29161 3372 29192
rect 3694 29180 3700 29192
rect 3752 29180 3758 29232
rect 4724 29220 4752 29260
rect 4798 29248 4804 29300
rect 4856 29288 4862 29300
rect 5813 29291 5871 29297
rect 5813 29288 5825 29291
rect 4856 29260 5825 29288
rect 4856 29248 4862 29260
rect 5813 29257 5825 29260
rect 5859 29257 5871 29291
rect 5813 29251 5871 29257
rect 7101 29291 7159 29297
rect 7101 29257 7113 29291
rect 7147 29288 7159 29291
rect 7466 29288 7472 29300
rect 7147 29260 7472 29288
rect 7147 29257 7159 29260
rect 7101 29251 7159 29257
rect 4890 29220 4896 29232
rect 4724 29192 4896 29220
rect 4890 29180 4896 29192
rect 4948 29180 4954 29232
rect 3329 29155 3387 29161
rect 3329 29121 3341 29155
rect 3375 29121 3387 29155
rect 3329 29115 3387 29121
rect 3605 29155 3663 29161
rect 3605 29121 3617 29155
rect 3651 29121 3663 29155
rect 3786 29152 3792 29164
rect 3747 29124 3792 29152
rect 3605 29115 3663 29121
rect 2731 29056 3280 29084
rect 3620 29084 3648 29115
rect 3786 29112 3792 29124
rect 3844 29112 3850 29164
rect 4246 29112 4252 29164
rect 4304 29152 4310 29164
rect 4433 29155 4491 29161
rect 4433 29152 4445 29155
rect 4304 29124 4445 29152
rect 4304 29112 4310 29124
rect 4433 29121 4445 29124
rect 4479 29121 4491 29155
rect 4433 29115 4491 29121
rect 4522 29112 4528 29164
rect 4580 29152 4586 29164
rect 4689 29155 4747 29161
rect 4689 29152 4701 29155
rect 4580 29124 4701 29152
rect 4580 29112 4586 29124
rect 4689 29121 4701 29124
rect 4735 29121 4747 29155
rect 4908 29152 4936 29180
rect 5828 29152 5856 29251
rect 7466 29248 7472 29260
rect 7524 29248 7530 29300
rect 7852 29260 8064 29288
rect 6641 29223 6699 29229
rect 6641 29189 6653 29223
rect 6687 29220 6699 29223
rect 7852 29220 7880 29260
rect 6687 29192 7880 29220
rect 8036 29220 8064 29260
rect 9214 29248 9220 29300
rect 9272 29288 9278 29300
rect 9272 29260 9904 29288
rect 9272 29248 9278 29260
rect 9766 29220 9772 29232
rect 8036 29192 8423 29220
rect 6687 29189 6699 29192
rect 6641 29183 6699 29189
rect 6917 29155 6975 29161
rect 6917 29152 6929 29155
rect 4908 29124 5764 29152
rect 5828 29124 6929 29152
rect 4689 29115 4747 29121
rect 4154 29084 4160 29096
rect 3620 29056 4160 29084
rect 2731 29053 2743 29056
rect 2685 29047 2743 29053
rect 4154 29044 4160 29056
rect 4212 29044 4218 29096
rect 2593 29019 2651 29025
rect 2593 28985 2605 29019
rect 2639 29016 2651 29019
rect 5736 29016 5764 29124
rect 6917 29121 6929 29124
rect 6963 29121 6975 29155
rect 6917 29115 6975 29121
rect 7285 29155 7343 29161
rect 7285 29121 7297 29155
rect 7331 29152 7343 29155
rect 7374 29152 7380 29164
rect 7331 29124 7380 29152
rect 7331 29121 7343 29124
rect 7285 29115 7343 29121
rect 7374 29112 7380 29124
rect 7432 29112 7438 29164
rect 7926 29152 7932 29164
rect 7887 29124 7932 29152
rect 7926 29112 7932 29124
rect 7984 29112 7990 29164
rect 8021 29155 8079 29161
rect 8021 29121 8033 29155
rect 8067 29121 8079 29155
rect 8021 29115 8079 29121
rect 8205 29155 8263 29161
rect 8205 29121 8217 29155
rect 8251 29121 8263 29155
rect 8205 29115 8263 29121
rect 8307 29155 8365 29161
rect 8307 29121 8319 29155
rect 8353 29152 8365 29155
rect 8395 29152 8423 29192
rect 9324 29192 9772 29220
rect 9324 29161 9352 29192
rect 9766 29180 9772 29192
rect 9824 29180 9830 29232
rect 9876 29220 9904 29260
rect 10226 29248 10232 29300
rect 10284 29288 10290 29300
rect 10689 29291 10747 29297
rect 10689 29288 10701 29291
rect 10284 29260 10701 29288
rect 10284 29248 10290 29260
rect 10689 29257 10701 29260
rect 10735 29257 10747 29291
rect 10689 29251 10747 29257
rect 11514 29248 11520 29300
rect 11572 29288 11578 29300
rect 12989 29291 13047 29297
rect 12989 29288 13001 29291
rect 11572 29260 13001 29288
rect 11572 29248 11578 29260
rect 12989 29257 13001 29260
rect 13035 29257 13047 29291
rect 12989 29251 13047 29257
rect 13096 29260 15792 29288
rect 9876 29192 11284 29220
rect 8353 29124 8423 29152
rect 9309 29155 9367 29161
rect 8353 29121 8365 29124
rect 8307 29115 8365 29121
rect 9309 29121 9321 29155
rect 9355 29121 9367 29155
rect 9309 29115 9367 29121
rect 9576 29155 9634 29161
rect 9576 29121 9588 29155
rect 9622 29152 9634 29155
rect 11146 29152 11152 29164
rect 9622 29124 11152 29152
rect 9622 29121 9634 29124
rect 9576 29115 9634 29121
rect 6822 29084 6828 29096
rect 6783 29056 6828 29084
rect 6822 29044 6828 29056
rect 6880 29044 6886 29096
rect 7006 29044 7012 29096
rect 7064 29084 7070 29096
rect 7193 29087 7251 29093
rect 7193 29084 7205 29087
rect 7064 29056 7205 29084
rect 7064 29044 7070 29056
rect 7193 29053 7205 29056
rect 7239 29084 7251 29087
rect 7466 29084 7472 29096
rect 7239 29056 7472 29084
rect 7239 29053 7251 29056
rect 7193 29047 7251 29053
rect 7466 29044 7472 29056
rect 7524 29044 7530 29096
rect 8036 29084 8064 29115
rect 7668 29056 8064 29084
rect 7668 29016 7696 29056
rect 8220 29028 8248 29115
rect 11146 29112 11152 29124
rect 11204 29112 11210 29164
rect 11256 29084 11284 29192
rect 12894 29180 12900 29232
rect 12952 29220 12958 29232
rect 13096 29220 13124 29260
rect 12952 29192 13124 29220
rect 12952 29180 12958 29192
rect 13630 29180 13636 29232
rect 13688 29220 13694 29232
rect 14826 29220 14832 29232
rect 13688 29192 14832 29220
rect 13688 29180 13694 29192
rect 14826 29180 14832 29192
rect 14884 29180 14890 29232
rect 15654 29220 15660 29232
rect 15396 29192 15660 29220
rect 11517 29155 11575 29161
rect 11517 29121 11529 29155
rect 11563 29152 11575 29155
rect 11563 29124 12020 29152
rect 11563 29121 11575 29124
rect 11517 29115 11575 29121
rect 11793 29087 11851 29093
rect 11793 29084 11805 29087
rect 11256 29056 11805 29084
rect 11793 29053 11805 29056
rect 11839 29053 11851 29087
rect 11992 29084 12020 29124
rect 12066 29112 12072 29164
rect 12124 29152 12130 29164
rect 13173 29155 13231 29161
rect 13173 29152 13185 29155
rect 12124 29124 13185 29152
rect 12124 29112 12130 29124
rect 13173 29121 13185 29124
rect 13219 29121 13231 29155
rect 13446 29152 13452 29164
rect 13407 29124 13452 29152
rect 13173 29115 13231 29121
rect 13446 29112 13452 29124
rect 13504 29112 13510 29164
rect 14185 29155 14243 29161
rect 14185 29121 14197 29155
rect 14231 29152 14243 29155
rect 14921 29155 14979 29161
rect 14921 29152 14933 29155
rect 14231 29124 14933 29152
rect 14231 29121 14243 29124
rect 14185 29115 14243 29121
rect 14921 29121 14933 29124
rect 14967 29121 14979 29155
rect 14921 29115 14979 29121
rect 15105 29155 15163 29161
rect 15105 29121 15117 29155
rect 15151 29152 15163 29155
rect 15286 29152 15292 29164
rect 15151 29124 15292 29152
rect 15151 29121 15163 29124
rect 15105 29115 15163 29121
rect 15286 29112 15292 29124
rect 15344 29112 15350 29164
rect 15396 29161 15424 29192
rect 15654 29180 15660 29192
rect 15712 29180 15718 29232
rect 15764 29220 15792 29260
rect 17126 29248 17132 29300
rect 17184 29288 17190 29300
rect 17770 29288 17776 29300
rect 17184 29260 17776 29288
rect 17184 29248 17190 29260
rect 17770 29248 17776 29260
rect 17828 29248 17834 29300
rect 20990 29248 20996 29300
rect 21048 29288 21054 29300
rect 21085 29291 21143 29297
rect 21085 29288 21097 29291
rect 21048 29260 21097 29288
rect 21048 29248 21054 29260
rect 21085 29257 21097 29260
rect 21131 29257 21143 29291
rect 21085 29251 21143 29257
rect 21821 29291 21879 29297
rect 21821 29257 21833 29291
rect 21867 29288 21879 29291
rect 21910 29288 21916 29300
rect 21867 29260 21916 29288
rect 21867 29257 21879 29260
rect 21821 29251 21879 29257
rect 21910 29248 21916 29260
rect 21968 29248 21974 29300
rect 22186 29288 22192 29300
rect 22020 29260 22192 29288
rect 15764 29192 21956 29220
rect 15381 29155 15439 29161
rect 15381 29121 15393 29155
rect 15427 29121 15439 29155
rect 15381 29115 15439 29121
rect 15565 29155 15623 29161
rect 15565 29121 15577 29155
rect 15611 29121 15623 29155
rect 15565 29115 15623 29121
rect 12526 29084 12532 29096
rect 11992 29056 12532 29084
rect 11793 29047 11851 29053
rect 12526 29044 12532 29056
rect 12584 29084 12590 29096
rect 12986 29084 12992 29096
rect 12584 29056 12992 29084
rect 12584 29044 12590 29056
rect 12986 29044 12992 29056
rect 13044 29044 13050 29096
rect 14090 29084 14096 29096
rect 13280 29056 14096 29084
rect 2639 28988 4200 29016
rect 5736 28988 7696 29016
rect 2639 28985 2651 28988
rect 2593 28979 2651 28985
rect 2222 28948 2228 28960
rect 2183 28920 2228 28948
rect 2222 28908 2228 28920
rect 2280 28908 2286 28960
rect 4172 28948 4200 28988
rect 8202 28976 8208 29028
rect 8260 28976 8266 29028
rect 10594 28976 10600 29028
rect 10652 29016 10658 29028
rect 13280 29016 13308 29056
rect 14090 29044 14096 29056
rect 14148 29044 14154 29096
rect 14366 29084 14372 29096
rect 14327 29056 14372 29084
rect 14366 29044 14372 29056
rect 14424 29044 14430 29096
rect 14461 29087 14519 29093
rect 14461 29053 14473 29087
rect 14507 29084 14519 29087
rect 14642 29084 14648 29096
rect 14507 29056 14648 29084
rect 14507 29053 14519 29056
rect 14461 29047 14519 29053
rect 14642 29044 14648 29056
rect 14700 29044 14706 29096
rect 15194 29044 15200 29096
rect 15252 29084 15258 29096
rect 15580 29084 15608 29115
rect 16666 29112 16672 29164
rect 16724 29152 16730 29164
rect 17129 29155 17187 29161
rect 17129 29152 17141 29155
rect 16724 29124 17141 29152
rect 16724 29112 16730 29124
rect 17129 29121 17141 29124
rect 17175 29121 17187 29155
rect 17310 29152 17316 29164
rect 17271 29124 17316 29152
rect 17129 29115 17187 29121
rect 17310 29112 17316 29124
rect 17368 29112 17374 29164
rect 17402 29112 17408 29164
rect 17460 29152 17466 29164
rect 17678 29152 17684 29164
rect 17460 29124 17684 29152
rect 17460 29112 17466 29124
rect 17678 29112 17684 29124
rect 17736 29112 17742 29164
rect 18601 29155 18659 29161
rect 18601 29121 18613 29155
rect 18647 29152 18659 29155
rect 19426 29152 19432 29164
rect 18647 29124 19432 29152
rect 18647 29121 18659 29124
rect 18601 29115 18659 29121
rect 19426 29112 19432 29124
rect 19484 29112 19490 29164
rect 20993 29155 21051 29161
rect 20993 29121 21005 29155
rect 21039 29121 21051 29155
rect 20993 29115 21051 29121
rect 15252 29056 15608 29084
rect 15252 29044 15258 29056
rect 17034 29044 17040 29096
rect 17092 29084 17098 29096
rect 17497 29087 17555 29093
rect 17497 29084 17509 29087
rect 17092 29056 17509 29084
rect 17092 29044 17098 29056
rect 17497 29053 17509 29056
rect 17543 29053 17555 29087
rect 17497 29047 17555 29053
rect 17589 29087 17647 29093
rect 17589 29053 17601 29087
rect 17635 29084 17647 29087
rect 17954 29084 17960 29096
rect 17635 29056 17960 29084
rect 17635 29053 17647 29056
rect 17589 29047 17647 29053
rect 17954 29044 17960 29056
rect 18012 29084 18018 29096
rect 18138 29084 18144 29096
rect 18012 29056 18144 29084
rect 18012 29044 18018 29056
rect 18138 29044 18144 29056
rect 18196 29044 18202 29096
rect 18690 29044 18696 29096
rect 18748 29084 18754 29096
rect 21008 29084 21036 29115
rect 18748 29056 21036 29084
rect 21928 29084 21956 29192
rect 22020 29161 22048 29260
rect 22186 29248 22192 29260
rect 22244 29248 22250 29300
rect 22465 29291 22523 29297
rect 22465 29257 22477 29291
rect 22511 29288 22523 29291
rect 22922 29288 22928 29300
rect 22511 29260 22928 29288
rect 22511 29257 22523 29260
rect 22465 29251 22523 29257
rect 22922 29248 22928 29260
rect 22980 29248 22986 29300
rect 24118 29248 24124 29300
rect 24176 29288 24182 29300
rect 28537 29291 28595 29297
rect 28537 29288 28549 29291
rect 24176 29260 28549 29288
rect 24176 29248 24182 29260
rect 28537 29257 28549 29260
rect 28583 29257 28595 29291
rect 32324 29288 32352 29736
rect 28537 29251 28595 29257
rect 28966 29260 32352 29288
rect 25777 29223 25835 29229
rect 22112 29192 25728 29220
rect 22005 29155 22063 29161
rect 22005 29121 22017 29155
rect 22051 29121 22063 29155
rect 22005 29115 22063 29121
rect 22112 29084 22140 29192
rect 22189 29155 22247 29161
rect 22189 29121 22201 29155
rect 22235 29152 22247 29155
rect 22462 29152 22468 29164
rect 22235 29124 22468 29152
rect 22235 29121 22247 29124
rect 22189 29115 22247 29121
rect 21928 29056 22140 29084
rect 18748 29044 18754 29056
rect 10652 28988 13308 29016
rect 13357 29019 13415 29025
rect 10652 28976 10658 28988
rect 13357 28985 13369 29019
rect 13403 29016 13415 29019
rect 13906 29016 13912 29028
rect 13403 28988 13912 29016
rect 13403 28985 13415 28988
rect 13357 28979 13415 28985
rect 13906 28976 13912 28988
rect 13964 28976 13970 29028
rect 14001 29019 14059 29025
rect 14001 28985 14013 29019
rect 14047 29016 14059 29019
rect 14734 29016 14740 29028
rect 14047 28988 14740 29016
rect 14047 28985 14059 28988
rect 14001 28979 14059 28985
rect 14734 28976 14740 28988
rect 14792 28976 14798 29028
rect 17126 28976 17132 29028
rect 17184 29016 17190 29028
rect 18782 29016 18788 29028
rect 17184 28988 18788 29016
rect 17184 28976 17190 28988
rect 18782 28976 18788 28988
rect 18840 28976 18846 29028
rect 19242 28976 19248 29028
rect 19300 29016 19306 29028
rect 19889 29019 19947 29025
rect 19889 29016 19901 29019
rect 19300 28988 19901 29016
rect 19300 28976 19306 28988
rect 19889 28985 19901 28988
rect 19935 28985 19947 29019
rect 19889 28979 19947 28985
rect 20990 28976 20996 29028
rect 21048 29016 21054 29028
rect 22204 29016 22232 29115
rect 22462 29112 22468 29124
rect 22520 29112 22526 29164
rect 22554 29112 22560 29164
rect 22612 29152 22618 29164
rect 22741 29155 22799 29161
rect 22741 29152 22753 29155
rect 22612 29124 22753 29152
rect 22612 29112 22618 29124
rect 22741 29121 22753 29124
rect 22787 29121 22799 29155
rect 22741 29115 22799 29121
rect 22833 29155 22891 29161
rect 22833 29121 22845 29155
rect 22879 29121 22891 29155
rect 23106 29152 23112 29164
rect 23067 29124 23112 29152
rect 22833 29115 22891 29121
rect 22281 29087 22339 29093
rect 22281 29053 22293 29087
rect 22327 29084 22339 29087
rect 22646 29084 22652 29096
rect 22327 29056 22652 29084
rect 22327 29053 22339 29056
rect 22281 29047 22339 29053
rect 22646 29044 22652 29056
rect 22704 29084 22710 29096
rect 22848 29084 22876 29115
rect 23106 29112 23112 29124
rect 23164 29112 23170 29164
rect 24118 29152 24124 29164
rect 24079 29124 24124 29152
rect 24118 29112 24124 29124
rect 24176 29112 24182 29164
rect 24397 29155 24455 29161
rect 24397 29121 24409 29155
rect 24443 29121 24455 29155
rect 24397 29115 24455 29121
rect 24489 29155 24547 29161
rect 24489 29121 24501 29155
rect 24535 29121 24547 29155
rect 24489 29115 24547 29121
rect 24581 29155 24639 29161
rect 24581 29121 24593 29155
rect 24627 29152 24639 29155
rect 24670 29152 24676 29164
rect 24627 29124 24676 29152
rect 24627 29121 24639 29124
rect 24581 29115 24639 29121
rect 22704 29056 22876 29084
rect 22925 29087 22983 29093
rect 22704 29044 22710 29056
rect 22925 29053 22937 29087
rect 22971 29084 22983 29087
rect 23014 29084 23020 29096
rect 22971 29056 23020 29084
rect 22971 29053 22983 29056
rect 22925 29047 22983 29053
rect 23014 29044 23020 29056
rect 23072 29044 23078 29096
rect 24210 29044 24216 29096
rect 24268 29084 24274 29096
rect 24412 29084 24440 29115
rect 24268 29056 24440 29084
rect 24504 29084 24532 29115
rect 24670 29112 24676 29124
rect 24728 29112 24734 29164
rect 24765 29155 24823 29161
rect 24765 29121 24777 29155
rect 24811 29152 24823 29155
rect 25700 29152 25728 29192
rect 25777 29189 25789 29223
rect 25823 29220 25835 29223
rect 25866 29220 25872 29232
rect 25823 29192 25872 29220
rect 25823 29189 25835 29192
rect 25777 29183 25835 29189
rect 25866 29180 25872 29192
rect 25924 29180 25930 29232
rect 28966 29220 28994 29260
rect 25976 29192 28994 29220
rect 25976 29152 26004 29192
rect 28074 29152 28080 29164
rect 24811 29124 25636 29152
rect 25700 29124 26004 29152
rect 27172 29124 28080 29152
rect 24811 29121 24823 29124
rect 24765 29115 24823 29121
rect 24857 29087 24915 29093
rect 24504 29056 24808 29084
rect 24268 29044 24274 29056
rect 21048 28988 22232 29016
rect 23109 29019 23167 29025
rect 21048 28976 21054 28988
rect 23109 28985 23121 29019
rect 23155 29016 23167 29019
rect 24670 29016 24676 29028
rect 23155 28988 24676 29016
rect 23155 28985 23167 28988
rect 23109 28979 23167 28985
rect 24670 28976 24676 28988
rect 24728 28976 24734 29028
rect 24780 29016 24808 29056
rect 24857 29053 24869 29087
rect 24903 29084 24915 29087
rect 24946 29084 24952 29096
rect 24903 29056 24952 29084
rect 24903 29053 24915 29056
rect 24857 29047 24915 29053
rect 24946 29044 24952 29056
rect 25004 29044 25010 29096
rect 25130 29044 25136 29096
rect 25188 29084 25194 29096
rect 25409 29087 25467 29093
rect 25409 29084 25421 29087
rect 25188 29056 25421 29084
rect 25188 29044 25194 29056
rect 25409 29053 25421 29056
rect 25455 29053 25467 29087
rect 25608 29084 25636 29124
rect 27172 29096 27200 29124
rect 28074 29112 28080 29124
rect 28132 29112 28138 29164
rect 28350 29152 28356 29164
rect 28311 29124 28356 29152
rect 28350 29112 28356 29124
rect 28408 29112 28414 29164
rect 29270 29112 29276 29164
rect 29328 29152 29334 29164
rect 29365 29155 29423 29161
rect 29365 29152 29377 29155
rect 29328 29124 29377 29152
rect 29328 29112 29334 29124
rect 29365 29121 29377 29124
rect 29411 29121 29423 29155
rect 29365 29115 29423 29121
rect 27065 29087 27123 29093
rect 25608 29056 27016 29084
rect 25409 29047 25467 29053
rect 26510 29016 26516 29028
rect 24780 28988 26516 29016
rect 26510 28976 26516 28988
rect 26568 28976 26574 29028
rect 26988 29016 27016 29056
rect 27065 29053 27077 29087
rect 27111 29084 27123 29087
rect 27154 29084 27160 29096
rect 27111 29056 27160 29084
rect 27111 29053 27123 29056
rect 27065 29047 27123 29053
rect 27154 29044 27160 29056
rect 27212 29044 27218 29096
rect 27338 29084 27344 29096
rect 27299 29056 27344 29084
rect 27338 29044 27344 29056
rect 27396 29044 27402 29096
rect 29178 29084 29184 29096
rect 29139 29056 29184 29084
rect 29178 29044 29184 29056
rect 29236 29044 29242 29096
rect 29380 29084 29408 29115
rect 30098 29112 30104 29164
rect 30156 29152 30162 29164
rect 30374 29152 30380 29164
rect 30156 29124 30201 29152
rect 30335 29124 30380 29152
rect 30156 29112 30162 29124
rect 30374 29112 30380 29124
rect 30432 29112 30438 29164
rect 29380 29056 29960 29084
rect 27798 29016 27804 29028
rect 26988 28988 27804 29016
rect 27798 28976 27804 28988
rect 27856 28976 27862 29028
rect 29822 29016 29828 29028
rect 29783 28988 29828 29016
rect 29822 28976 29828 28988
rect 29880 28976 29886 29028
rect 4430 28948 4436 28960
rect 4172 28920 4436 28948
rect 4430 28908 4436 28920
rect 4488 28948 4494 28960
rect 5166 28948 5172 28960
rect 4488 28920 5172 28948
rect 4488 28908 4494 28920
rect 5166 28908 5172 28920
rect 5224 28908 5230 28960
rect 7745 28951 7803 28957
rect 7745 28917 7757 28951
rect 7791 28948 7803 28951
rect 8110 28948 8116 28960
rect 7791 28920 8116 28948
rect 7791 28917 7803 28920
rect 7745 28911 7803 28917
rect 8110 28908 8116 28920
rect 8168 28908 8174 28960
rect 9122 28908 9128 28960
rect 9180 28948 9186 28960
rect 9490 28948 9496 28960
rect 9180 28920 9496 28948
rect 9180 28908 9186 28920
rect 9490 28908 9496 28920
rect 9548 28908 9554 28960
rect 10502 28908 10508 28960
rect 10560 28948 10566 28960
rect 11514 28948 11520 28960
rect 10560 28920 11520 28948
rect 10560 28908 10566 28920
rect 11514 28908 11520 28920
rect 11572 28908 11578 28960
rect 12710 28908 12716 28960
rect 12768 28948 12774 28960
rect 20254 28948 20260 28960
rect 12768 28920 20260 28948
rect 12768 28908 12774 28920
rect 20254 28908 20260 28920
rect 20312 28908 20318 28960
rect 21174 28908 21180 28960
rect 21232 28948 21238 28960
rect 22186 28948 22192 28960
rect 21232 28920 22192 28948
rect 21232 28908 21238 28920
rect 22186 28908 22192 28920
rect 22244 28908 22250 28960
rect 22462 28948 22468 28960
rect 22423 28920 22468 28948
rect 22462 28908 22468 28920
rect 22520 28908 22526 28960
rect 24210 28908 24216 28960
rect 24268 28948 24274 28960
rect 24578 28948 24584 28960
rect 24268 28920 24584 28948
rect 24268 28908 24274 28920
rect 24578 28908 24584 28920
rect 24636 28908 24642 28960
rect 25682 28908 25688 28960
rect 25740 28948 25746 28960
rect 25777 28951 25835 28957
rect 25777 28948 25789 28951
rect 25740 28920 25789 28948
rect 25740 28908 25746 28920
rect 25777 28917 25789 28920
rect 25823 28917 25835 28951
rect 25958 28948 25964 28960
rect 25919 28920 25964 28948
rect 25777 28911 25835 28917
rect 25958 28908 25964 28920
rect 26016 28908 26022 28960
rect 26878 28908 26884 28960
rect 26936 28948 26942 28960
rect 29730 28948 29736 28960
rect 26936 28920 29736 28948
rect 26936 28908 26942 28920
rect 29730 28908 29736 28920
rect 29788 28908 29794 28960
rect 29932 28948 29960 29056
rect 30190 29044 30196 29096
rect 30248 29093 30254 29096
rect 30248 29087 30276 29093
rect 30264 29053 30276 29087
rect 30248 29047 30276 29053
rect 30248 29044 30254 29047
rect 30834 28948 30840 28960
rect 29932 28920 30840 28948
rect 30834 28908 30840 28920
rect 30892 28908 30898 28960
rect 31018 28948 31024 28960
rect 30979 28920 31024 28948
rect 31018 28908 31024 28920
rect 31076 28908 31082 28960
rect 1104 28858 32016 28880
rect 1104 28806 2136 28858
rect 2188 28806 12440 28858
rect 12492 28806 22744 28858
rect 22796 28806 32016 28858
rect 1104 28784 32016 28806
rect 4157 28747 4215 28753
rect 4157 28713 4169 28747
rect 4203 28744 4215 28747
rect 4522 28744 4528 28756
rect 4203 28716 4528 28744
rect 4203 28713 4215 28716
rect 4157 28707 4215 28713
rect 4522 28704 4528 28716
rect 4580 28704 4586 28756
rect 6917 28747 6975 28753
rect 6917 28713 6929 28747
rect 6963 28744 6975 28747
rect 8202 28744 8208 28756
rect 6963 28716 8208 28744
rect 6963 28713 6975 28716
rect 6917 28707 6975 28713
rect 8202 28704 8208 28716
rect 8260 28704 8266 28756
rect 8938 28744 8944 28756
rect 8899 28716 8944 28744
rect 8938 28704 8944 28716
rect 8996 28704 9002 28756
rect 10042 28744 10048 28756
rect 10003 28716 10048 28744
rect 10042 28704 10048 28716
rect 10100 28704 10106 28756
rect 11146 28744 11152 28756
rect 11107 28716 11152 28744
rect 11146 28704 11152 28716
rect 11204 28704 11210 28756
rect 11514 28744 11520 28756
rect 11475 28716 11520 28744
rect 11514 28704 11520 28716
rect 11572 28704 11578 28756
rect 12066 28744 12072 28756
rect 12027 28716 12072 28744
rect 12066 28704 12072 28716
rect 12124 28704 12130 28756
rect 12342 28704 12348 28756
rect 12400 28744 12406 28756
rect 12618 28744 12624 28756
rect 12400 28716 12624 28744
rect 12400 28704 12406 28716
rect 12618 28704 12624 28716
rect 12676 28704 12682 28756
rect 13265 28747 13323 28753
rect 13265 28713 13277 28747
rect 13311 28744 13323 28747
rect 14458 28744 14464 28756
rect 13311 28716 14464 28744
rect 13311 28713 13323 28716
rect 13265 28707 13323 28713
rect 14458 28704 14464 28716
rect 14516 28704 14522 28756
rect 14826 28704 14832 28756
rect 14884 28744 14890 28756
rect 15565 28747 15623 28753
rect 14884 28716 15332 28744
rect 14884 28704 14890 28716
rect 3050 28636 3056 28688
rect 3108 28676 3114 28688
rect 3237 28679 3295 28685
rect 3237 28676 3249 28679
rect 3108 28648 3249 28676
rect 3108 28636 3114 28648
rect 3237 28645 3249 28648
rect 3283 28676 3295 28679
rect 3786 28676 3792 28688
rect 3283 28648 3792 28676
rect 3283 28645 3295 28648
rect 3237 28639 3295 28645
rect 3786 28636 3792 28648
rect 3844 28676 3850 28688
rect 6365 28679 6423 28685
rect 6365 28676 6377 28679
rect 3844 28648 6377 28676
rect 3844 28636 3850 28648
rect 6365 28645 6377 28648
rect 6411 28645 6423 28679
rect 6365 28639 6423 28645
rect 7926 28636 7932 28688
rect 7984 28676 7990 28688
rect 7984 28648 8524 28676
rect 7984 28636 7990 28648
rect 4430 28568 4436 28620
rect 4488 28608 4494 28620
rect 4525 28611 4583 28617
rect 4525 28608 4537 28611
rect 4488 28580 4537 28608
rect 4488 28568 4494 28580
rect 4525 28577 4537 28580
rect 4571 28577 4583 28611
rect 5350 28608 5356 28620
rect 4525 28571 4583 28577
rect 4632 28580 5212 28608
rect 5311 28580 5356 28608
rect 1394 28500 1400 28552
rect 1452 28540 1458 28552
rect 1857 28543 1915 28549
rect 1857 28540 1869 28543
rect 1452 28512 1869 28540
rect 1452 28500 1458 28512
rect 1857 28509 1869 28512
rect 1903 28540 1915 28543
rect 2682 28540 2688 28552
rect 1903 28512 2688 28540
rect 1903 28509 1915 28512
rect 1857 28503 1915 28509
rect 2682 28500 2688 28512
rect 2740 28500 2746 28552
rect 4338 28540 4344 28552
rect 4299 28512 4344 28540
rect 4338 28500 4344 28512
rect 4396 28500 4402 28552
rect 4632 28549 4660 28580
rect 4617 28543 4675 28549
rect 4617 28509 4629 28543
rect 4663 28509 4675 28543
rect 4617 28503 4675 28509
rect 5077 28543 5135 28549
rect 5077 28509 5089 28543
rect 5123 28509 5135 28543
rect 5184 28540 5212 28580
rect 5350 28568 5356 28580
rect 5408 28568 5414 28620
rect 8110 28608 8116 28620
rect 6288 28580 8116 28608
rect 6288 28540 6316 28580
rect 8110 28568 8116 28580
rect 8168 28608 8174 28620
rect 8168 28580 8432 28608
rect 8168 28568 8174 28580
rect 5184 28512 6316 28540
rect 5077 28503 5135 28509
rect 2124 28475 2182 28481
rect 2124 28441 2136 28475
rect 2170 28472 2182 28475
rect 2222 28472 2228 28484
rect 2170 28444 2228 28472
rect 2170 28441 2182 28444
rect 2124 28435 2182 28441
rect 2222 28432 2228 28444
rect 2280 28432 2286 28484
rect 5092 28404 5120 28503
rect 6362 28500 6368 28552
rect 6420 28540 6426 28552
rect 6549 28543 6607 28549
rect 6549 28540 6561 28543
rect 6420 28512 6561 28540
rect 6420 28500 6426 28512
rect 6549 28509 6561 28512
rect 6595 28509 6607 28543
rect 6549 28503 6607 28509
rect 6638 28500 6644 28552
rect 6696 28540 6702 28552
rect 7926 28540 7932 28552
rect 6696 28512 6741 28540
rect 7887 28512 7932 28540
rect 6696 28500 6702 28512
rect 7926 28500 7932 28512
rect 7984 28500 7990 28552
rect 8202 28540 8208 28552
rect 8163 28512 8208 28540
rect 8202 28500 8208 28512
rect 8260 28500 8266 28552
rect 8404 28549 8432 28580
rect 8389 28543 8447 28549
rect 8389 28509 8401 28543
rect 8435 28509 8447 28543
rect 8496 28540 8524 28648
rect 9582 28636 9588 28688
rect 9640 28676 9646 28688
rect 9766 28676 9772 28688
rect 9640 28648 9772 28676
rect 9640 28636 9646 28648
rect 9766 28636 9772 28648
rect 9824 28636 9830 28688
rect 10962 28636 10968 28688
rect 11020 28676 11026 28688
rect 15194 28676 15200 28688
rect 11020 28648 15200 28676
rect 11020 28636 11026 28648
rect 15194 28636 15200 28648
rect 15252 28636 15258 28688
rect 15304 28676 15332 28716
rect 15565 28713 15577 28747
rect 15611 28744 15623 28747
rect 15746 28744 15752 28756
rect 15611 28716 15752 28744
rect 15611 28713 15623 28716
rect 15565 28707 15623 28713
rect 15746 28704 15752 28716
rect 15804 28704 15810 28756
rect 17865 28747 17923 28753
rect 15856 28716 17540 28744
rect 15856 28676 15884 28716
rect 15304 28648 15884 28676
rect 8754 28568 8760 28620
rect 8812 28608 8818 28620
rect 11146 28608 11152 28620
rect 8812 28580 9536 28608
rect 8812 28568 8818 28580
rect 9125 28543 9183 28549
rect 9125 28540 9137 28543
rect 8496 28512 9137 28540
rect 8389 28503 8447 28509
rect 9125 28509 9137 28512
rect 9171 28509 9183 28543
rect 9125 28503 9183 28509
rect 6178 28432 6184 28484
rect 6236 28472 6242 28484
rect 6733 28475 6791 28481
rect 6733 28472 6745 28475
rect 6236 28444 6745 28472
rect 6236 28432 6242 28444
rect 6733 28441 6745 28444
rect 6779 28441 6791 28475
rect 8404 28472 8432 28503
rect 9214 28500 9220 28552
rect 9272 28540 9278 28552
rect 9398 28540 9404 28552
rect 9272 28512 9317 28540
rect 9359 28512 9404 28540
rect 9272 28500 9278 28512
rect 9398 28500 9404 28512
rect 9456 28500 9462 28552
rect 9508 28549 9536 28580
rect 10704 28580 11152 28608
rect 9493 28543 9551 28549
rect 9493 28509 9505 28543
rect 9539 28509 9551 28543
rect 9493 28503 9551 28509
rect 9674 28500 9680 28552
rect 9732 28540 9738 28552
rect 10229 28543 10287 28549
rect 10229 28540 10241 28543
rect 9732 28512 10241 28540
rect 9732 28500 9738 28512
rect 10229 28509 10241 28512
rect 10275 28509 10287 28543
rect 10502 28540 10508 28552
rect 10463 28512 10508 28540
rect 10229 28503 10287 28509
rect 10502 28500 10508 28512
rect 10560 28500 10566 28552
rect 10704 28549 10732 28580
rect 11146 28568 11152 28580
rect 11204 28608 11210 28620
rect 11609 28611 11667 28617
rect 11609 28608 11621 28611
rect 11204 28580 11621 28608
rect 11204 28568 11210 28580
rect 11609 28577 11621 28580
rect 11655 28577 11667 28611
rect 11609 28571 11667 28577
rect 12406 28580 14320 28608
rect 10689 28543 10747 28549
rect 10689 28509 10701 28543
rect 10735 28509 10747 28543
rect 10689 28503 10747 28509
rect 10781 28543 10839 28549
rect 10781 28509 10793 28543
rect 10827 28540 10839 28543
rect 11333 28543 11391 28549
rect 11333 28540 11345 28543
rect 10827 28512 11345 28540
rect 10827 28509 10839 28512
rect 10781 28503 10839 28509
rect 11333 28509 11345 28512
rect 11379 28509 11391 28543
rect 11974 28540 11980 28552
rect 11333 28503 11391 28509
rect 11440 28512 11980 28540
rect 11440 28472 11468 28512
rect 11974 28500 11980 28512
rect 12032 28500 12038 28552
rect 12066 28500 12072 28552
rect 12124 28540 12130 28552
rect 12253 28543 12311 28549
rect 12253 28540 12265 28543
rect 12124 28512 12265 28540
rect 12124 28500 12130 28512
rect 12253 28509 12265 28512
rect 12299 28540 12311 28543
rect 12406 28540 12434 28580
rect 12526 28540 12532 28552
rect 12299 28512 12434 28540
rect 12487 28512 12532 28540
rect 12299 28509 12311 28512
rect 12253 28503 12311 28509
rect 12526 28500 12532 28512
rect 12584 28500 12590 28552
rect 12713 28543 12771 28549
rect 12713 28509 12725 28543
rect 12759 28509 12771 28543
rect 12713 28503 12771 28509
rect 6733 28435 6791 28441
rect 7300 28444 8340 28472
rect 8404 28444 11468 28472
rect 7300 28404 7328 28444
rect 5092 28376 7328 28404
rect 7374 28364 7380 28416
rect 7432 28404 7438 28416
rect 7745 28407 7803 28413
rect 7745 28404 7757 28407
rect 7432 28376 7757 28404
rect 7432 28364 7438 28376
rect 7745 28373 7757 28376
rect 7791 28373 7803 28407
rect 8312 28404 8340 28444
rect 11882 28432 11888 28484
rect 11940 28472 11946 28484
rect 12728 28472 12756 28503
rect 12802 28500 12808 28552
rect 12860 28540 12866 28552
rect 14292 28549 14320 28580
rect 13541 28543 13599 28549
rect 13541 28540 13553 28543
rect 12860 28512 13553 28540
rect 12860 28500 12866 28512
rect 13541 28509 13553 28512
rect 13587 28540 13599 28543
rect 14277 28543 14335 28549
rect 13587 28512 14228 28540
rect 13587 28509 13599 28512
rect 13541 28503 13599 28509
rect 11940 28444 12756 28472
rect 11940 28432 11946 28444
rect 13170 28432 13176 28484
rect 13228 28472 13234 28484
rect 13265 28475 13323 28481
rect 13265 28472 13277 28475
rect 13228 28444 13277 28472
rect 13228 28432 13234 28444
rect 13265 28441 13277 28444
rect 13311 28441 13323 28475
rect 13906 28472 13912 28484
rect 13265 28435 13323 28441
rect 13464 28444 13912 28472
rect 9490 28404 9496 28416
rect 8312 28376 9496 28404
rect 7745 28367 7803 28373
rect 9490 28364 9496 28376
rect 9548 28364 9554 28416
rect 9674 28364 9680 28416
rect 9732 28404 9738 28416
rect 10781 28407 10839 28413
rect 10781 28404 10793 28407
rect 9732 28376 10793 28404
rect 9732 28364 9738 28376
rect 10781 28373 10793 28376
rect 10827 28373 10839 28407
rect 10781 28367 10839 28373
rect 11054 28364 11060 28416
rect 11112 28404 11118 28416
rect 11698 28404 11704 28416
rect 11112 28376 11704 28404
rect 11112 28364 11118 28376
rect 11698 28364 11704 28376
rect 11756 28364 11762 28416
rect 12158 28364 12164 28416
rect 12216 28404 12222 28416
rect 13188 28404 13216 28432
rect 13464 28413 13492 28444
rect 13906 28432 13912 28444
rect 13964 28432 13970 28484
rect 12216 28376 13216 28404
rect 13449 28407 13507 28413
rect 12216 28364 12222 28376
rect 13449 28373 13461 28407
rect 13495 28373 13507 28407
rect 13449 28367 13507 28373
rect 13722 28364 13728 28416
rect 13780 28404 13786 28416
rect 14093 28407 14151 28413
rect 14093 28404 14105 28407
rect 13780 28376 14105 28404
rect 13780 28364 13786 28376
rect 14093 28373 14105 28376
rect 14139 28373 14151 28407
rect 14200 28404 14228 28512
rect 14277 28509 14289 28543
rect 14323 28509 14335 28543
rect 14277 28503 14335 28509
rect 14366 28500 14372 28552
rect 14424 28540 14430 28552
rect 14553 28543 14611 28549
rect 14553 28540 14565 28543
rect 14424 28512 14565 28540
rect 14424 28500 14430 28512
rect 14553 28509 14565 28512
rect 14599 28509 14611 28543
rect 14553 28503 14611 28509
rect 14642 28500 14648 28552
rect 14700 28540 14706 28552
rect 14737 28543 14795 28549
rect 14737 28540 14749 28543
rect 14700 28512 14749 28540
rect 14700 28500 14706 28512
rect 14737 28509 14749 28512
rect 14783 28509 14795 28543
rect 15212 28540 15240 28636
rect 17512 28608 17540 28716
rect 17865 28713 17877 28747
rect 17911 28744 17923 28747
rect 18322 28744 18328 28756
rect 17911 28716 18328 28744
rect 17911 28713 17923 28716
rect 17865 28707 17923 28713
rect 18322 28704 18328 28716
rect 18380 28704 18386 28756
rect 20625 28747 20683 28753
rect 20625 28713 20637 28747
rect 20671 28744 20683 28747
rect 20714 28744 20720 28756
rect 20671 28716 20720 28744
rect 20671 28713 20683 28716
rect 20625 28707 20683 28713
rect 20714 28704 20720 28716
rect 20772 28744 20778 28756
rect 21453 28747 21511 28753
rect 21453 28744 21465 28747
rect 20772 28716 21465 28744
rect 20772 28704 20778 28716
rect 21453 28713 21465 28716
rect 21499 28744 21511 28747
rect 21542 28744 21548 28756
rect 21499 28716 21548 28744
rect 21499 28713 21511 28716
rect 21453 28707 21511 28713
rect 21542 28704 21548 28716
rect 21600 28704 21606 28756
rect 21729 28747 21787 28753
rect 21729 28713 21741 28747
rect 21775 28744 21787 28747
rect 22370 28744 22376 28756
rect 21775 28716 22376 28744
rect 21775 28713 21787 28716
rect 21729 28707 21787 28713
rect 22370 28704 22376 28716
rect 22428 28704 22434 28756
rect 22649 28747 22707 28753
rect 22649 28713 22661 28747
rect 22695 28744 22707 28747
rect 23106 28744 23112 28756
rect 22695 28716 23112 28744
rect 22695 28713 22707 28716
rect 22649 28707 22707 28713
rect 23106 28704 23112 28716
rect 23164 28704 23170 28756
rect 25498 28704 25504 28756
rect 25556 28744 25562 28756
rect 25961 28747 26019 28753
rect 25961 28744 25973 28747
rect 25556 28716 25973 28744
rect 25556 28704 25562 28716
rect 25961 28713 25973 28716
rect 26007 28713 26019 28747
rect 26878 28744 26884 28756
rect 26839 28716 26884 28744
rect 25961 28707 26019 28713
rect 26878 28704 26884 28716
rect 26936 28704 26942 28756
rect 28994 28744 29000 28756
rect 27633 28716 28580 28744
rect 28955 28716 29000 28744
rect 18690 28676 18696 28688
rect 18651 28648 18696 28676
rect 18690 28636 18696 28648
rect 18748 28636 18754 28688
rect 20254 28636 20260 28688
rect 20312 28676 20318 28688
rect 20312 28648 22591 28676
rect 20312 28636 20318 28648
rect 17512 28580 19380 28608
rect 15746 28540 15752 28552
rect 15212 28512 15752 28540
rect 14737 28503 14795 28509
rect 14752 28472 14780 28503
rect 15746 28500 15752 28512
rect 15804 28500 15810 28552
rect 16025 28543 16083 28549
rect 16025 28509 16037 28543
rect 16071 28540 16083 28543
rect 16298 28540 16304 28552
rect 16071 28512 16304 28540
rect 16071 28509 16083 28512
rect 16025 28503 16083 28509
rect 16298 28500 16304 28512
rect 16356 28500 16362 28552
rect 16485 28543 16543 28549
rect 16485 28509 16497 28543
rect 16531 28540 16543 28543
rect 17310 28540 17316 28552
rect 16531 28512 17316 28540
rect 16531 28509 16543 28512
rect 16485 28503 16543 28509
rect 17310 28500 17316 28512
rect 17368 28540 17374 28552
rect 18046 28540 18052 28552
rect 17368 28512 18052 28540
rect 17368 28500 17374 28512
rect 18046 28500 18052 28512
rect 18104 28540 18110 28552
rect 19242 28540 19248 28552
rect 18104 28512 19248 28540
rect 18104 28500 18110 28512
rect 19242 28500 19248 28512
rect 19300 28500 19306 28552
rect 19352 28540 19380 28580
rect 21910 28568 21916 28620
rect 21968 28608 21974 28620
rect 22462 28608 22468 28620
rect 21968 28580 22468 28608
rect 21968 28568 21974 28580
rect 22462 28568 22468 28580
rect 22520 28568 22526 28620
rect 22563 28608 22591 28648
rect 22922 28636 22928 28688
rect 22980 28676 22986 28688
rect 22980 28648 23336 28676
rect 22980 28636 22986 28648
rect 22563 28580 23060 28608
rect 19501 28543 19559 28549
rect 19501 28540 19513 28543
rect 19352 28512 19513 28540
rect 19501 28509 19513 28512
rect 19547 28509 19559 28543
rect 19501 28503 19559 28509
rect 21085 28543 21143 28549
rect 21085 28509 21097 28543
rect 21131 28540 21143 28543
rect 21174 28540 21180 28552
rect 21131 28512 21180 28540
rect 21131 28509 21143 28512
rect 21085 28503 21143 28509
rect 21174 28500 21180 28512
rect 21232 28500 21238 28552
rect 21729 28543 21787 28549
rect 21729 28540 21741 28543
rect 21284 28512 21741 28540
rect 16758 28481 16764 28484
rect 15933 28475 15991 28481
rect 15933 28472 15945 28475
rect 14752 28444 15945 28472
rect 15933 28441 15945 28444
rect 15979 28441 15991 28475
rect 15933 28435 15991 28441
rect 16752 28435 16764 28481
rect 16816 28472 16822 28484
rect 16816 28444 16852 28472
rect 16758 28432 16764 28435
rect 16816 28432 16822 28444
rect 18506 28432 18512 28484
rect 18564 28472 18570 28484
rect 18564 28444 18609 28472
rect 18564 28432 18570 28444
rect 20162 28432 20168 28484
rect 20220 28472 20226 28484
rect 21284 28472 21312 28512
rect 21729 28509 21741 28512
rect 21775 28509 21787 28543
rect 21729 28503 21787 28509
rect 22646 28500 22652 28552
rect 22704 28540 22710 28552
rect 23032 28549 23060 28580
rect 23308 28549 23336 28648
rect 24302 28636 24308 28688
rect 24360 28676 24366 28688
rect 25314 28676 25320 28688
rect 24360 28648 25320 28676
rect 24360 28636 24366 28648
rect 25314 28636 25320 28648
rect 25372 28636 25378 28688
rect 25682 28636 25688 28688
rect 25740 28676 25746 28688
rect 27633 28676 27661 28716
rect 25740 28648 27661 28676
rect 28552 28676 28580 28716
rect 28994 28704 29000 28716
rect 29052 28744 29058 28756
rect 29730 28744 29736 28756
rect 29052 28716 29736 28744
rect 29052 28704 29058 28716
rect 29730 28704 29736 28716
rect 29788 28744 29794 28756
rect 30190 28744 30196 28756
rect 29788 28716 30196 28744
rect 29788 28704 29794 28716
rect 30190 28704 30196 28716
rect 30248 28704 30254 28756
rect 29086 28676 29092 28688
rect 28552 28648 29092 28676
rect 25740 28636 25746 28648
rect 29086 28636 29092 28648
rect 29144 28636 29150 28688
rect 24210 28568 24216 28620
rect 24268 28608 24274 28620
rect 24762 28608 24768 28620
rect 24268 28580 24532 28608
rect 24723 28580 24768 28608
rect 24268 28568 24274 28580
rect 22925 28543 22983 28549
rect 22925 28540 22937 28543
rect 22704 28512 22937 28540
rect 22704 28500 22710 28512
rect 22925 28509 22937 28512
rect 22971 28509 22983 28543
rect 22925 28503 22983 28509
rect 23017 28543 23075 28549
rect 23017 28509 23029 28543
rect 23063 28509 23075 28543
rect 23130 28543 23188 28549
rect 23130 28540 23142 28543
rect 23017 28503 23075 28509
rect 23113 28509 23142 28540
rect 23176 28509 23188 28543
rect 23113 28503 23188 28509
rect 23293 28543 23351 28549
rect 23293 28509 23305 28543
rect 23339 28509 23351 28543
rect 23293 28503 23351 28509
rect 20220 28444 21312 28472
rect 21453 28475 21511 28481
rect 20220 28432 20226 28444
rect 21453 28441 21465 28475
rect 21499 28441 21511 28475
rect 22373 28475 22431 28481
rect 22373 28472 22385 28475
rect 21453 28435 21511 28441
rect 21652 28444 22385 28472
rect 14826 28404 14832 28416
rect 14200 28376 14832 28404
rect 14093 28367 14151 28373
rect 14826 28364 14832 28376
rect 14884 28404 14890 28416
rect 21468 28404 21496 28435
rect 21652 28413 21680 28444
rect 22373 28441 22385 28444
rect 22419 28441 22431 28475
rect 22373 28435 22431 28441
rect 22830 28432 22836 28484
rect 22888 28472 22894 28484
rect 23113 28472 23141 28503
rect 23842 28500 23848 28552
rect 23900 28540 23906 28552
rect 24397 28543 24455 28549
rect 23900 28538 24348 28540
rect 24397 28538 24409 28543
rect 23900 28512 24409 28538
rect 23900 28500 23906 28512
rect 24320 28510 24409 28512
rect 24397 28509 24409 28510
rect 24443 28509 24455 28543
rect 24504 28542 24532 28580
rect 24762 28568 24768 28580
rect 24820 28568 24826 28620
rect 27614 28608 27620 28620
rect 27575 28580 27620 28608
rect 27614 28568 27620 28580
rect 27672 28568 27678 28620
rect 24581 28543 24639 28549
rect 24581 28542 24593 28543
rect 24504 28514 24593 28542
rect 24397 28503 24455 28509
rect 24581 28509 24593 28514
rect 24627 28509 24639 28543
rect 24581 28503 24639 28509
rect 24673 28543 24731 28549
rect 24673 28509 24685 28543
rect 24719 28509 24731 28543
rect 24673 28503 24731 28509
rect 24949 28543 25007 28549
rect 24949 28509 24961 28543
rect 24995 28540 25007 28543
rect 25038 28540 25044 28552
rect 24995 28512 25044 28540
rect 24995 28509 25007 28512
rect 24949 28503 25007 28509
rect 22888 28444 23141 28472
rect 24688 28472 24716 28503
rect 25038 28500 25044 28512
rect 25096 28500 25102 28552
rect 25406 28500 25412 28552
rect 25464 28540 25470 28552
rect 25590 28540 25596 28552
rect 25464 28512 25596 28540
rect 25464 28500 25470 28512
rect 25590 28500 25596 28512
rect 25648 28500 25654 28552
rect 25774 28540 25780 28552
rect 25735 28512 25780 28540
rect 25774 28500 25780 28512
rect 25832 28500 25838 28552
rect 26142 28500 26148 28552
rect 26200 28540 26206 28552
rect 26513 28543 26571 28549
rect 26513 28540 26525 28543
rect 26200 28512 26525 28540
rect 26200 28500 26206 28512
rect 26513 28509 26525 28512
rect 26559 28509 26571 28543
rect 27632 28540 27660 28568
rect 29914 28540 29920 28552
rect 27632 28512 29920 28540
rect 26513 28503 26571 28509
rect 29914 28500 29920 28512
rect 29972 28500 29978 28552
rect 30006 28500 30012 28552
rect 30064 28540 30070 28552
rect 30173 28543 30231 28549
rect 30173 28540 30185 28543
rect 30064 28512 30185 28540
rect 30064 28500 30070 28512
rect 30173 28509 30185 28512
rect 30219 28509 30231 28543
rect 30173 28503 30231 28509
rect 25222 28472 25228 28484
rect 24688 28444 25228 28472
rect 22888 28432 22894 28444
rect 25222 28432 25228 28444
rect 25280 28432 25286 28484
rect 25958 28432 25964 28484
rect 26016 28472 26022 28484
rect 27884 28475 27942 28481
rect 26016 28444 27200 28472
rect 26016 28432 26022 28444
rect 14884 28376 21496 28404
rect 21637 28407 21695 28413
rect 14884 28364 14890 28376
rect 21637 28373 21649 28407
rect 21683 28373 21695 28407
rect 21637 28367 21695 28373
rect 22002 28364 22008 28416
rect 22060 28404 22066 28416
rect 22462 28404 22468 28416
rect 22060 28376 22468 28404
rect 22060 28364 22066 28376
rect 22462 28364 22468 28376
rect 22520 28364 22526 28416
rect 22557 28407 22615 28413
rect 22557 28373 22569 28407
rect 22603 28404 22615 28407
rect 24486 28404 24492 28416
rect 22603 28376 24492 28404
rect 22603 28373 22615 28376
rect 22557 28367 22615 28373
rect 24486 28364 24492 28376
rect 24544 28404 24550 28416
rect 24762 28404 24768 28416
rect 24544 28376 24768 28404
rect 24544 28364 24550 28376
rect 24762 28364 24768 28376
rect 24820 28364 24826 28416
rect 24854 28364 24860 28416
rect 24912 28404 24918 28416
rect 25133 28407 25191 28413
rect 25133 28404 25145 28407
rect 24912 28376 25145 28404
rect 24912 28364 24918 28376
rect 25133 28373 25145 28376
rect 25179 28373 25191 28407
rect 25133 28367 25191 28373
rect 26418 28364 26424 28416
rect 26476 28404 26482 28416
rect 26881 28407 26939 28413
rect 26881 28404 26893 28407
rect 26476 28376 26893 28404
rect 26476 28364 26482 28376
rect 26881 28373 26893 28376
rect 26927 28373 26939 28407
rect 27062 28404 27068 28416
rect 27023 28376 27068 28404
rect 26881 28367 26939 28373
rect 27062 28364 27068 28376
rect 27120 28364 27126 28416
rect 27172 28404 27200 28444
rect 27884 28441 27896 28475
rect 27930 28472 27942 28475
rect 28534 28472 28540 28484
rect 27930 28444 28540 28472
rect 27930 28441 27942 28444
rect 27884 28435 27942 28441
rect 28534 28432 28540 28444
rect 28592 28432 28598 28484
rect 28966 28444 32352 28472
rect 28966 28404 28994 28444
rect 27172 28376 28994 28404
rect 29178 28364 29184 28416
rect 29236 28404 29242 28416
rect 31110 28404 31116 28416
rect 29236 28376 31116 28404
rect 29236 28364 29242 28376
rect 31110 28364 31116 28376
rect 31168 28404 31174 28416
rect 31297 28407 31355 28413
rect 31297 28404 31309 28407
rect 31168 28376 31309 28404
rect 31168 28364 31174 28376
rect 31297 28373 31309 28376
rect 31343 28373 31355 28407
rect 31297 28367 31355 28373
rect 1104 28314 32016 28336
rect 1104 28262 7288 28314
rect 7340 28262 17592 28314
rect 17644 28262 27896 28314
rect 27948 28262 32016 28314
rect 32324 28268 32352 28444
rect 1104 28240 32016 28262
rect 32232 28240 32352 28268
rect 1946 28160 1952 28212
rect 2004 28200 2010 28212
rect 2406 28200 2412 28212
rect 2004 28172 2412 28200
rect 2004 28160 2010 28172
rect 2406 28160 2412 28172
rect 2464 28160 2470 28212
rect 8202 28160 8208 28212
rect 8260 28200 8266 28212
rect 8260 28172 8708 28200
rect 8260 28160 8266 28172
rect 0 28132 800 28146
rect 2961 28135 3019 28141
rect 0 28104 1440 28132
rect 0 28090 800 28104
rect 1412 28073 1440 28104
rect 2961 28101 2973 28135
rect 3007 28132 3019 28135
rect 7742 28132 7748 28144
rect 3007 28104 7748 28132
rect 3007 28101 3019 28104
rect 2961 28095 3019 28101
rect 7742 28092 7748 28104
rect 7800 28092 7806 28144
rect 1397 28067 1455 28073
rect 1397 28033 1409 28067
rect 1443 28033 1455 28067
rect 1397 28027 1455 28033
rect 2406 28024 2412 28076
rect 2464 28064 2470 28076
rect 2501 28067 2559 28073
rect 2501 28064 2513 28067
rect 2464 28036 2513 28064
rect 2464 28024 2470 28036
rect 2501 28033 2513 28036
rect 2547 28033 2559 28067
rect 2501 28027 2559 28033
rect 5353 28067 5411 28073
rect 5353 28033 5365 28067
rect 5399 28064 5411 28067
rect 5534 28064 5540 28076
rect 5399 28036 5540 28064
rect 5399 28033 5411 28036
rect 5353 28027 5411 28033
rect 5534 28024 5540 28036
rect 5592 28024 5598 28076
rect 6632 28067 6690 28073
rect 6632 28033 6644 28067
rect 6678 28064 6690 28067
rect 7190 28064 7196 28076
rect 6678 28036 7196 28064
rect 6678 28033 6690 28036
rect 6632 28027 6690 28033
rect 7190 28024 7196 28036
rect 7248 28024 7254 28076
rect 7926 28024 7932 28076
rect 7984 28064 7990 28076
rect 8680 28073 8708 28172
rect 9674 28160 9680 28212
rect 9732 28200 9738 28212
rect 11054 28200 11060 28212
rect 9732 28172 9777 28200
rect 9876 28172 11060 28200
rect 9732 28160 9738 28172
rect 8754 28092 8760 28144
rect 8812 28132 8818 28144
rect 9876 28132 9904 28172
rect 11054 28160 11060 28172
rect 11112 28160 11118 28212
rect 11606 28160 11612 28212
rect 11664 28200 11670 28212
rect 11974 28200 11980 28212
rect 11664 28172 11980 28200
rect 11664 28160 11670 28172
rect 11974 28160 11980 28172
rect 12032 28160 12038 28212
rect 12342 28160 12348 28212
rect 12400 28200 12406 28212
rect 12710 28200 12716 28212
rect 12400 28172 12716 28200
rect 12400 28160 12406 28172
rect 12710 28160 12716 28172
rect 12768 28160 12774 28212
rect 14642 28200 14648 28212
rect 12820 28172 14648 28200
rect 10502 28132 10508 28144
rect 8812 28104 9904 28132
rect 10152 28104 10508 28132
rect 8812 28092 8818 28104
rect 8389 28067 8447 28073
rect 8389 28064 8401 28067
rect 7984 28036 8401 28064
rect 7984 28024 7990 28036
rect 8389 28033 8401 28036
rect 8435 28064 8447 28067
rect 8665 28067 8723 28073
rect 8435 28036 8616 28064
rect 8435 28033 8447 28036
rect 8389 28027 8447 28033
rect 2314 27956 2320 28008
rect 2372 27996 2378 28008
rect 5442 27996 5448 28008
rect 2372 27968 5448 27996
rect 2372 27956 2378 27968
rect 5442 27956 5448 27968
rect 5500 27956 5506 28008
rect 5629 27999 5687 28005
rect 5629 27965 5641 27999
rect 5675 27996 5687 27999
rect 5718 27996 5724 28008
rect 5675 27968 5724 27996
rect 5675 27965 5687 27968
rect 5629 27959 5687 27965
rect 5718 27956 5724 27968
rect 5776 27956 5782 28008
rect 6362 27996 6368 28008
rect 6323 27968 6368 27996
rect 6362 27956 6368 27968
rect 6420 27956 6426 28008
rect 7466 27956 7472 28008
rect 7524 27996 7530 28008
rect 8478 27996 8484 28008
rect 7524 27968 8484 27996
rect 7524 27956 7530 27968
rect 8478 27956 8484 27968
rect 8536 27956 8542 28008
rect 4338 27888 4344 27940
rect 4396 27928 4402 27940
rect 5350 27928 5356 27940
rect 4396 27900 5356 27928
rect 4396 27888 4402 27900
rect 5350 27888 5356 27900
rect 5408 27928 5414 27940
rect 5537 27931 5595 27937
rect 5537 27928 5549 27931
rect 5408 27900 5549 27928
rect 5408 27888 5414 27900
rect 5537 27897 5549 27900
rect 5583 27897 5595 27931
rect 5537 27891 5595 27897
rect 7745 27931 7803 27937
rect 7745 27897 7757 27931
rect 7791 27928 7803 27931
rect 8110 27928 8116 27940
rect 7791 27900 8116 27928
rect 7791 27897 7803 27900
rect 7745 27891 7803 27897
rect 8110 27888 8116 27900
rect 8168 27888 8174 27940
rect 8588 27928 8616 28036
rect 8665 28033 8677 28067
rect 8711 28033 8723 28067
rect 8665 28027 8723 28033
rect 8849 28067 8907 28073
rect 8849 28033 8861 28067
rect 8895 28064 8907 28067
rect 8941 28067 8999 28073
rect 8941 28064 8953 28067
rect 8895 28036 8953 28064
rect 8895 28033 8907 28036
rect 8849 28027 8907 28033
rect 8941 28033 8953 28036
rect 8987 28033 8999 28067
rect 8941 28027 8999 28033
rect 8680 27996 8708 28027
rect 9766 28024 9772 28076
rect 9824 28064 9830 28076
rect 10152 28073 10180 28104
rect 10502 28092 10508 28104
rect 10560 28092 10566 28144
rect 12820 28132 12848 28172
rect 14642 28160 14648 28172
rect 14700 28200 14706 28212
rect 14921 28203 14979 28209
rect 14921 28200 14933 28203
rect 14700 28172 14933 28200
rect 14700 28160 14706 28172
rect 14921 28169 14933 28172
rect 14967 28200 14979 28203
rect 16117 28203 16175 28209
rect 14967 28172 15976 28200
rect 14967 28169 14979 28172
rect 14921 28163 14979 28169
rect 10796 28104 12848 28132
rect 13556 28104 15608 28132
rect 9861 28067 9919 28073
rect 9861 28064 9873 28067
rect 9824 28036 9873 28064
rect 9824 28024 9830 28036
rect 9861 28033 9873 28036
rect 9907 28033 9919 28067
rect 9861 28027 9919 28033
rect 10137 28067 10195 28073
rect 10137 28033 10149 28067
rect 10183 28033 10195 28067
rect 10137 28027 10195 28033
rect 10152 27996 10180 28027
rect 10226 28024 10232 28076
rect 10284 28064 10290 28076
rect 10796 28073 10824 28104
rect 10321 28067 10379 28073
rect 10321 28064 10333 28067
rect 10284 28036 10333 28064
rect 10284 28024 10290 28036
rect 10321 28033 10333 28036
rect 10367 28033 10379 28067
rect 10321 28027 10379 28033
rect 10781 28067 10839 28073
rect 10781 28033 10793 28067
rect 10827 28033 10839 28067
rect 10962 28064 10968 28076
rect 10923 28036 10968 28064
rect 10781 28027 10839 28033
rect 10962 28024 10968 28036
rect 11020 28024 11026 28076
rect 11606 28024 11612 28076
rect 11664 28064 11670 28076
rect 11957 28067 12015 28073
rect 11957 28064 11969 28067
rect 11664 28036 11969 28064
rect 11664 28024 11670 28036
rect 11957 28033 11969 28036
rect 12003 28033 12015 28067
rect 13556 28064 13584 28104
rect 11957 28027 12015 28033
rect 12728 28036 13584 28064
rect 8680 27968 10180 27996
rect 11514 27956 11520 28008
rect 11572 27996 11578 28008
rect 11701 27999 11759 28005
rect 11701 27996 11713 27999
rect 11572 27968 11713 27996
rect 11572 27956 11578 27968
rect 11701 27965 11713 27968
rect 11747 27965 11759 27999
rect 11701 27959 11759 27965
rect 9766 27928 9772 27940
rect 8588 27900 9772 27928
rect 9766 27888 9772 27900
rect 9824 27888 9830 27940
rect 1394 27820 1400 27872
rect 1452 27860 1458 27872
rect 1581 27863 1639 27869
rect 1581 27860 1593 27863
rect 1452 27832 1593 27860
rect 1452 27820 1458 27832
rect 1581 27829 1593 27832
rect 1627 27829 1639 27863
rect 2314 27860 2320 27872
rect 2275 27832 2320 27860
rect 1581 27823 1639 27829
rect 2314 27820 2320 27832
rect 2372 27820 2378 27872
rect 2682 27820 2688 27872
rect 2740 27860 2746 27872
rect 4246 27860 4252 27872
rect 2740 27832 4252 27860
rect 2740 27820 2746 27832
rect 4246 27820 4252 27832
rect 4304 27820 4310 27872
rect 5166 27860 5172 27872
rect 5127 27832 5172 27860
rect 5166 27820 5172 27832
rect 5224 27820 5230 27872
rect 7834 27820 7840 27872
rect 7892 27860 7898 27872
rect 8205 27863 8263 27869
rect 8205 27860 8217 27863
rect 7892 27832 8217 27860
rect 7892 27820 7898 27832
rect 8205 27829 8217 27832
rect 8251 27829 8263 27863
rect 8205 27823 8263 27829
rect 8386 27820 8392 27872
rect 8444 27860 8450 27872
rect 8941 27863 8999 27869
rect 8941 27860 8953 27863
rect 8444 27832 8953 27860
rect 8444 27820 8450 27832
rect 8941 27829 8953 27832
rect 8987 27829 8999 27863
rect 8941 27823 8999 27829
rect 10873 27863 10931 27869
rect 10873 27829 10885 27863
rect 10919 27860 10931 27863
rect 12728 27860 12756 28036
rect 13630 28024 13636 28076
rect 13688 28064 13694 28076
rect 13797 28067 13855 28073
rect 13797 28064 13809 28067
rect 13688 28036 13809 28064
rect 13688 28024 13694 28036
rect 13797 28033 13809 28036
rect 13843 28033 13855 28067
rect 13797 28027 13855 28033
rect 14090 28024 14096 28076
rect 14148 28064 14154 28076
rect 15378 28064 15384 28076
rect 14148 28036 15240 28064
rect 15339 28036 15384 28064
rect 14148 28024 14154 28036
rect 13541 27999 13599 28005
rect 13541 27965 13553 27999
rect 13587 27965 13599 27999
rect 13541 27959 13599 27965
rect 12802 27888 12808 27940
rect 12860 27928 12866 27940
rect 13446 27928 13452 27940
rect 12860 27900 13452 27928
rect 12860 27888 12866 27900
rect 13446 27888 13452 27900
rect 13504 27888 13510 27940
rect 13078 27860 13084 27872
rect 10919 27832 12756 27860
rect 13039 27832 13084 27860
rect 10919 27829 10931 27832
rect 10873 27823 10931 27829
rect 13078 27820 13084 27832
rect 13136 27820 13142 27872
rect 13556 27860 13584 27959
rect 15212 27928 15240 28036
rect 15378 28024 15384 28036
rect 15436 28024 15442 28076
rect 15580 28073 15608 28104
rect 15948 28073 15976 28172
rect 16117 28169 16129 28203
rect 16163 28200 16175 28203
rect 16206 28200 16212 28212
rect 16163 28172 16212 28200
rect 16163 28169 16175 28172
rect 16117 28163 16175 28169
rect 16206 28160 16212 28172
rect 16264 28160 16270 28212
rect 17126 28160 17132 28212
rect 17184 28200 17190 28212
rect 17221 28203 17279 28209
rect 17221 28200 17233 28203
rect 17184 28172 17233 28200
rect 17184 28160 17190 28172
rect 17221 28169 17233 28172
rect 17267 28169 17279 28203
rect 17954 28200 17960 28212
rect 17221 28163 17279 28169
rect 17512 28172 17960 28200
rect 17512 28141 17540 28172
rect 17954 28160 17960 28172
rect 18012 28200 18018 28212
rect 18012 28172 18552 28200
rect 18012 28160 18018 28172
rect 17497 28135 17555 28141
rect 17497 28101 17509 28135
rect 17543 28101 17555 28135
rect 17497 28095 17555 28101
rect 17589 28135 17647 28141
rect 17589 28101 17601 28135
rect 17635 28132 17647 28135
rect 18322 28132 18328 28144
rect 17635 28104 18328 28132
rect 17635 28101 17647 28104
rect 17589 28095 17647 28101
rect 18322 28092 18328 28104
rect 18380 28092 18386 28144
rect 18524 28141 18552 28172
rect 19334 28160 19340 28212
rect 19392 28200 19398 28212
rect 19613 28203 19671 28209
rect 19613 28200 19625 28203
rect 19392 28172 19625 28200
rect 19392 28160 19398 28172
rect 19613 28169 19625 28172
rect 19659 28169 19671 28203
rect 21637 28203 21695 28209
rect 21637 28200 21649 28203
rect 19613 28163 19671 28169
rect 20364 28172 21649 28200
rect 18509 28135 18567 28141
rect 18509 28101 18521 28135
rect 18555 28132 18567 28135
rect 18690 28132 18696 28144
rect 18555 28104 18696 28132
rect 18555 28101 18567 28104
rect 18509 28095 18567 28101
rect 18690 28092 18696 28104
rect 18748 28092 18754 28144
rect 19518 28092 19524 28144
rect 19576 28132 19582 28144
rect 20364 28132 20392 28172
rect 21637 28169 21649 28172
rect 21683 28169 21695 28203
rect 21637 28163 21695 28169
rect 22462 28160 22468 28212
rect 22520 28200 22526 28212
rect 23845 28203 23903 28209
rect 23845 28200 23857 28203
rect 22520 28172 23857 28200
rect 22520 28160 22526 28172
rect 23845 28169 23857 28172
rect 23891 28169 23903 28203
rect 24210 28200 24216 28212
rect 24171 28172 24216 28200
rect 23845 28163 23903 28169
rect 24210 28160 24216 28172
rect 24268 28160 24274 28212
rect 24302 28160 24308 28212
rect 24360 28200 24366 28212
rect 24578 28200 24584 28212
rect 24360 28172 24584 28200
rect 24360 28160 24366 28172
rect 24578 28160 24584 28172
rect 24636 28160 24642 28212
rect 24762 28160 24768 28212
rect 24820 28200 24826 28212
rect 24857 28203 24915 28209
rect 24857 28200 24869 28203
rect 24820 28172 24869 28200
rect 24820 28160 24826 28172
rect 24857 28169 24869 28172
rect 24903 28169 24915 28203
rect 25038 28200 25044 28212
rect 24857 28163 24915 28169
rect 24964 28172 25044 28200
rect 19576 28104 20392 28132
rect 20625 28135 20683 28141
rect 19576 28092 19582 28104
rect 20625 28101 20637 28135
rect 20671 28132 20683 28135
rect 24394 28132 24400 28144
rect 20671 28104 24400 28132
rect 20671 28101 20683 28104
rect 20625 28095 20683 28101
rect 24394 28092 24400 28104
rect 24452 28132 24458 28144
rect 24964 28132 24992 28172
rect 25038 28160 25044 28172
rect 25096 28160 25102 28212
rect 25222 28160 25228 28212
rect 25280 28200 25286 28212
rect 25869 28203 25927 28209
rect 25869 28200 25881 28203
rect 25280 28172 25881 28200
rect 25280 28160 25286 28172
rect 25869 28169 25881 28172
rect 25915 28169 25927 28203
rect 27525 28203 27583 28209
rect 27525 28200 27537 28203
rect 25869 28163 25927 28169
rect 27172 28172 27537 28200
rect 24452 28104 24992 28132
rect 24452 28092 24458 28104
rect 15565 28067 15623 28073
rect 15565 28033 15577 28067
rect 15611 28033 15623 28067
rect 15565 28027 15623 28033
rect 15657 28067 15715 28073
rect 15657 28033 15669 28067
rect 15703 28064 15715 28067
rect 15933 28067 15991 28073
rect 15703 28036 15884 28064
rect 15703 28033 15715 28036
rect 15657 28027 15715 28033
rect 15286 27956 15292 28008
rect 15344 27996 15350 28008
rect 15749 27999 15807 28005
rect 15749 27996 15761 27999
rect 15344 27968 15761 27996
rect 15344 27956 15350 27968
rect 15749 27965 15761 27968
rect 15795 27965 15807 27999
rect 15856 27996 15884 28036
rect 15933 28033 15945 28067
rect 15979 28033 15991 28067
rect 15933 28027 15991 28033
rect 16942 28024 16948 28076
rect 17000 28064 17006 28076
rect 17405 28067 17463 28073
rect 17405 28064 17417 28067
rect 17000 28036 17417 28064
rect 17000 28024 17006 28036
rect 17405 28033 17417 28036
rect 17451 28033 17463 28067
rect 17405 28027 17463 28033
rect 17681 28067 17739 28073
rect 17681 28033 17693 28067
rect 17727 28033 17739 28067
rect 17681 28027 17739 28033
rect 17865 28067 17923 28073
rect 17865 28033 17877 28067
rect 17911 28064 17923 28067
rect 18230 28064 18236 28076
rect 17911 28036 18236 28064
rect 17911 28033 17923 28036
rect 17865 28027 17923 28033
rect 16114 27996 16120 28008
rect 15856 27968 16120 27996
rect 15749 27959 15807 27965
rect 16114 27956 16120 27968
rect 16172 27956 16178 28008
rect 17696 27996 17724 28027
rect 18230 28024 18236 28036
rect 18288 28024 18294 28076
rect 18601 28067 18659 28073
rect 18601 28033 18613 28067
rect 18647 28064 18659 28067
rect 18966 28064 18972 28076
rect 18647 28036 18972 28064
rect 18647 28033 18659 28036
rect 18601 28027 18659 28033
rect 18966 28024 18972 28036
rect 19024 28024 19030 28076
rect 19705 28067 19763 28073
rect 19705 28033 19717 28067
rect 19751 28064 19763 28067
rect 20901 28067 20959 28073
rect 20901 28064 20913 28067
rect 19751 28036 20913 28064
rect 19751 28033 19763 28036
rect 19705 28027 19763 28033
rect 20901 28033 20913 28036
rect 20947 28033 20959 28067
rect 20901 28027 20959 28033
rect 20993 28067 21051 28073
rect 20993 28033 21005 28067
rect 21039 28033 21051 28067
rect 20993 28027 21051 28033
rect 18397 27999 18455 28005
rect 18397 27996 18409 27999
rect 17696 27968 18409 27996
rect 18397 27965 18409 27968
rect 18443 27965 18455 27999
rect 19794 27996 19800 28008
rect 19755 27968 19800 27996
rect 18397 27959 18455 27965
rect 19794 27956 19800 27968
rect 19852 27956 19858 28008
rect 19245 27931 19303 27937
rect 19245 27928 19257 27931
rect 15212 27900 19257 27928
rect 19245 27897 19257 27900
rect 19291 27897 19303 27931
rect 20916 27928 20944 28027
rect 21008 27996 21036 28027
rect 21082 28024 21088 28076
rect 21140 28064 21146 28076
rect 21269 28067 21327 28073
rect 21140 28036 21185 28064
rect 21140 28024 21146 28036
rect 21269 28033 21281 28067
rect 21315 28033 21327 28067
rect 21269 28027 21327 28033
rect 21637 28067 21695 28073
rect 21637 28033 21649 28067
rect 21683 28064 21695 28067
rect 21913 28067 21971 28073
rect 21913 28064 21925 28067
rect 21683 28036 21925 28064
rect 21683 28033 21695 28036
rect 21637 28027 21695 28033
rect 21913 28033 21925 28036
rect 21959 28033 21971 28067
rect 22554 28064 22560 28076
rect 22467 28036 22560 28064
rect 21913 28027 21971 28033
rect 21008 27968 21128 27996
rect 21100 27928 21128 27968
rect 21174 27956 21180 28008
rect 21232 27996 21238 28008
rect 21284 27996 21312 28027
rect 21232 27968 21312 27996
rect 21232 27956 21238 27968
rect 21542 27956 21548 28008
rect 21600 27996 21606 28008
rect 22480 27996 22508 28036
rect 22554 28024 22560 28036
rect 22612 28064 22618 28076
rect 22899 28067 22957 28073
rect 22899 28064 22911 28067
rect 22612 28036 22911 28064
rect 22612 28024 22618 28036
rect 22899 28033 22911 28036
rect 22945 28033 22957 28067
rect 23198 28064 23204 28076
rect 23159 28036 23204 28064
rect 22899 28027 22957 28033
rect 23198 28024 23204 28036
rect 23256 28024 23262 28076
rect 24578 28064 24584 28076
rect 24539 28036 24584 28064
rect 24578 28024 24584 28036
rect 24636 28024 24642 28076
rect 24670 28024 24676 28076
rect 24728 28064 24734 28076
rect 24949 28067 25007 28073
rect 24728 28036 24773 28064
rect 24728 28024 24734 28036
rect 24949 28033 24961 28067
rect 24995 28064 25007 28067
rect 25682 28064 25688 28076
rect 24995 28036 25688 28064
rect 24995 28033 25007 28036
rect 24949 28027 25007 28033
rect 25682 28024 25688 28036
rect 25740 28024 25746 28076
rect 25866 28024 25872 28076
rect 25924 28064 25930 28076
rect 26145 28067 26203 28073
rect 26145 28064 26157 28067
rect 25924 28036 26157 28064
rect 25924 28024 25930 28036
rect 26145 28033 26157 28036
rect 26191 28033 26203 28067
rect 26145 28027 26203 28033
rect 26329 28067 26387 28073
rect 26329 28033 26341 28067
rect 26375 28064 26387 28067
rect 27062 28064 27068 28076
rect 26375 28036 27068 28064
rect 26375 28033 26387 28036
rect 26329 28027 26387 28033
rect 27062 28024 27068 28036
rect 27120 28024 27126 28076
rect 27172 28073 27200 28172
rect 27525 28169 27537 28172
rect 27571 28169 27583 28203
rect 27525 28163 27583 28169
rect 27798 28160 27804 28212
rect 27856 28200 27862 28212
rect 27893 28203 27951 28209
rect 27893 28200 27905 28203
rect 27856 28172 27905 28200
rect 27856 28160 27862 28172
rect 27893 28169 27905 28172
rect 27939 28169 27951 28203
rect 27893 28163 27951 28169
rect 28261 28203 28319 28209
rect 28261 28169 28273 28203
rect 28307 28200 28319 28203
rect 28442 28200 28448 28212
rect 28307 28172 28448 28200
rect 28307 28169 28319 28172
rect 28261 28163 28319 28169
rect 28442 28160 28448 28172
rect 28500 28160 28506 28212
rect 28813 28203 28871 28209
rect 28813 28169 28825 28203
rect 28859 28200 28871 28203
rect 31202 28200 31208 28212
rect 28859 28172 31208 28200
rect 28859 28169 28871 28172
rect 28813 28163 28871 28169
rect 31202 28160 31208 28172
rect 31260 28160 31266 28212
rect 27338 28092 27344 28144
rect 27396 28132 27402 28144
rect 28166 28132 28172 28144
rect 27396 28104 28172 28132
rect 27396 28092 27402 28104
rect 28166 28092 28172 28104
rect 28224 28092 28230 28144
rect 28353 28135 28411 28141
rect 28353 28101 28365 28135
rect 28399 28132 28411 28135
rect 31018 28132 31024 28144
rect 28399 28104 31024 28132
rect 28399 28101 28411 28104
rect 28353 28095 28411 28101
rect 31018 28092 31024 28104
rect 31076 28092 31082 28144
rect 32232 28132 32260 28240
rect 32320 28132 33120 28146
rect 32232 28104 33120 28132
rect 32320 28090 33120 28104
rect 27157 28067 27215 28073
rect 28813 28067 28871 28073
rect 27157 28033 27169 28067
rect 27203 28033 27215 28067
rect 27157 28027 27215 28033
rect 28276 28064 28580 28067
rect 28813 28064 28825 28067
rect 28276 28039 28825 28064
rect 21600 27968 22508 27996
rect 21600 27956 21606 27968
rect 22646 27956 22652 28008
rect 22704 27996 22710 28008
rect 23017 27999 23075 28005
rect 23017 27996 23029 27999
rect 22704 27968 23029 27996
rect 22704 27956 22710 27968
rect 23017 27965 23029 27968
rect 23063 27965 23075 27999
rect 23017 27959 23075 27965
rect 23109 27999 23167 28005
rect 23109 27965 23121 27999
rect 23155 27996 23167 27999
rect 23382 27996 23388 28008
rect 23155 27968 23388 27996
rect 23155 27965 23167 27968
rect 23109 27959 23167 27965
rect 23382 27956 23388 27968
rect 23440 27956 23446 28008
rect 24118 27956 24124 28008
rect 24176 27996 24182 28008
rect 25774 27996 25780 28008
rect 24176 27968 25780 27996
rect 24176 27956 24182 27968
rect 25774 27956 25780 27968
rect 25832 27956 25838 28008
rect 26053 27999 26111 28005
rect 26053 27965 26065 27999
rect 26099 27965 26111 27999
rect 26053 27959 26111 27965
rect 21266 27928 21272 27940
rect 20916 27900 21036 27928
rect 21100 27900 21272 27928
rect 19245 27891 19303 27897
rect 14550 27860 14556 27872
rect 13556 27832 14556 27860
rect 14550 27820 14556 27832
rect 14608 27820 14614 27872
rect 16298 27820 16304 27872
rect 16356 27860 16362 27872
rect 18966 27860 18972 27872
rect 16356 27832 18972 27860
rect 16356 27820 16362 27832
rect 18966 27820 18972 27832
rect 19024 27820 19030 27872
rect 19058 27820 19064 27872
rect 19116 27860 19122 27872
rect 20070 27860 20076 27872
rect 19116 27832 20076 27860
rect 19116 27820 19122 27832
rect 20070 27820 20076 27832
rect 20128 27820 20134 27872
rect 21008 27860 21036 27900
rect 21266 27888 21272 27900
rect 21324 27888 21330 27940
rect 22097 27931 22155 27937
rect 22097 27897 22109 27931
rect 22143 27928 22155 27931
rect 22462 27928 22468 27940
rect 22143 27900 22468 27928
rect 22143 27897 22155 27900
rect 22097 27891 22155 27897
rect 22462 27888 22468 27900
rect 22520 27888 22526 27940
rect 22741 27931 22799 27937
rect 22741 27897 22753 27931
rect 22787 27928 22799 27931
rect 24946 27928 24952 27940
rect 22787 27900 24952 27928
rect 22787 27897 22799 27900
rect 22741 27891 22799 27897
rect 24946 27888 24952 27900
rect 25004 27888 25010 27940
rect 25590 27888 25596 27940
rect 25648 27928 25654 27940
rect 26068 27928 26096 27959
rect 26234 27956 26240 28008
rect 26292 27996 26298 28008
rect 27433 27999 27491 28005
rect 26292 27968 26337 27996
rect 26292 27956 26298 27968
rect 27433 27965 27445 27999
rect 27479 27996 27491 27999
rect 28276 27996 28304 28039
rect 28552 28036 28825 28039
rect 28813 28033 28825 28036
rect 28859 28033 28871 28067
rect 28813 28027 28871 28033
rect 29273 28067 29331 28073
rect 29273 28033 29285 28067
rect 29319 28033 29331 28067
rect 29273 28027 29331 28033
rect 29549 28067 29607 28073
rect 29549 28033 29561 28067
rect 29595 28033 29607 28067
rect 29730 28064 29736 28076
rect 29691 28036 29736 28064
rect 29549 28027 29607 28033
rect 27479 27968 28304 27996
rect 27479 27965 27491 27968
rect 27433 27959 27491 27965
rect 28442 27956 28448 28008
rect 28500 27996 28506 28008
rect 29288 27996 29316 28027
rect 28500 27968 28545 27996
rect 29288 27968 29500 27996
rect 28500 27956 28506 27968
rect 26878 27928 26884 27940
rect 25648 27900 26884 27928
rect 25648 27888 25654 27900
rect 26878 27888 26884 27900
rect 26936 27888 26942 27940
rect 26973 27931 27031 27937
rect 26973 27897 26985 27931
rect 27019 27928 27031 27931
rect 29270 27928 29276 27940
rect 27019 27900 29276 27928
rect 27019 27897 27031 27900
rect 26973 27891 27031 27897
rect 29270 27888 29276 27900
rect 29328 27888 29334 27940
rect 23750 27860 23756 27872
rect 21008 27832 23756 27860
rect 23750 27820 23756 27832
rect 23808 27820 23814 27872
rect 23845 27863 23903 27869
rect 23845 27829 23857 27863
rect 23891 27860 23903 27863
rect 24489 27863 24547 27869
rect 24489 27860 24501 27863
rect 23891 27832 24501 27860
rect 23891 27829 23903 27832
rect 23845 27823 23903 27829
rect 24489 27829 24501 27832
rect 24535 27860 24547 27863
rect 24578 27860 24584 27872
rect 24535 27832 24584 27860
rect 24535 27829 24547 27832
rect 24489 27823 24547 27829
rect 24578 27820 24584 27832
rect 24636 27820 24642 27872
rect 24670 27820 24676 27872
rect 24728 27860 24734 27872
rect 24854 27860 24860 27872
rect 24728 27832 24860 27860
rect 24728 27820 24734 27832
rect 24854 27820 24860 27832
rect 24912 27820 24918 27872
rect 27338 27860 27344 27872
rect 27299 27832 27344 27860
rect 27338 27820 27344 27832
rect 27396 27820 27402 27872
rect 27525 27863 27583 27869
rect 27525 27829 27537 27863
rect 27571 27860 27583 27863
rect 28626 27860 28632 27872
rect 27571 27832 28632 27860
rect 27571 27829 27583 27832
rect 27525 27823 27583 27829
rect 28626 27820 28632 27832
rect 28684 27820 28690 27872
rect 28718 27820 28724 27872
rect 28776 27860 28782 27872
rect 29089 27863 29147 27869
rect 29089 27860 29101 27863
rect 28776 27832 29101 27860
rect 28776 27820 28782 27832
rect 29089 27829 29101 27832
rect 29135 27829 29147 27863
rect 29472 27860 29500 27968
rect 29564 27928 29592 28027
rect 29730 28024 29736 28036
rect 29788 28024 29794 28076
rect 30193 28067 30251 28073
rect 30193 28033 30205 28067
rect 30239 28064 30251 28067
rect 30469 28067 30527 28073
rect 30469 28064 30481 28067
rect 30239 28036 30481 28064
rect 30239 28033 30251 28036
rect 30193 28027 30251 28033
rect 30469 28033 30481 28036
rect 30515 28064 30527 28067
rect 30650 28064 30656 28076
rect 30515 28036 30656 28064
rect 30515 28033 30527 28036
rect 30469 28027 30527 28033
rect 30650 28024 30656 28036
rect 30708 28024 30714 28076
rect 30742 28024 30748 28076
rect 30800 28064 30806 28076
rect 30800 28036 30893 28064
rect 30800 28024 30806 28036
rect 30926 28024 30932 28076
rect 30984 28064 30990 28076
rect 31294 28064 31300 28076
rect 30984 28036 31300 28064
rect 30984 28024 30990 28036
rect 31294 28024 31300 28036
rect 31352 28024 31358 28076
rect 30760 27928 30788 28024
rect 29564 27900 30788 27928
rect 30193 27863 30251 27869
rect 30193 27860 30205 27863
rect 29472 27832 30205 27860
rect 29089 27823 29147 27829
rect 30193 27829 30205 27832
rect 30239 27829 30251 27863
rect 30193 27823 30251 27829
rect 30285 27863 30343 27869
rect 30285 27829 30297 27863
rect 30331 27860 30343 27863
rect 30558 27860 30564 27872
rect 30331 27832 30564 27860
rect 30331 27829 30343 27832
rect 30285 27823 30343 27829
rect 30558 27820 30564 27832
rect 30616 27820 30622 27872
rect 1104 27770 32016 27792
rect 1104 27718 2136 27770
rect 2188 27718 12440 27770
rect 12492 27718 22744 27770
rect 22796 27718 32016 27770
rect 1104 27696 32016 27718
rect 4430 27656 4436 27668
rect 4172 27628 4436 27656
rect 2590 27588 2596 27600
rect 2551 27560 2596 27588
rect 2590 27548 2596 27560
rect 2648 27548 2654 27600
rect 2961 27591 3019 27597
rect 2961 27557 2973 27591
rect 3007 27588 3019 27591
rect 4172 27588 4200 27628
rect 4430 27616 4436 27628
rect 4488 27616 4494 27668
rect 7852 27628 8064 27656
rect 4338 27588 4344 27600
rect 3007 27560 4200 27588
rect 4299 27560 4344 27588
rect 3007 27557 3019 27560
rect 2961 27551 3019 27557
rect 4338 27548 4344 27560
rect 4396 27548 4402 27600
rect 6273 27591 6331 27597
rect 6273 27557 6285 27591
rect 6319 27588 6331 27591
rect 6914 27588 6920 27600
rect 6319 27560 6920 27588
rect 6319 27557 6331 27560
rect 6273 27551 6331 27557
rect 6914 27548 6920 27560
rect 6972 27548 6978 27600
rect 7193 27591 7251 27597
rect 7193 27557 7205 27591
rect 7239 27588 7251 27591
rect 7466 27588 7472 27600
rect 7239 27560 7472 27588
rect 7239 27557 7251 27560
rect 7193 27551 7251 27557
rect 7466 27548 7472 27560
rect 7524 27588 7530 27600
rect 7852 27588 7880 27628
rect 7524 27560 7880 27588
rect 8036 27588 8064 27628
rect 8478 27616 8484 27668
rect 8536 27656 8542 27668
rect 9122 27656 9128 27668
rect 8536 27628 9128 27656
rect 8536 27616 8542 27628
rect 9122 27616 9128 27628
rect 9180 27616 9186 27668
rect 11517 27659 11575 27665
rect 11517 27625 11529 27659
rect 11563 27656 11575 27659
rect 11606 27656 11612 27668
rect 11563 27628 11612 27656
rect 11563 27625 11575 27628
rect 11517 27619 11575 27625
rect 11606 27616 11612 27628
rect 11664 27616 11670 27668
rect 11790 27616 11796 27668
rect 11848 27656 11854 27668
rect 11848 27628 15700 27656
rect 11848 27616 11854 27628
rect 9309 27591 9367 27597
rect 9309 27588 9321 27591
rect 8036 27560 9321 27588
rect 7524 27548 7530 27560
rect 9309 27557 9321 27560
rect 9355 27588 9367 27591
rect 10410 27588 10416 27600
rect 9355 27560 10416 27588
rect 9355 27557 9367 27560
rect 9309 27551 9367 27557
rect 10410 27548 10416 27560
rect 10468 27548 10474 27600
rect 11885 27591 11943 27597
rect 11885 27557 11897 27591
rect 11931 27588 11943 27591
rect 13906 27588 13912 27600
rect 11931 27560 13912 27588
rect 11931 27557 11943 27560
rect 11885 27551 11943 27557
rect 13906 27548 13912 27560
rect 13964 27588 13970 27600
rect 14182 27588 14188 27600
rect 13964 27560 14188 27588
rect 13964 27548 13970 27560
rect 14182 27548 14188 27560
rect 14240 27548 14246 27600
rect 15672 27588 15700 27628
rect 15746 27616 15752 27668
rect 15804 27656 15810 27668
rect 16025 27659 16083 27665
rect 16025 27656 16037 27659
rect 15804 27628 16037 27656
rect 15804 27616 15810 27628
rect 16025 27625 16037 27628
rect 16071 27625 16083 27659
rect 20901 27659 20959 27665
rect 16025 27619 16083 27625
rect 16546 27628 19748 27656
rect 16546 27588 16574 27628
rect 19720 27588 19748 27628
rect 20901 27625 20913 27659
rect 20947 27656 20959 27659
rect 21082 27656 21088 27668
rect 20947 27628 21088 27656
rect 20947 27625 20959 27628
rect 20901 27619 20959 27625
rect 21082 27616 21088 27628
rect 21140 27616 21146 27668
rect 21453 27659 21511 27665
rect 21453 27625 21465 27659
rect 21499 27656 21511 27659
rect 23014 27656 23020 27668
rect 21499 27628 23020 27656
rect 21499 27625 21511 27628
rect 21453 27619 21511 27625
rect 23014 27616 23020 27628
rect 23072 27616 23078 27668
rect 23290 27616 23296 27668
rect 23348 27656 23354 27668
rect 23566 27656 23572 27668
rect 23348 27628 23572 27656
rect 23348 27616 23354 27628
rect 23566 27616 23572 27628
rect 23624 27616 23630 27668
rect 24486 27656 24492 27668
rect 24447 27628 24492 27656
rect 24486 27616 24492 27628
rect 24544 27616 24550 27668
rect 25866 27616 25872 27668
rect 25924 27656 25930 27668
rect 26145 27659 26203 27665
rect 26145 27656 26157 27659
rect 25924 27628 26157 27656
rect 25924 27616 25930 27628
rect 26145 27625 26157 27628
rect 26191 27625 26203 27659
rect 26145 27619 26203 27625
rect 26234 27616 26240 27668
rect 26292 27656 26298 27668
rect 27430 27656 27436 27668
rect 26292 27628 27436 27656
rect 26292 27616 26298 27628
rect 27430 27616 27436 27628
rect 27488 27656 27494 27668
rect 28534 27656 28540 27668
rect 27488 27628 27660 27656
rect 28495 27628 28540 27656
rect 27488 27616 27494 27628
rect 21266 27588 21272 27600
rect 15672 27560 16574 27588
rect 18340 27560 19656 27588
rect 19720 27560 21272 27588
rect 1578 27480 1584 27532
rect 1636 27520 1642 27532
rect 2041 27523 2099 27529
rect 2041 27520 2053 27523
rect 1636 27492 2053 27520
rect 1636 27480 1642 27492
rect 2041 27489 2053 27492
rect 2087 27489 2099 27523
rect 2041 27483 2099 27489
rect 2133 27523 2191 27529
rect 2133 27489 2145 27523
rect 2179 27520 2191 27523
rect 2866 27520 2872 27532
rect 2179 27492 2872 27520
rect 2179 27489 2191 27492
rect 2133 27483 2191 27489
rect 2866 27480 2872 27492
rect 2924 27480 2930 27532
rect 3050 27520 3056 27532
rect 3011 27492 3056 27520
rect 3050 27480 3056 27492
rect 3108 27480 3114 27532
rect 4246 27480 4252 27532
rect 4304 27520 4310 27532
rect 4893 27523 4951 27529
rect 4893 27520 4905 27523
rect 4304 27492 4905 27520
rect 4304 27480 4310 27492
rect 4893 27489 4905 27492
rect 4939 27489 4951 27523
rect 7834 27520 7840 27532
rect 4893 27483 4951 27489
rect 7024 27492 7840 27520
rect 1857 27455 1915 27461
rect 1857 27421 1869 27455
rect 1903 27452 1915 27455
rect 1903 27424 2728 27452
rect 1903 27421 1915 27424
rect 1857 27415 1915 27421
rect 2700 27384 2728 27424
rect 2774 27412 2780 27464
rect 2832 27452 2838 27464
rect 4154 27452 4160 27464
rect 2832 27424 2877 27452
rect 4115 27424 4160 27452
rect 2832 27412 2838 27424
rect 4154 27412 4160 27424
rect 4212 27412 4218 27464
rect 5166 27461 5172 27464
rect 4433 27455 4491 27461
rect 4433 27421 4445 27455
rect 4479 27421 4491 27455
rect 5160 27452 5172 27461
rect 5127 27424 5172 27452
rect 4433 27415 4491 27421
rect 5160 27415 5172 27424
rect 4338 27384 4344 27396
rect 2700 27356 4344 27384
rect 4338 27344 4344 27356
rect 4396 27344 4402 27396
rect 4448 27384 4476 27415
rect 5166 27412 5172 27415
rect 5224 27412 5230 27464
rect 7024 27461 7052 27492
rect 7834 27480 7840 27492
rect 7892 27480 7898 27532
rect 8481 27523 8539 27529
rect 8481 27520 8493 27523
rect 8391 27492 8493 27520
rect 7009 27455 7067 27461
rect 7009 27421 7021 27455
rect 7055 27421 7067 27455
rect 7009 27415 7067 27421
rect 7285 27455 7343 27461
rect 7285 27421 7297 27455
rect 7331 27421 7343 27455
rect 7285 27415 7343 27421
rect 5074 27384 5080 27396
rect 4448 27356 5080 27384
rect 5074 27344 5080 27356
rect 5132 27344 5138 27396
rect 1673 27319 1731 27325
rect 1673 27285 1685 27319
rect 1719 27316 1731 27319
rect 2774 27316 2780 27328
rect 1719 27288 2780 27316
rect 1719 27285 1731 27288
rect 1673 27279 1731 27285
rect 2774 27276 2780 27288
rect 2832 27276 2838 27328
rect 3973 27319 4031 27325
rect 3973 27285 3985 27319
rect 4019 27316 4031 27319
rect 4062 27316 4068 27328
rect 4019 27288 4068 27316
rect 4019 27285 4031 27288
rect 3973 27279 4031 27285
rect 4062 27276 4068 27288
rect 4120 27276 4126 27328
rect 6825 27319 6883 27325
rect 6825 27285 6837 27319
rect 6871 27316 6883 27319
rect 7006 27316 7012 27328
rect 6871 27288 7012 27316
rect 6871 27285 6883 27288
rect 6825 27279 6883 27285
rect 7006 27276 7012 27288
rect 7064 27276 7070 27328
rect 7300 27316 7328 27415
rect 7926 27412 7932 27464
rect 7984 27452 7990 27464
rect 8202 27452 8208 27464
rect 7984 27424 8029 27452
rect 8163 27424 8208 27452
rect 7984 27412 7990 27424
rect 8202 27412 8208 27424
rect 8260 27412 8266 27464
rect 8404 27461 8432 27492
rect 8481 27489 8493 27492
rect 8527 27520 8539 27523
rect 9214 27520 9220 27532
rect 8527 27492 9220 27520
rect 8527 27489 8539 27492
rect 8481 27483 8539 27489
rect 9214 27480 9220 27492
rect 9272 27480 9278 27532
rect 9401 27523 9459 27529
rect 9401 27489 9413 27523
rect 9447 27520 9459 27523
rect 10226 27520 10232 27532
rect 9447 27492 10232 27520
rect 9447 27489 9459 27492
rect 9401 27483 9459 27489
rect 10226 27480 10232 27492
rect 10284 27480 10290 27532
rect 12802 27520 12808 27532
rect 11624 27492 12808 27520
rect 8389 27455 8447 27461
rect 8389 27421 8401 27455
rect 8435 27421 8447 27455
rect 8389 27415 8447 27421
rect 9125 27455 9183 27461
rect 9125 27421 9137 27455
rect 9171 27421 9183 27455
rect 9125 27415 9183 27421
rect 7745 27387 7803 27393
rect 7745 27353 7757 27387
rect 7791 27384 7803 27387
rect 9140 27384 9168 27415
rect 9490 27412 9496 27464
rect 9548 27452 9554 27464
rect 9861 27455 9919 27461
rect 9861 27452 9873 27455
rect 9548 27424 9873 27452
rect 9548 27412 9554 27424
rect 9861 27421 9873 27424
rect 9907 27421 9919 27455
rect 9861 27415 9919 27421
rect 10137 27455 10195 27461
rect 10137 27421 10149 27455
rect 10183 27452 10195 27455
rect 10502 27452 10508 27464
rect 10183 27424 10508 27452
rect 10183 27421 10195 27424
rect 10137 27415 10195 27421
rect 7791 27356 9168 27384
rect 9876 27384 9904 27415
rect 10502 27412 10508 27424
rect 10560 27412 10566 27464
rect 11624 27384 11652 27492
rect 12802 27480 12808 27492
rect 12860 27480 12866 27532
rect 14366 27520 14372 27532
rect 12912 27492 14372 27520
rect 12912 27464 12940 27492
rect 14366 27480 14372 27492
rect 14424 27480 14430 27532
rect 11701 27455 11759 27461
rect 11701 27421 11713 27455
rect 11747 27421 11759 27455
rect 11701 27415 11759 27421
rect 9876 27356 11652 27384
rect 11716 27384 11744 27415
rect 11882 27412 11888 27464
rect 11940 27452 11946 27464
rect 11977 27455 12035 27461
rect 11977 27452 11989 27455
rect 11940 27424 11989 27452
rect 11940 27412 11946 27424
rect 11977 27421 11989 27424
rect 12023 27421 12035 27455
rect 11977 27415 12035 27421
rect 12066 27412 12072 27464
rect 12124 27452 12130 27464
rect 12621 27455 12679 27461
rect 12621 27452 12633 27455
rect 12124 27424 12633 27452
rect 12124 27412 12130 27424
rect 12621 27421 12633 27424
rect 12667 27421 12679 27455
rect 12894 27452 12900 27464
rect 12855 27424 12900 27452
rect 12621 27415 12679 27421
rect 12894 27412 12900 27424
rect 12952 27412 12958 27464
rect 13078 27452 13084 27464
rect 13039 27424 13084 27452
rect 13078 27412 13084 27424
rect 13136 27412 13142 27464
rect 13170 27412 13176 27464
rect 13228 27452 13234 27464
rect 13998 27452 14004 27464
rect 13228 27424 14004 27452
rect 13228 27412 13234 27424
rect 13998 27412 14004 27424
rect 14056 27412 14062 27464
rect 14550 27412 14556 27464
rect 14608 27452 14614 27464
rect 14645 27455 14703 27461
rect 14645 27452 14657 27455
rect 14608 27424 14657 27452
rect 14608 27412 14614 27424
rect 14645 27421 14657 27424
rect 14691 27421 14703 27455
rect 14645 27415 14703 27421
rect 14734 27412 14740 27464
rect 14792 27452 14798 27464
rect 14901 27455 14959 27461
rect 14901 27452 14913 27455
rect 14792 27424 14913 27452
rect 14792 27412 14798 27424
rect 14901 27421 14913 27424
rect 14947 27421 14959 27455
rect 14901 27415 14959 27421
rect 15194 27412 15200 27464
rect 15252 27452 15258 27464
rect 16577 27455 16635 27461
rect 16577 27452 16589 27455
rect 15252 27424 16589 27452
rect 15252 27412 15258 27424
rect 16577 27421 16589 27424
rect 16623 27421 16635 27455
rect 17310 27452 17316 27464
rect 17271 27424 17316 27452
rect 16577 27415 16635 27421
rect 17310 27412 17316 27424
rect 17368 27412 17374 27464
rect 18340 27452 18368 27560
rect 18877 27523 18935 27529
rect 18877 27489 18889 27523
rect 18923 27520 18935 27523
rect 19058 27520 19064 27532
rect 18923 27492 19064 27520
rect 18923 27489 18935 27492
rect 18877 27483 18935 27489
rect 19058 27480 19064 27492
rect 19116 27480 19122 27532
rect 17512 27424 18368 27452
rect 12437 27387 12495 27393
rect 12437 27384 12449 27387
rect 11716 27356 12449 27384
rect 7791 27353 7803 27356
rect 7745 27347 7803 27353
rect 12437 27353 12449 27356
rect 12483 27353 12495 27387
rect 12437 27347 12495 27353
rect 12802 27344 12808 27396
rect 12860 27384 12866 27396
rect 13096 27384 13124 27412
rect 12860 27356 13124 27384
rect 12860 27344 12866 27356
rect 15102 27344 15108 27396
rect 15160 27384 15166 27396
rect 17512 27384 17540 27424
rect 18598 27412 18604 27464
rect 18656 27452 18662 27464
rect 19628 27461 19656 27560
rect 21266 27548 21272 27560
rect 21324 27548 21330 27600
rect 22005 27591 22063 27597
rect 22005 27557 22017 27591
rect 22051 27588 22063 27591
rect 22554 27588 22560 27600
rect 22051 27560 22560 27588
rect 22051 27557 22063 27560
rect 22005 27551 22063 27557
rect 22554 27548 22560 27560
rect 22612 27548 22618 27600
rect 23198 27548 23204 27600
rect 23256 27588 23262 27600
rect 24302 27588 24308 27600
rect 23256 27560 24308 27588
rect 23256 27548 23262 27560
rect 24302 27548 24308 27560
rect 24360 27548 24366 27600
rect 25501 27591 25559 27597
rect 25501 27557 25513 27591
rect 25547 27588 25559 27591
rect 25590 27588 25596 27600
rect 25547 27560 25596 27588
rect 25547 27557 25559 27560
rect 25501 27551 25559 27557
rect 25590 27548 25596 27560
rect 25648 27548 25654 27600
rect 27632 27588 27660 27628
rect 28534 27616 28540 27628
rect 28592 27616 28598 27668
rect 28626 27616 28632 27668
rect 28684 27656 28690 27668
rect 29822 27656 29828 27668
rect 28684 27628 29828 27656
rect 28684 27616 28690 27628
rect 29822 27616 29828 27628
rect 29880 27616 29886 27668
rect 31294 27656 31300 27668
rect 31255 27628 31300 27656
rect 31294 27616 31300 27628
rect 31352 27616 31358 27668
rect 28077 27591 28135 27597
rect 28077 27588 28089 27591
rect 27632 27560 28089 27588
rect 28077 27557 28089 27560
rect 28123 27557 28135 27591
rect 28077 27551 28135 27557
rect 22646 27480 22652 27532
rect 22704 27520 22710 27532
rect 23017 27523 23075 27529
rect 23017 27520 23029 27523
rect 22704 27492 23029 27520
rect 22704 27480 22710 27492
rect 23017 27489 23029 27492
rect 23063 27489 23075 27523
rect 23017 27483 23075 27489
rect 23842 27480 23848 27532
rect 23900 27520 23906 27532
rect 24673 27523 24731 27529
rect 24673 27520 24685 27523
rect 23900 27492 24685 27520
rect 23900 27480 23906 27492
rect 24673 27489 24685 27492
rect 24719 27520 24731 27523
rect 25682 27520 25688 27532
rect 24719 27492 25688 27520
rect 24719 27489 24731 27492
rect 24673 27483 24731 27489
rect 25682 27480 25688 27492
rect 25740 27480 25746 27532
rect 28997 27523 29055 27529
rect 28997 27489 29009 27523
rect 29043 27520 29055 27523
rect 29178 27520 29184 27532
rect 29043 27492 29184 27520
rect 29043 27489 29055 27492
rect 28997 27483 29055 27489
rect 29178 27480 29184 27492
rect 29236 27480 29242 27532
rect 29914 27520 29920 27532
rect 29875 27492 29920 27520
rect 29914 27480 29920 27492
rect 29972 27480 29978 27532
rect 19521 27455 19579 27461
rect 19521 27452 19533 27455
rect 18656 27424 19533 27452
rect 18656 27412 18662 27424
rect 19521 27421 19533 27424
rect 19567 27421 19579 27455
rect 19521 27415 19579 27421
rect 19610 27455 19668 27461
rect 19610 27421 19622 27455
rect 19656 27421 19668 27455
rect 19610 27415 19668 27421
rect 19705 27455 19763 27461
rect 19705 27421 19717 27455
rect 19751 27421 19763 27455
rect 19705 27415 19763 27421
rect 19889 27455 19947 27461
rect 19889 27421 19901 27455
rect 19935 27452 19947 27455
rect 20070 27452 20076 27464
rect 19935 27424 20076 27452
rect 19935 27421 19947 27424
rect 19889 27415 19947 27421
rect 15160 27356 17540 27384
rect 17580 27387 17638 27393
rect 15160 27344 15166 27356
rect 17580 27353 17592 27387
rect 17626 27384 17638 27387
rect 17678 27384 17684 27396
rect 17626 27356 17684 27384
rect 17626 27353 17638 27356
rect 17580 27347 17638 27353
rect 17678 27344 17684 27356
rect 17736 27344 17742 27396
rect 18782 27344 18788 27396
rect 18840 27384 18846 27396
rect 19720 27384 19748 27415
rect 20070 27412 20076 27424
rect 20128 27412 20134 27464
rect 20714 27452 20720 27464
rect 20675 27424 20720 27452
rect 20714 27412 20720 27424
rect 20772 27412 20778 27464
rect 21361 27455 21419 27461
rect 21361 27421 21373 27455
rect 21407 27452 21419 27455
rect 21910 27452 21916 27464
rect 21407 27424 21916 27452
rect 21407 27421 21419 27424
rect 21361 27415 21419 27421
rect 21910 27412 21916 27424
rect 21968 27412 21974 27464
rect 22281 27455 22339 27461
rect 22281 27421 22293 27455
rect 22327 27452 22339 27455
rect 22370 27452 22376 27464
rect 22327 27424 22376 27452
rect 22327 27421 22339 27424
rect 22281 27415 22339 27421
rect 22370 27412 22376 27424
rect 22428 27412 22434 27464
rect 22741 27455 22799 27461
rect 22741 27421 22753 27455
rect 22787 27452 22799 27455
rect 22922 27452 22928 27464
rect 22787 27424 22928 27452
rect 22787 27421 22799 27424
rect 22741 27415 22799 27421
rect 22922 27412 22928 27424
rect 22980 27412 22986 27464
rect 23382 27412 23388 27464
rect 23440 27452 23446 27464
rect 24118 27452 24124 27464
rect 23440 27424 24124 27452
rect 23440 27412 23446 27424
rect 24118 27412 24124 27424
rect 24176 27412 24182 27464
rect 24394 27452 24400 27464
rect 24355 27424 24400 27452
rect 24394 27412 24400 27424
rect 24452 27412 24458 27464
rect 25317 27455 25375 27461
rect 25317 27421 25329 27455
rect 25363 27452 25375 27455
rect 25498 27452 25504 27464
rect 25363 27424 25504 27452
rect 25363 27421 25375 27424
rect 25317 27415 25375 27421
rect 25498 27412 25504 27424
rect 25556 27412 25562 27464
rect 26694 27452 26700 27464
rect 26655 27424 26700 27452
rect 26694 27412 26700 27424
rect 26752 27412 26758 27464
rect 28718 27452 28724 27464
rect 28679 27424 28724 27452
rect 28718 27412 28724 27424
rect 28776 27412 28782 27464
rect 28902 27452 28908 27464
rect 28863 27424 28908 27452
rect 28902 27412 28908 27424
rect 28960 27412 28966 27464
rect 18840 27356 19748 27384
rect 18840 27344 18846 27356
rect 19978 27344 19984 27396
rect 20036 27384 20042 27396
rect 20533 27387 20591 27393
rect 20533 27384 20545 27387
rect 20036 27356 20545 27384
rect 20036 27344 20042 27356
rect 20533 27353 20545 27356
rect 20579 27353 20591 27387
rect 20533 27347 20591 27353
rect 20898 27344 20904 27396
rect 20956 27384 20962 27396
rect 21726 27384 21732 27396
rect 20956 27356 21732 27384
rect 20956 27344 20962 27356
rect 21726 27344 21732 27356
rect 21784 27384 21790 27396
rect 22005 27387 22063 27393
rect 22005 27384 22017 27387
rect 21784 27356 22017 27384
rect 21784 27344 21790 27356
rect 22005 27353 22017 27356
rect 22051 27353 22063 27387
rect 22005 27347 22063 27353
rect 25130 27344 25136 27396
rect 25188 27384 25194 27396
rect 26053 27387 26111 27393
rect 26053 27384 26065 27387
rect 25188 27356 26065 27384
rect 25188 27344 25194 27356
rect 26053 27353 26065 27356
rect 26099 27384 26111 27387
rect 26142 27384 26148 27396
rect 26099 27356 26148 27384
rect 26099 27353 26111 27356
rect 26053 27347 26111 27353
rect 26142 27344 26148 27356
rect 26200 27344 26206 27396
rect 26786 27344 26792 27396
rect 26844 27384 26850 27396
rect 26942 27387 27000 27393
rect 26942 27384 26954 27387
rect 26844 27356 26954 27384
rect 26844 27344 26850 27356
rect 26942 27353 26954 27356
rect 26988 27353 27000 27387
rect 26942 27347 27000 27353
rect 30184 27387 30242 27393
rect 30184 27353 30196 27387
rect 30230 27384 30242 27387
rect 30374 27384 30380 27396
rect 30230 27356 30380 27384
rect 30230 27353 30242 27356
rect 30184 27347 30242 27353
rect 30374 27344 30380 27356
rect 30432 27344 30438 27396
rect 8481 27319 8539 27325
rect 8481 27316 8493 27319
rect 7300 27288 8493 27316
rect 8481 27285 8493 27288
rect 8527 27285 8539 27319
rect 8938 27316 8944 27328
rect 8899 27288 8944 27316
rect 8481 27279 8539 27285
rect 8938 27276 8944 27288
rect 8996 27276 9002 27328
rect 9490 27276 9496 27328
rect 9548 27316 9554 27328
rect 16761 27319 16819 27325
rect 16761 27316 16773 27319
rect 9548 27288 16773 27316
rect 9548 27276 9554 27288
rect 16761 27285 16773 27288
rect 16807 27316 16819 27319
rect 18414 27316 18420 27328
rect 16807 27288 18420 27316
rect 16807 27285 16819 27288
rect 16761 27279 16819 27285
rect 18414 27276 18420 27288
rect 18472 27276 18478 27328
rect 18693 27319 18751 27325
rect 18693 27285 18705 27319
rect 18739 27316 18751 27319
rect 18877 27319 18935 27325
rect 18877 27316 18889 27319
rect 18739 27288 18889 27316
rect 18739 27285 18751 27288
rect 18693 27279 18751 27285
rect 18877 27285 18889 27288
rect 18923 27285 18935 27319
rect 18877 27279 18935 27285
rect 19058 27276 19064 27328
rect 19116 27316 19122 27328
rect 19245 27319 19303 27325
rect 19245 27316 19257 27319
rect 19116 27288 19257 27316
rect 19116 27276 19122 27288
rect 19245 27285 19257 27288
rect 19291 27285 19303 27319
rect 19245 27279 19303 27285
rect 22189 27319 22247 27325
rect 22189 27285 22201 27319
rect 22235 27316 22247 27319
rect 23566 27316 23572 27328
rect 22235 27288 23572 27316
rect 22235 27285 22247 27288
rect 22189 27279 22247 27285
rect 23566 27276 23572 27288
rect 23624 27276 23630 27328
rect 24673 27319 24731 27325
rect 24673 27285 24685 27319
rect 24719 27316 24731 27319
rect 24762 27316 24768 27328
rect 24719 27288 24768 27316
rect 24719 27285 24731 27288
rect 24673 27279 24731 27285
rect 24762 27276 24768 27288
rect 24820 27316 24826 27328
rect 28442 27316 28448 27328
rect 24820 27288 28448 27316
rect 24820 27276 24826 27288
rect 28442 27276 28448 27288
rect 28500 27276 28506 27328
rect 29362 27276 29368 27328
rect 29420 27316 29426 27328
rect 30098 27316 30104 27328
rect 29420 27288 30104 27316
rect 29420 27276 29426 27288
rect 30098 27276 30104 27288
rect 30156 27276 30162 27328
rect 1104 27226 32016 27248
rect 1104 27174 7288 27226
rect 7340 27174 17592 27226
rect 17644 27174 27896 27226
rect 27948 27174 32016 27226
rect 1104 27152 32016 27174
rect 1854 27072 1860 27124
rect 1912 27112 1918 27124
rect 2590 27112 2596 27124
rect 1912 27084 2596 27112
rect 1912 27072 1918 27084
rect 2590 27072 2596 27084
rect 2648 27072 2654 27124
rect 7190 27112 7196 27124
rect 7151 27084 7196 27112
rect 7190 27072 7196 27084
rect 7248 27072 7254 27124
rect 9490 27112 9496 27124
rect 8312 27084 9496 27112
rect 2682 27044 2688 27056
rect 1412 27016 2688 27044
rect 1412 26920 1440 27016
rect 2682 27004 2688 27016
rect 2740 27044 2746 27056
rect 8312 27044 8340 27084
rect 9490 27072 9496 27084
rect 9548 27072 9554 27124
rect 10318 27072 10324 27124
rect 10376 27112 10382 27124
rect 10965 27115 11023 27121
rect 10965 27112 10977 27115
rect 10376 27084 10977 27112
rect 10376 27072 10382 27084
rect 10965 27081 10977 27084
rect 11011 27081 11023 27115
rect 10965 27075 11023 27081
rect 11238 27072 11244 27124
rect 11296 27112 11302 27124
rect 11517 27115 11575 27121
rect 11517 27112 11529 27115
rect 11296 27084 11529 27112
rect 11296 27072 11302 27084
rect 11517 27081 11529 27084
rect 11563 27081 11575 27115
rect 11517 27075 11575 27081
rect 11606 27072 11612 27124
rect 11664 27112 11670 27124
rect 12526 27112 12532 27124
rect 11664 27084 12532 27112
rect 11664 27072 11670 27084
rect 12526 27072 12532 27084
rect 12584 27112 12590 27124
rect 12894 27112 12900 27124
rect 12584 27084 12900 27112
rect 12584 27072 12590 27084
rect 12894 27072 12900 27084
rect 12952 27112 12958 27124
rect 13170 27112 13176 27124
rect 12952 27084 13176 27112
rect 12952 27072 12958 27084
rect 13170 27072 13176 27084
rect 13228 27072 13234 27124
rect 13541 27115 13599 27121
rect 13541 27081 13553 27115
rect 13587 27112 13599 27115
rect 13630 27112 13636 27124
rect 13587 27084 13636 27112
rect 13587 27081 13599 27084
rect 13541 27075 13599 27081
rect 13630 27072 13636 27084
rect 13688 27072 13694 27124
rect 14093 27115 14151 27121
rect 14093 27081 14105 27115
rect 14139 27112 14151 27115
rect 17034 27112 17040 27124
rect 14139 27084 17040 27112
rect 14139 27081 14151 27084
rect 14093 27075 14151 27081
rect 17034 27072 17040 27084
rect 17092 27072 17098 27124
rect 17678 27112 17684 27124
rect 17639 27084 17684 27112
rect 17678 27072 17684 27084
rect 17736 27072 17742 27124
rect 18601 27115 18659 27121
rect 18601 27081 18613 27115
rect 18647 27112 18659 27115
rect 18647 27084 22232 27112
rect 18647 27081 18659 27084
rect 18601 27075 18659 27081
rect 2740 27016 3832 27044
rect 2740 27004 2746 27016
rect 1670 26985 1676 26988
rect 1664 26939 1676 26985
rect 1728 26976 1734 26988
rect 3804 26985 3832 27016
rect 6748 27016 8340 27044
rect 8380 27047 8438 27053
rect 4062 26985 4068 26988
rect 3789 26979 3847 26985
rect 1728 26948 1764 26976
rect 1670 26936 1676 26939
rect 1728 26936 1734 26948
rect 3789 26945 3801 26979
rect 3835 26945 3847 26979
rect 4056 26976 4068 26985
rect 4023 26948 4068 26976
rect 3789 26939 3847 26945
rect 4056 26939 4068 26948
rect 4062 26936 4068 26939
rect 4120 26936 4126 26988
rect 6748 26985 6776 27016
rect 8380 27013 8392 27047
rect 8426 27044 8438 27047
rect 8938 27044 8944 27056
rect 8426 27016 8944 27044
rect 8426 27013 8438 27016
rect 8380 27007 8438 27013
rect 8938 27004 8944 27016
rect 8996 27004 9002 27056
rect 10781 27047 10839 27053
rect 10781 27013 10793 27047
rect 10827 27044 10839 27047
rect 11149 27047 11207 27053
rect 11149 27044 11161 27047
rect 10827 27016 11161 27044
rect 10827 27013 10839 27016
rect 10781 27007 10839 27013
rect 11149 27013 11161 27016
rect 11195 27013 11207 27047
rect 11149 27007 11207 27013
rect 12621 27047 12679 27053
rect 12621 27013 12633 27047
rect 12667 27044 12679 27047
rect 12667 27016 13032 27044
rect 12667 27013 12679 27016
rect 12621 27007 12679 27013
rect 5813 26979 5871 26985
rect 5813 26945 5825 26979
rect 5859 26945 5871 26979
rect 5813 26939 5871 26945
rect 6549 26979 6607 26985
rect 6549 26945 6561 26979
rect 6595 26945 6607 26979
rect 6549 26939 6607 26945
rect 6733 26979 6791 26985
rect 6733 26945 6745 26979
rect 6779 26945 6791 26979
rect 7374 26976 7380 26988
rect 7335 26948 7380 26976
rect 6733 26939 6791 26945
rect 1394 26908 1400 26920
rect 1355 26880 1400 26908
rect 1394 26868 1400 26880
rect 1452 26868 1458 26920
rect 5828 26908 5856 26939
rect 4816 26880 5856 26908
rect 1762 26732 1768 26784
rect 1820 26772 1826 26784
rect 2682 26772 2688 26784
rect 1820 26744 2688 26772
rect 1820 26732 1826 26744
rect 2682 26732 2688 26744
rect 2740 26732 2746 26784
rect 2777 26775 2835 26781
rect 2777 26741 2789 26775
rect 2823 26772 2835 26775
rect 2866 26772 2872 26784
rect 2823 26744 2872 26772
rect 2823 26741 2835 26744
rect 2777 26735 2835 26741
rect 2866 26732 2872 26744
rect 2924 26732 2930 26784
rect 3142 26732 3148 26784
rect 3200 26772 3206 26784
rect 4816 26772 4844 26880
rect 5169 26843 5227 26849
rect 5169 26809 5181 26843
rect 5215 26840 5227 26843
rect 5718 26840 5724 26852
rect 5215 26812 5724 26840
rect 5215 26809 5227 26812
rect 5169 26803 5227 26809
rect 5718 26800 5724 26812
rect 5776 26800 5782 26852
rect 6564 26840 6592 26939
rect 7374 26936 7380 26948
rect 7432 26936 7438 26988
rect 7466 26936 7472 26988
rect 7524 26976 7530 26988
rect 7561 26979 7619 26985
rect 7561 26976 7573 26979
rect 7524 26948 7573 26976
rect 7524 26936 7530 26948
rect 7561 26945 7573 26948
rect 7607 26945 7619 26979
rect 7561 26939 7619 26945
rect 7653 26979 7711 26985
rect 7653 26945 7665 26979
rect 7699 26976 7711 26979
rect 7834 26976 7840 26988
rect 7699 26948 7840 26976
rect 7699 26945 7711 26948
rect 7653 26939 7711 26945
rect 7834 26936 7840 26948
rect 7892 26936 7898 26988
rect 8754 26936 8760 26988
rect 8812 26976 8818 26988
rect 11422 26976 11428 26988
rect 8812 26948 11428 26976
rect 8812 26936 8818 26948
rect 11422 26936 11428 26948
rect 11480 26936 11486 26988
rect 11698 26936 11704 26988
rect 11756 26976 11762 26988
rect 11793 26979 11851 26985
rect 11793 26976 11805 26979
rect 11756 26948 11805 26976
rect 11756 26936 11762 26948
rect 11793 26945 11805 26948
rect 11839 26945 11851 26979
rect 11885 26979 11943 26985
rect 11885 26972 11897 26979
rect 11931 26972 11943 26979
rect 11998 26979 12056 26985
rect 11793 26939 11851 26945
rect 11882 26920 11888 26972
rect 11940 26920 11946 26972
rect 11998 26945 12010 26979
rect 12044 26945 12056 26979
rect 11998 26939 12056 26945
rect 12161 26980 12219 26985
rect 12250 26980 12256 26988
rect 12161 26979 12256 26980
rect 12161 26945 12173 26979
rect 12207 26952 12256 26979
rect 12207 26945 12219 26952
rect 12161 26939 12219 26945
rect 8110 26908 8116 26920
rect 8071 26880 8116 26908
rect 8110 26868 8116 26880
rect 8168 26868 8174 26920
rect 10413 26911 10471 26917
rect 10413 26877 10425 26911
rect 10459 26908 10471 26911
rect 10870 26908 10876 26920
rect 10459 26880 10876 26908
rect 10459 26877 10471 26880
rect 10413 26871 10471 26877
rect 10870 26868 10876 26880
rect 10928 26908 10934 26920
rect 10928 26880 11836 26908
rect 10928 26868 10934 26880
rect 6564 26812 8156 26840
rect 5626 26772 5632 26784
rect 3200 26744 4844 26772
rect 5587 26744 5632 26772
rect 3200 26732 3206 26744
rect 5626 26732 5632 26744
rect 5684 26732 5690 26784
rect 6454 26732 6460 26784
rect 6512 26772 6518 26784
rect 6549 26775 6607 26781
rect 6549 26772 6561 26775
rect 6512 26744 6561 26772
rect 6512 26732 6518 26744
rect 6549 26741 6561 26744
rect 6595 26741 6607 26775
rect 6549 26735 6607 26741
rect 7374 26732 7380 26784
rect 7432 26772 7438 26784
rect 7650 26772 7656 26784
rect 7432 26744 7656 26772
rect 7432 26732 7438 26744
rect 7650 26732 7656 26744
rect 7708 26732 7714 26784
rect 8128 26772 8156 26812
rect 9214 26800 9220 26852
rect 9272 26840 9278 26852
rect 9493 26843 9551 26849
rect 9493 26840 9505 26843
rect 9272 26812 9505 26840
rect 9272 26800 9278 26812
rect 9493 26809 9505 26812
rect 9539 26809 9551 26843
rect 9493 26803 9551 26809
rect 9766 26800 9772 26852
rect 9824 26840 9830 26852
rect 10594 26840 10600 26852
rect 9824 26812 10600 26840
rect 9824 26800 9830 26812
rect 10594 26800 10600 26812
rect 10652 26800 10658 26852
rect 11238 26840 11244 26852
rect 10704 26812 11244 26840
rect 10704 26772 10732 26812
rect 11238 26800 11244 26812
rect 11296 26800 11302 26852
rect 11808 26840 11836 26880
rect 11882 26840 11888 26852
rect 11808 26812 11888 26840
rect 11882 26800 11888 26812
rect 11940 26800 11946 26852
rect 12013 26840 12041 26939
rect 12250 26936 12256 26952
rect 12308 26936 12314 26988
rect 12529 26979 12587 26985
rect 12529 26945 12541 26979
rect 12575 26976 12587 26979
rect 12710 26976 12716 26988
rect 12575 26948 12716 26976
rect 12575 26945 12587 26948
rect 12529 26939 12587 26945
rect 12710 26936 12716 26948
rect 12768 26936 12774 26988
rect 12805 26979 12863 26985
rect 12805 26945 12817 26979
rect 12851 26976 12863 26979
rect 12894 26976 12900 26988
rect 12851 26948 12900 26976
rect 12851 26945 12863 26948
rect 12805 26939 12863 26945
rect 12894 26936 12900 26948
rect 12952 26936 12958 26988
rect 13004 26908 13032 27016
rect 13446 27004 13452 27056
rect 13504 27044 13510 27056
rect 15286 27044 15292 27056
rect 13504 27016 15292 27044
rect 13504 27004 13510 27016
rect 15286 27004 15292 27016
rect 15344 27044 15350 27056
rect 19978 27044 19984 27056
rect 15344 27016 19984 27044
rect 15344 27004 15350 27016
rect 19978 27004 19984 27016
rect 20036 27004 20042 27056
rect 20809 27047 20867 27053
rect 20809 27013 20821 27047
rect 20855 27044 20867 27047
rect 22066 27047 22124 27053
rect 22066 27044 22078 27047
rect 20855 27016 22078 27044
rect 20855 27013 20867 27016
rect 20809 27007 20867 27013
rect 22066 27013 22078 27016
rect 22112 27013 22124 27047
rect 22204 27044 22232 27084
rect 22922 27072 22928 27124
rect 22980 27112 22986 27124
rect 23201 27115 23259 27121
rect 23201 27112 23213 27115
rect 22980 27084 23213 27112
rect 22980 27072 22986 27084
rect 23201 27081 23213 27084
rect 23247 27081 23259 27115
rect 23201 27075 23259 27081
rect 23474 27072 23480 27124
rect 23532 27112 23538 27124
rect 25038 27112 25044 27124
rect 23532 27084 25044 27112
rect 23532 27072 23538 27084
rect 25038 27072 25044 27084
rect 25096 27112 25102 27124
rect 25501 27115 25559 27121
rect 25501 27112 25513 27115
rect 25096 27084 25513 27112
rect 25096 27072 25102 27084
rect 25501 27081 25513 27084
rect 25547 27081 25559 27115
rect 25501 27075 25559 27081
rect 25961 27115 26019 27121
rect 25961 27081 25973 27115
rect 26007 27112 26019 27115
rect 26786 27112 26792 27124
rect 26007 27084 26792 27112
rect 26007 27081 26019 27084
rect 25961 27075 26019 27081
rect 26786 27072 26792 27084
rect 26844 27072 26850 27124
rect 27338 27072 27344 27124
rect 27396 27112 27402 27124
rect 30374 27112 30380 27124
rect 27396 27084 29408 27112
rect 30335 27084 30380 27112
rect 27396 27072 27402 27084
rect 23382 27044 23388 27056
rect 22204 27016 23388 27044
rect 22066 27007 22124 27013
rect 23382 27004 23388 27016
rect 23440 27004 23446 27056
rect 23569 27047 23627 27053
rect 23569 27013 23581 27047
rect 23615 27044 23627 27047
rect 25866 27044 25872 27056
rect 23615 27016 25872 27044
rect 23615 27013 23627 27016
rect 23569 27007 23627 27013
rect 25866 27004 25872 27016
rect 25924 27004 25930 27056
rect 26326 27004 26332 27056
rect 26384 27044 26390 27056
rect 26384 27016 27476 27044
rect 26384 27004 26390 27016
rect 13722 26976 13728 26988
rect 13683 26948 13728 26976
rect 13722 26936 13728 26948
rect 13780 26936 13786 26988
rect 13998 26976 14004 26988
rect 13959 26948 14004 26976
rect 13998 26936 14004 26948
rect 14056 26936 14062 26988
rect 14366 26936 14372 26988
rect 14424 26976 14430 26988
rect 14461 26979 14519 26985
rect 14461 26976 14473 26979
rect 14424 26948 14473 26976
rect 14424 26936 14430 26948
rect 14461 26945 14473 26948
rect 14507 26945 14519 26979
rect 14461 26939 14519 26945
rect 14645 26979 14703 26985
rect 14645 26945 14657 26979
rect 14691 26945 14703 26979
rect 14645 26939 14703 26945
rect 14737 26979 14795 26985
rect 14737 26945 14749 26979
rect 14783 26976 14795 26979
rect 14783 26948 15332 26976
rect 14783 26945 14795 26948
rect 14737 26939 14795 26945
rect 14093 26911 14151 26917
rect 14093 26908 14105 26911
rect 13004 26880 14105 26908
rect 14093 26877 14105 26880
rect 14139 26877 14151 26911
rect 14093 26871 14151 26877
rect 14182 26868 14188 26920
rect 14240 26908 14246 26920
rect 14660 26908 14688 26939
rect 14240 26880 14688 26908
rect 14240 26868 14246 26880
rect 12989 26843 13047 26849
rect 12989 26840 13001 26843
rect 12013 26812 13001 26840
rect 12989 26809 13001 26812
rect 13035 26809 13047 26843
rect 15304 26840 15332 26948
rect 15378 26936 15384 26988
rect 15436 26976 15442 26988
rect 15749 26979 15807 26985
rect 15749 26976 15761 26979
rect 15436 26948 15761 26976
rect 15436 26936 15442 26948
rect 15749 26945 15761 26948
rect 15795 26945 15807 26979
rect 15749 26939 15807 26945
rect 15933 26979 15991 26985
rect 15933 26945 15945 26979
rect 15979 26976 15991 26979
rect 16206 26976 16212 26988
rect 15979 26948 16212 26976
rect 15979 26945 15991 26948
rect 15933 26939 15991 26945
rect 16206 26936 16212 26948
rect 16264 26936 16270 26988
rect 16942 26976 16948 26988
rect 16903 26948 16948 26976
rect 16942 26936 16948 26948
rect 17000 26936 17006 26988
rect 17862 26976 17868 26988
rect 17823 26948 17868 26976
rect 17862 26936 17868 26948
rect 17920 26936 17926 26988
rect 18141 26979 18199 26985
rect 18141 26945 18153 26979
rect 18187 26976 18199 26979
rect 18598 26976 18604 26988
rect 18187 26948 18604 26976
rect 18187 26945 18199 26948
rect 18141 26939 18199 26945
rect 18598 26936 18604 26948
rect 18656 26976 18662 26988
rect 18877 26979 18935 26985
rect 18877 26976 18889 26979
rect 18656 26948 18889 26976
rect 18656 26936 18662 26948
rect 18877 26945 18889 26948
rect 18923 26945 18935 26979
rect 19058 26976 19064 26988
rect 19019 26948 19064 26976
rect 18877 26939 18935 26945
rect 19058 26936 19064 26948
rect 19116 26936 19122 26988
rect 20070 26976 20076 26988
rect 20031 26948 20076 26976
rect 20070 26936 20076 26948
rect 20128 26936 20134 26988
rect 20349 26979 20407 26985
rect 20349 26945 20361 26979
rect 20395 26976 20407 26979
rect 20714 26976 20720 26988
rect 20395 26948 20720 26976
rect 20395 26945 20407 26948
rect 20349 26939 20407 26945
rect 20714 26936 20720 26948
rect 20772 26936 20778 26988
rect 20990 26976 20996 26988
rect 20951 26948 20996 26976
rect 20990 26936 20996 26948
rect 21048 26936 21054 26988
rect 21818 26976 21824 26988
rect 21779 26948 21824 26976
rect 21818 26936 21824 26948
rect 21876 26936 21882 26988
rect 22370 26936 22376 26988
rect 22428 26976 22434 26988
rect 22830 26976 22836 26988
rect 22428 26948 22836 26976
rect 22428 26936 22434 26948
rect 22830 26936 22836 26948
rect 22888 26936 22894 26988
rect 23474 26936 23480 26988
rect 23532 26976 23538 26988
rect 27448 26985 27476 27016
rect 24377 26979 24435 26985
rect 24377 26976 24389 26979
rect 23532 26948 24389 26976
rect 23532 26936 23538 26948
rect 24377 26945 24389 26948
rect 24423 26945 24435 26979
rect 24377 26939 24435 26945
rect 26145 26979 26203 26985
rect 26145 26945 26157 26979
rect 26191 26976 26203 26979
rect 26973 26979 27031 26985
rect 26973 26976 26985 26979
rect 26191 26948 26985 26976
rect 26191 26945 26203 26948
rect 26145 26939 26203 26945
rect 26973 26945 26985 26948
rect 27019 26945 27031 26979
rect 26973 26939 27031 26945
rect 27157 26979 27215 26985
rect 27157 26945 27169 26979
rect 27203 26945 27215 26979
rect 27157 26939 27215 26945
rect 27433 26979 27491 26985
rect 27433 26945 27445 26979
rect 27479 26945 27491 26979
rect 27433 26939 27491 26945
rect 16482 26868 16488 26920
rect 16540 26908 16546 26920
rect 18785 26911 18843 26917
rect 18785 26908 18797 26911
rect 16540 26880 18797 26908
rect 16540 26868 16546 26880
rect 18785 26877 18797 26880
rect 18831 26877 18843 26911
rect 18785 26871 18843 26877
rect 18969 26911 19027 26917
rect 18969 26877 18981 26911
rect 19015 26908 19027 26911
rect 19334 26908 19340 26920
rect 19015 26880 19340 26908
rect 19015 26877 19027 26880
rect 18969 26871 19027 26877
rect 16574 26840 16580 26852
rect 15304 26812 16580 26840
rect 12989 26803 13047 26809
rect 16574 26800 16580 26812
rect 16632 26800 16638 26852
rect 18800 26840 18828 26871
rect 19334 26868 19340 26880
rect 19392 26868 19398 26920
rect 19702 26868 19708 26920
rect 19760 26908 19766 26920
rect 20806 26908 20812 26920
rect 19760 26880 20812 26908
rect 19760 26868 19766 26880
rect 20806 26868 20812 26880
rect 20864 26868 20870 26920
rect 21174 26868 21180 26920
rect 21232 26908 21238 26920
rect 21269 26911 21327 26917
rect 21269 26908 21281 26911
rect 21232 26880 21281 26908
rect 21232 26868 21238 26880
rect 21269 26877 21281 26880
rect 21315 26877 21327 26911
rect 24118 26908 24124 26920
rect 24079 26880 24124 26908
rect 21269 26871 21327 26877
rect 24118 26868 24124 26880
rect 24176 26868 24182 26920
rect 26418 26908 26424 26920
rect 26379 26880 26424 26908
rect 26418 26868 26424 26880
rect 26476 26868 26482 26920
rect 19058 26840 19064 26852
rect 18800 26812 19064 26840
rect 19058 26800 19064 26812
rect 19116 26800 19122 26852
rect 20257 26843 20315 26849
rect 20257 26840 20269 26843
rect 19306 26812 20269 26840
rect 8128 26744 10732 26772
rect 10781 26775 10839 26781
rect 10781 26741 10793 26775
rect 10827 26772 10839 26775
rect 11054 26772 11060 26784
rect 10827 26744 11060 26772
rect 10827 26741 10839 26744
rect 10781 26735 10839 26741
rect 11054 26732 11060 26744
rect 11112 26732 11118 26784
rect 11149 26775 11207 26781
rect 11149 26741 11161 26775
rect 11195 26772 11207 26775
rect 12529 26775 12587 26781
rect 12529 26772 12541 26775
rect 11195 26744 12541 26772
rect 11195 26741 11207 26744
rect 11149 26735 11207 26741
rect 12529 26741 12541 26744
rect 12575 26741 12587 26775
rect 13906 26772 13912 26784
rect 13867 26744 13912 26772
rect 12529 26735 12587 26741
rect 13906 26732 13912 26744
rect 13964 26732 13970 26784
rect 13998 26732 14004 26784
rect 14056 26772 14062 26784
rect 14461 26775 14519 26781
rect 14461 26772 14473 26775
rect 14056 26744 14473 26772
rect 14056 26732 14062 26744
rect 14461 26741 14473 26744
rect 14507 26741 14519 26775
rect 14461 26735 14519 26741
rect 16117 26775 16175 26781
rect 16117 26741 16129 26775
rect 16163 26772 16175 26775
rect 16666 26772 16672 26784
rect 16163 26744 16672 26772
rect 16163 26741 16175 26744
rect 16117 26735 16175 26741
rect 16666 26732 16672 26744
rect 16724 26732 16730 26784
rect 17126 26772 17132 26784
rect 17087 26744 17132 26772
rect 17126 26732 17132 26744
rect 17184 26732 17190 26784
rect 18049 26775 18107 26781
rect 18049 26741 18061 26775
rect 18095 26772 18107 26775
rect 18414 26772 18420 26784
rect 18095 26744 18420 26772
rect 18095 26741 18107 26744
rect 18049 26735 18107 26741
rect 18414 26732 18420 26744
rect 18472 26772 18478 26784
rect 19306 26772 19334 26812
rect 20257 26809 20269 26812
rect 20303 26809 20315 26843
rect 26329 26843 26387 26849
rect 26329 26840 26341 26843
rect 20257 26803 20315 26809
rect 25148 26812 26341 26840
rect 19886 26772 19892 26784
rect 18472 26744 19334 26772
rect 19847 26744 19892 26772
rect 18472 26732 18478 26744
rect 19886 26732 19892 26744
rect 19944 26732 19950 26784
rect 21082 26732 21088 26784
rect 21140 26772 21146 26784
rect 21177 26775 21235 26781
rect 21177 26772 21189 26775
rect 21140 26744 21189 26772
rect 21140 26732 21146 26744
rect 21177 26741 21189 26744
rect 21223 26741 21235 26775
rect 21177 26735 21235 26741
rect 22186 26732 22192 26784
rect 22244 26772 22250 26784
rect 23569 26775 23627 26781
rect 23569 26772 23581 26775
rect 22244 26744 23581 26772
rect 22244 26732 22250 26744
rect 23569 26741 23581 26744
rect 23615 26741 23627 26775
rect 23569 26735 23627 26741
rect 23750 26732 23756 26784
rect 23808 26772 23814 26784
rect 24762 26772 24768 26784
rect 23808 26744 24768 26772
rect 23808 26732 23814 26744
rect 24762 26732 24768 26744
rect 24820 26772 24826 26784
rect 25148 26772 25176 26812
rect 26329 26809 26341 26812
rect 26375 26809 26387 26843
rect 26329 26803 26387 26809
rect 24820 26744 25176 26772
rect 24820 26732 24826 26744
rect 25222 26732 25228 26784
rect 25280 26772 25286 26784
rect 27172 26772 27200 26939
rect 27522 26936 27528 26988
rect 27580 26976 27586 26988
rect 27617 26979 27675 26985
rect 27617 26976 27629 26979
rect 27580 26948 27629 26976
rect 27580 26936 27586 26948
rect 27617 26945 27629 26948
rect 27663 26945 27675 26979
rect 27617 26939 27675 26945
rect 27982 26936 27988 26988
rect 28040 26976 28046 26988
rect 28261 26979 28319 26985
rect 28261 26976 28273 26979
rect 28040 26948 28273 26976
rect 28040 26936 28046 26948
rect 28261 26945 28273 26948
rect 28307 26945 28319 26979
rect 29178 26976 29184 26988
rect 29139 26948 29184 26976
rect 28261 26939 28319 26945
rect 29178 26936 29184 26948
rect 29236 26936 29242 26988
rect 29380 26985 29408 27084
rect 30374 27072 30380 27084
rect 30432 27072 30438 27124
rect 29365 26979 29423 26985
rect 29365 26945 29377 26979
rect 29411 26976 29423 26979
rect 29914 26976 29920 26988
rect 29411 26948 29920 26976
rect 29411 26945 29423 26948
rect 29365 26939 29423 26945
rect 29914 26936 29920 26948
rect 29972 26936 29978 26988
rect 30558 26976 30564 26988
rect 30519 26948 30564 26976
rect 30558 26936 30564 26948
rect 30616 26936 30622 26988
rect 28534 26908 28540 26920
rect 28495 26880 28540 26908
rect 28534 26868 28540 26880
rect 28592 26868 28598 26920
rect 29454 26908 29460 26920
rect 29415 26880 29460 26908
rect 29454 26868 29460 26880
rect 29512 26868 29518 26920
rect 30837 26911 30895 26917
rect 30837 26877 30849 26911
rect 30883 26908 30895 26911
rect 31018 26908 31024 26920
rect 30883 26880 31024 26908
rect 30883 26877 30895 26880
rect 30837 26871 30895 26877
rect 31018 26868 31024 26880
rect 31076 26868 31082 26920
rect 28902 26800 28908 26852
rect 28960 26840 28966 26852
rect 30745 26843 30803 26849
rect 30745 26840 30757 26843
rect 28960 26812 30757 26840
rect 28960 26800 28966 26812
rect 30745 26809 30757 26812
rect 30791 26809 30803 26843
rect 30745 26803 30803 26809
rect 28074 26772 28080 26784
rect 25280 26744 27200 26772
rect 28035 26744 28080 26772
rect 25280 26732 25286 26744
rect 28074 26732 28080 26744
rect 28132 26732 28138 26784
rect 28442 26772 28448 26784
rect 28403 26744 28448 26772
rect 28442 26732 28448 26744
rect 28500 26732 28506 26784
rect 28626 26732 28632 26784
rect 28684 26772 28690 26784
rect 28997 26775 29055 26781
rect 28997 26772 29009 26775
rect 28684 26744 29009 26772
rect 28684 26732 28690 26744
rect 28997 26741 29009 26744
rect 29043 26741 29055 26775
rect 28997 26735 29055 26741
rect 1104 26682 32016 26704
rect 1104 26630 2136 26682
rect 2188 26630 12440 26682
rect 12492 26630 22744 26682
rect 22796 26630 32016 26682
rect 1104 26608 32016 26630
rect 4154 26528 4160 26580
rect 4212 26568 4218 26580
rect 4433 26571 4491 26577
rect 4433 26568 4445 26571
rect 4212 26540 4445 26568
rect 4212 26528 4218 26540
rect 4433 26537 4445 26540
rect 4479 26537 4491 26571
rect 5534 26568 5540 26580
rect 5495 26540 5540 26568
rect 4433 26531 4491 26537
rect 5534 26528 5540 26540
rect 5592 26528 5598 26580
rect 5718 26568 5724 26580
rect 5644 26540 5724 26568
rect 3053 26503 3111 26509
rect 3053 26469 3065 26503
rect 3099 26500 3111 26503
rect 3326 26500 3332 26512
rect 3099 26472 3332 26500
rect 3099 26469 3111 26472
rect 3053 26463 3111 26469
rect 3326 26460 3332 26472
rect 3384 26460 3390 26512
rect 2498 26392 2504 26444
rect 2556 26432 2562 26444
rect 4522 26432 4528 26444
rect 2556 26404 4528 26432
rect 2556 26392 2562 26404
rect 4522 26392 4528 26404
rect 4580 26392 4586 26444
rect 1854 26324 1860 26376
rect 1912 26364 1918 26376
rect 2133 26367 2191 26373
rect 2133 26364 2145 26367
rect 1912 26336 2145 26364
rect 1912 26324 1918 26336
rect 2133 26333 2145 26336
rect 2179 26333 2191 26367
rect 2133 26327 2191 26333
rect 2409 26367 2467 26373
rect 2409 26333 2421 26367
rect 2455 26333 2467 26367
rect 2409 26327 2467 26333
rect 2593 26367 2651 26373
rect 2593 26333 2605 26367
rect 2639 26364 2651 26367
rect 2866 26364 2872 26376
rect 2639 26336 2872 26364
rect 2639 26333 2651 26336
rect 2593 26327 2651 26333
rect 0 26296 800 26310
rect 1486 26296 1492 26308
rect 0 26268 1492 26296
rect 0 26254 800 26268
rect 1486 26256 1492 26268
rect 1544 26256 1550 26308
rect 2424 26296 2452 26327
rect 2866 26324 2872 26336
rect 2924 26324 2930 26376
rect 3234 26364 3240 26376
rect 3195 26336 3240 26364
rect 3234 26324 3240 26336
rect 3292 26324 3298 26376
rect 3973 26367 4031 26373
rect 3973 26333 3985 26367
rect 4019 26364 4031 26367
rect 4062 26364 4068 26376
rect 4019 26336 4068 26364
rect 4019 26333 4031 26336
rect 3973 26327 4031 26333
rect 4062 26324 4068 26336
rect 4120 26324 4126 26376
rect 4617 26367 4675 26373
rect 4617 26333 4629 26367
rect 4663 26364 4675 26367
rect 4706 26364 4712 26376
rect 4663 26336 4712 26364
rect 4663 26333 4675 26336
rect 4617 26327 4675 26333
rect 4706 26324 4712 26336
rect 4764 26324 4770 26376
rect 4893 26367 4951 26373
rect 4893 26333 4905 26367
rect 4939 26364 4951 26367
rect 4982 26364 4988 26376
rect 4939 26336 4988 26364
rect 4939 26333 4951 26336
rect 4893 26327 4951 26333
rect 4982 26324 4988 26336
rect 5040 26324 5046 26376
rect 5077 26367 5135 26373
rect 5077 26333 5089 26367
rect 5123 26364 5135 26367
rect 5644 26364 5672 26540
rect 5718 26528 5724 26540
rect 5776 26568 5782 26580
rect 7098 26568 7104 26580
rect 5776 26540 7104 26568
rect 5776 26528 5782 26540
rect 7098 26528 7104 26540
rect 7156 26528 7162 26580
rect 7834 26528 7840 26580
rect 7892 26568 7898 26580
rect 8113 26571 8171 26577
rect 8113 26568 8125 26571
rect 7892 26540 8125 26568
rect 7892 26528 7898 26540
rect 8113 26537 8125 26540
rect 8159 26568 8171 26571
rect 8386 26568 8392 26580
rect 8159 26540 8392 26568
rect 8159 26537 8171 26540
rect 8113 26531 8171 26537
rect 8386 26528 8392 26540
rect 8444 26528 8450 26580
rect 9125 26571 9183 26577
rect 9125 26537 9137 26571
rect 9171 26568 9183 26571
rect 11606 26568 11612 26580
rect 9171 26540 11612 26568
rect 9171 26537 9183 26540
rect 9125 26531 9183 26537
rect 11606 26528 11612 26540
rect 11664 26528 11670 26580
rect 11885 26571 11943 26577
rect 11885 26537 11897 26571
rect 11931 26568 11943 26571
rect 12805 26571 12863 26577
rect 12805 26568 12817 26571
rect 11931 26540 12817 26568
rect 11931 26537 11943 26540
rect 11885 26531 11943 26537
rect 12805 26537 12817 26540
rect 12851 26568 12863 26571
rect 13081 26571 13139 26577
rect 13081 26568 13093 26571
rect 12851 26540 13093 26568
rect 12851 26537 12863 26540
rect 12805 26531 12863 26537
rect 13081 26537 13093 26540
rect 13127 26537 13139 26571
rect 13081 26531 13139 26537
rect 13449 26571 13507 26577
rect 13449 26537 13461 26571
rect 13495 26568 13507 26571
rect 16942 26568 16948 26580
rect 13495 26540 16948 26568
rect 13495 26537 13507 26540
rect 13449 26531 13507 26537
rect 16942 26528 16948 26540
rect 17000 26528 17006 26580
rect 17126 26528 17132 26580
rect 17184 26568 17190 26580
rect 17184 26540 20760 26568
rect 17184 26528 17190 26540
rect 11790 26460 11796 26512
rect 11848 26500 11854 26512
rect 13998 26500 14004 26512
rect 11848 26472 14004 26500
rect 11848 26460 11854 26472
rect 13998 26460 14004 26472
rect 14056 26460 14062 26512
rect 14090 26460 14096 26512
rect 14148 26500 14154 26512
rect 15470 26500 15476 26512
rect 14148 26472 15476 26500
rect 14148 26460 14154 26472
rect 15470 26460 15476 26472
rect 15528 26460 15534 26512
rect 18230 26460 18236 26512
rect 18288 26500 18294 26512
rect 18509 26503 18567 26509
rect 18509 26500 18521 26503
rect 18288 26472 18521 26500
rect 18288 26460 18294 26472
rect 18509 26469 18521 26472
rect 18555 26469 18567 26503
rect 20732 26500 20760 26540
rect 20990 26528 20996 26580
rect 21048 26568 21054 26580
rect 21637 26571 21695 26577
rect 21637 26568 21649 26571
rect 21048 26540 21649 26568
rect 21048 26528 21054 26540
rect 21637 26537 21649 26540
rect 21683 26537 21695 26571
rect 21637 26531 21695 26537
rect 22833 26571 22891 26577
rect 22833 26537 22845 26571
rect 22879 26568 22891 26571
rect 23014 26568 23020 26580
rect 22879 26540 23020 26568
rect 22879 26537 22891 26540
rect 22833 26531 22891 26537
rect 23014 26528 23020 26540
rect 23072 26528 23078 26580
rect 23385 26571 23443 26577
rect 23385 26537 23397 26571
rect 23431 26568 23443 26571
rect 23474 26568 23480 26580
rect 23431 26540 23480 26568
rect 23431 26537 23443 26540
rect 23385 26531 23443 26537
rect 23474 26528 23480 26540
rect 23532 26528 23538 26580
rect 26694 26568 26700 26580
rect 24044 26540 26700 26568
rect 22557 26503 22615 26509
rect 22557 26500 22569 26503
rect 20732 26472 22569 26500
rect 18509 26463 18567 26469
rect 22557 26469 22569 26472
rect 22603 26469 22615 26503
rect 23750 26500 23756 26512
rect 23711 26472 23756 26500
rect 22557 26463 22615 26469
rect 23750 26460 23756 26472
rect 23808 26460 23814 26512
rect 11977 26435 12035 26441
rect 11977 26401 11989 26435
rect 12023 26432 12035 26435
rect 12526 26432 12532 26444
rect 12023 26404 12532 26432
rect 12023 26401 12035 26404
rect 11977 26395 12035 26401
rect 12526 26392 12532 26404
rect 12584 26392 12590 26444
rect 12710 26392 12716 26444
rect 12768 26392 12774 26444
rect 12894 26432 12900 26444
rect 12855 26404 12900 26432
rect 12894 26392 12900 26404
rect 12952 26392 12958 26444
rect 13538 26392 13544 26444
rect 13596 26432 13602 26444
rect 18141 26435 18199 26441
rect 13596 26404 15608 26432
rect 13596 26392 13602 26404
rect 5123 26336 5672 26364
rect 5721 26367 5779 26373
rect 5123 26333 5135 26336
rect 5077 26327 5135 26333
rect 5721 26333 5733 26367
rect 5767 26364 5779 26367
rect 5810 26364 5816 26376
rect 5767 26336 5816 26364
rect 5767 26333 5779 26336
rect 5721 26327 5779 26333
rect 5810 26324 5816 26336
rect 5868 26324 5874 26376
rect 5997 26367 6055 26373
rect 5997 26333 6009 26367
rect 6043 26333 6055 26367
rect 5997 26327 6055 26333
rect 6181 26367 6239 26373
rect 6181 26333 6193 26367
rect 6227 26333 6239 26367
rect 6181 26327 6239 26333
rect 4798 26296 4804 26308
rect 2424 26268 4804 26296
rect 4798 26256 4804 26268
rect 4856 26256 4862 26308
rect 5000 26296 5028 26324
rect 6012 26296 6040 26327
rect 5000 26268 6040 26296
rect 6196 26296 6224 26327
rect 6362 26324 6368 26376
rect 6420 26364 6426 26376
rect 6733 26367 6791 26373
rect 6733 26364 6745 26367
rect 6420 26336 6745 26364
rect 6420 26324 6426 26336
rect 6733 26333 6745 26336
rect 6779 26364 6791 26367
rect 6822 26364 6828 26376
rect 6779 26336 6828 26364
rect 6779 26333 6791 26336
rect 6733 26327 6791 26333
rect 6822 26324 6828 26336
rect 6880 26324 6886 26376
rect 7006 26373 7012 26376
rect 7000 26364 7012 26373
rect 6967 26336 7012 26364
rect 7000 26327 7012 26336
rect 7006 26324 7012 26327
rect 7064 26324 7070 26376
rect 8110 26324 8116 26376
rect 8168 26364 8174 26376
rect 9677 26367 9735 26373
rect 9677 26364 9689 26367
rect 8168 26336 9689 26364
rect 8168 26324 8174 26336
rect 9677 26333 9689 26336
rect 9723 26364 9735 26367
rect 11514 26364 11520 26376
rect 9723 26336 11520 26364
rect 9723 26333 9735 26336
rect 9677 26327 9735 26333
rect 11514 26324 11520 26336
rect 11572 26324 11578 26376
rect 11701 26367 11759 26373
rect 11701 26333 11713 26367
rect 11747 26364 11759 26367
rect 11790 26364 11796 26376
rect 11747 26336 11796 26364
rect 11747 26333 11759 26336
rect 11701 26327 11759 26333
rect 11790 26324 11796 26336
rect 11848 26324 11854 26376
rect 11882 26324 11888 26376
rect 11940 26364 11946 26376
rect 12250 26364 12256 26376
rect 11940 26336 12256 26364
rect 11940 26324 11946 26336
rect 12250 26324 12256 26336
rect 12308 26324 12314 26376
rect 12621 26367 12679 26373
rect 12621 26333 12633 26367
rect 12667 26333 12679 26367
rect 12728 26364 12756 26392
rect 13357 26367 13415 26373
rect 13357 26364 13369 26367
rect 12728 26336 13369 26364
rect 12621 26327 12679 26333
rect 13357 26333 13369 26336
rect 13403 26364 13415 26367
rect 13630 26364 13636 26376
rect 13403 26336 13636 26364
rect 13403 26333 13415 26336
rect 13357 26327 13415 26333
rect 6914 26296 6920 26308
rect 6196 26268 6920 26296
rect 6914 26256 6920 26268
rect 6972 26256 6978 26308
rect 9033 26299 9091 26305
rect 9033 26265 9045 26299
rect 9079 26296 9091 26299
rect 9766 26296 9772 26308
rect 9079 26268 9772 26296
rect 9079 26265 9091 26268
rect 9033 26259 9091 26265
rect 9766 26256 9772 26268
rect 9824 26256 9830 26308
rect 9944 26299 10002 26305
rect 9944 26265 9956 26299
rect 9990 26296 10002 26299
rect 12437 26299 12495 26305
rect 12437 26296 12449 26299
rect 9990 26268 12449 26296
rect 9990 26265 10002 26268
rect 9944 26259 10002 26265
rect 12437 26265 12449 26268
rect 12483 26265 12495 26299
rect 12636 26296 12664 26327
rect 13630 26324 13636 26336
rect 13688 26324 13694 26376
rect 13814 26324 13820 26376
rect 13872 26364 13878 26376
rect 14645 26367 14703 26373
rect 14645 26364 14657 26367
rect 13872 26336 14657 26364
rect 13872 26324 13878 26336
rect 14645 26333 14657 26336
rect 14691 26333 14703 26367
rect 15286 26364 15292 26376
rect 15247 26336 15292 26364
rect 14645 26327 14703 26333
rect 15286 26324 15292 26336
rect 15344 26324 15350 26376
rect 15580 26373 15608 26404
rect 18141 26401 18153 26435
rect 18187 26432 18199 26435
rect 19702 26432 19708 26444
rect 18187 26404 19708 26432
rect 18187 26401 18199 26404
rect 18141 26395 18199 26401
rect 19702 26392 19708 26404
rect 19760 26392 19766 26444
rect 21634 26392 21640 26444
rect 21692 26432 21698 26444
rect 24044 26432 24072 26540
rect 26694 26528 26700 26540
rect 26752 26528 26758 26580
rect 29914 26568 29920 26580
rect 29875 26540 29920 26568
rect 29914 26528 29920 26540
rect 29972 26568 29978 26580
rect 30837 26571 30895 26577
rect 30837 26568 30849 26571
rect 29972 26540 30849 26568
rect 29972 26528 29978 26540
rect 30837 26537 30849 26540
rect 30883 26568 30895 26571
rect 30926 26568 30932 26580
rect 30883 26540 30932 26568
rect 30883 26537 30895 26540
rect 30837 26531 30895 26537
rect 30926 26528 30932 26540
rect 30984 26528 30990 26580
rect 29730 26460 29736 26512
rect 29788 26500 29794 26512
rect 29788 26472 30972 26500
rect 29788 26460 29794 26472
rect 21692 26404 21864 26432
rect 21692 26392 21698 26404
rect 15565 26367 15623 26373
rect 15565 26333 15577 26367
rect 15611 26364 15623 26367
rect 15654 26364 15660 26376
rect 15611 26336 15660 26364
rect 15611 26333 15623 26336
rect 15565 26327 15623 26333
rect 15654 26324 15660 26336
rect 15712 26324 15718 26376
rect 15749 26367 15807 26373
rect 15749 26333 15761 26367
rect 15795 26364 15807 26367
rect 15838 26364 15844 26376
rect 15795 26336 15844 26364
rect 15795 26333 15807 26336
rect 15749 26327 15807 26333
rect 15838 26324 15844 26336
rect 15896 26324 15902 26376
rect 16666 26324 16672 26376
rect 16724 26364 16730 26376
rect 16761 26367 16819 26373
rect 16761 26364 16773 26367
rect 16724 26336 16773 26364
rect 16724 26324 16730 26336
rect 16761 26333 16773 26336
rect 16807 26333 16819 26367
rect 16761 26327 16819 26333
rect 17126 26324 17132 26376
rect 17184 26364 17190 26376
rect 17402 26364 17408 26376
rect 17184 26336 17408 26364
rect 17184 26324 17190 26336
rect 17402 26324 17408 26336
rect 17460 26324 17466 26376
rect 17494 26324 17500 26376
rect 17552 26364 17558 26376
rect 17681 26367 17739 26373
rect 17681 26364 17693 26367
rect 17552 26336 17693 26364
rect 17552 26324 17558 26336
rect 17681 26333 17693 26336
rect 17727 26333 17739 26367
rect 17681 26327 17739 26333
rect 17954 26324 17960 26376
rect 18012 26364 18018 26376
rect 18509 26367 18567 26373
rect 18509 26364 18521 26367
rect 18012 26336 18521 26364
rect 18012 26324 18018 26336
rect 18509 26333 18521 26336
rect 18555 26333 18567 26367
rect 18690 26364 18696 26376
rect 18651 26336 18696 26364
rect 18509 26327 18567 26333
rect 18690 26324 18696 26336
rect 18748 26324 18754 26376
rect 19797 26367 19855 26373
rect 19797 26333 19809 26367
rect 19843 26364 19855 26367
rect 20806 26364 20812 26376
rect 19843 26336 20812 26364
rect 19843 26333 19855 26336
rect 19797 26327 19855 26333
rect 20806 26324 20812 26336
rect 20864 26364 20870 26376
rect 21726 26364 21732 26376
rect 20864 26336 21732 26364
rect 20864 26324 20870 26336
rect 21726 26324 21732 26336
rect 21784 26324 21790 26376
rect 21836 26373 21864 26404
rect 23492 26404 24072 26432
rect 21821 26367 21879 26373
rect 21821 26333 21833 26367
rect 21867 26333 21879 26367
rect 21821 26327 21879 26333
rect 22097 26367 22155 26373
rect 22097 26333 22109 26367
rect 22143 26333 22155 26367
rect 22097 26327 22155 26333
rect 22281 26367 22339 26373
rect 22281 26333 22293 26367
rect 22327 26364 22339 26367
rect 22646 26364 22652 26376
rect 22327 26336 22652 26364
rect 22327 26333 22339 26336
rect 22281 26327 22339 26333
rect 12710 26296 12716 26308
rect 12636 26268 12716 26296
rect 12437 26259 12495 26265
rect 12710 26256 12716 26268
rect 12768 26256 12774 26308
rect 13081 26299 13139 26305
rect 13081 26265 13093 26299
rect 13127 26296 13139 26299
rect 13832 26296 13860 26324
rect 14458 26296 14464 26308
rect 13127 26268 13860 26296
rect 14419 26268 14464 26296
rect 13127 26265 13139 26268
rect 13081 26259 13139 26265
rect 14458 26256 14464 26268
rect 14516 26296 14522 26308
rect 14918 26296 14924 26308
rect 14516 26268 14924 26296
rect 14516 26256 14522 26268
rect 14918 26256 14924 26268
rect 14976 26256 14982 26308
rect 15105 26299 15163 26305
rect 15105 26265 15117 26299
rect 15151 26296 15163 26299
rect 15378 26296 15384 26308
rect 15151 26268 15384 26296
rect 15151 26265 15163 26268
rect 15105 26259 15163 26265
rect 15378 26256 15384 26268
rect 15436 26256 15442 26308
rect 16574 26256 16580 26308
rect 16632 26296 16638 26308
rect 18049 26299 18107 26305
rect 18049 26296 18061 26299
rect 16632 26268 18061 26296
rect 16632 26256 16638 26268
rect 18049 26265 18061 26268
rect 18095 26296 18107 26299
rect 18230 26296 18236 26308
rect 18095 26268 18236 26296
rect 18095 26265 18107 26268
rect 18049 26259 18107 26265
rect 18230 26256 18236 26268
rect 18288 26296 18294 26308
rect 18288 26268 19334 26296
rect 18288 26256 18294 26268
rect 1762 26188 1768 26240
rect 1820 26228 1826 26240
rect 1949 26231 2007 26237
rect 1949 26228 1961 26231
rect 1820 26200 1961 26228
rect 1820 26188 1826 26200
rect 1949 26197 1961 26200
rect 1995 26197 2007 26231
rect 3786 26228 3792 26240
rect 3747 26200 3792 26228
rect 1949 26191 2007 26197
rect 3786 26188 3792 26200
rect 3844 26188 3850 26240
rect 5074 26188 5080 26240
rect 5132 26228 5138 26240
rect 9674 26228 9680 26240
rect 5132 26200 9680 26228
rect 5132 26188 5138 26200
rect 9674 26188 9680 26200
rect 9732 26188 9738 26240
rect 10870 26188 10876 26240
rect 10928 26228 10934 26240
rect 11057 26231 11115 26237
rect 11057 26228 11069 26231
rect 10928 26200 11069 26228
rect 10928 26188 10934 26200
rect 11057 26197 11069 26200
rect 11103 26197 11115 26231
rect 11057 26191 11115 26197
rect 11517 26231 11575 26237
rect 11517 26197 11529 26231
rect 11563 26228 11575 26231
rect 11606 26228 11612 26240
rect 11563 26200 11612 26228
rect 11563 26197 11575 26200
rect 11517 26191 11575 26197
rect 11606 26188 11612 26200
rect 11664 26188 11670 26240
rect 11698 26188 11704 26240
rect 11756 26228 11762 26240
rect 14182 26228 14188 26240
rect 11756 26200 14188 26228
rect 11756 26188 11762 26200
rect 14182 26188 14188 26200
rect 14240 26188 14246 26240
rect 16666 26188 16672 26240
rect 16724 26228 16730 26240
rect 16853 26231 16911 26237
rect 16853 26228 16865 26231
rect 16724 26200 16865 26228
rect 16724 26188 16730 26200
rect 16853 26197 16865 26200
rect 16899 26228 16911 26231
rect 18141 26231 18199 26237
rect 18141 26228 18153 26231
rect 16899 26200 18153 26228
rect 16899 26197 16911 26200
rect 16853 26191 16911 26197
rect 18141 26197 18153 26200
rect 18187 26197 18199 26231
rect 19306 26228 19334 26268
rect 19886 26256 19892 26308
rect 19944 26296 19950 26308
rect 20042 26299 20100 26305
rect 20042 26296 20054 26299
rect 19944 26268 20054 26296
rect 19944 26256 19950 26268
rect 20042 26265 20054 26268
rect 20088 26265 20100 26299
rect 22112 26296 22140 26327
rect 22646 26324 22652 26336
rect 22704 26324 22710 26376
rect 22741 26367 22799 26373
rect 22741 26333 22753 26367
rect 22787 26333 22799 26367
rect 22922 26364 22928 26376
rect 22883 26336 22928 26364
rect 22741 26327 22799 26333
rect 22462 26296 22468 26308
rect 20042 26259 20100 26265
rect 20180 26268 21404 26296
rect 22112 26268 22468 26296
rect 20180 26228 20208 26268
rect 21174 26228 21180 26240
rect 19306 26200 20208 26228
rect 21135 26200 21180 26228
rect 18141 26191 18199 26197
rect 21174 26188 21180 26200
rect 21232 26188 21238 26240
rect 21376 26228 21404 26268
rect 22462 26256 22468 26268
rect 22520 26256 22526 26308
rect 22557 26299 22615 26305
rect 22557 26265 22569 26299
rect 22603 26296 22615 26299
rect 22756 26296 22784 26327
rect 22922 26324 22928 26336
rect 22980 26324 22986 26376
rect 23492 26296 23520 26404
rect 24118 26392 24124 26444
rect 24176 26432 24182 26444
rect 24176 26404 25544 26432
rect 24176 26392 24182 26404
rect 23569 26367 23627 26373
rect 23569 26333 23581 26367
rect 23615 26333 23627 26367
rect 23569 26327 23627 26333
rect 23845 26367 23903 26373
rect 23845 26333 23857 26367
rect 23891 26364 23903 26367
rect 24486 26364 24492 26376
rect 23891 26336 24492 26364
rect 23891 26333 23903 26336
rect 23845 26327 23903 26333
rect 22603 26268 23520 26296
rect 23584 26296 23612 26327
rect 24486 26324 24492 26336
rect 24544 26324 24550 26376
rect 24581 26367 24639 26373
rect 24581 26333 24593 26367
rect 24627 26333 24639 26367
rect 24581 26327 24639 26333
rect 24857 26367 24915 26373
rect 24857 26333 24869 26367
rect 24903 26333 24915 26367
rect 25038 26364 25044 26376
rect 24999 26336 25044 26364
rect 24857 26327 24915 26333
rect 24397 26299 24455 26305
rect 24397 26296 24409 26299
rect 23584 26268 24409 26296
rect 22603 26265 22615 26268
rect 22557 26259 22615 26265
rect 24397 26265 24409 26268
rect 24443 26265 24455 26299
rect 24397 26259 24455 26265
rect 22830 26228 22836 26240
rect 21376 26200 22836 26228
rect 22830 26188 22836 26200
rect 22888 26188 22894 26240
rect 24596 26228 24624 26327
rect 24872 26296 24900 26327
rect 25038 26324 25044 26336
rect 25096 26324 25102 26376
rect 25516 26373 25544 26404
rect 28994 26392 29000 26444
rect 29052 26432 29058 26444
rect 30009 26435 30067 26441
rect 30009 26432 30021 26435
rect 29052 26404 30021 26432
rect 29052 26392 29058 26404
rect 30009 26401 30021 26404
rect 30055 26401 30067 26435
rect 30009 26395 30067 26401
rect 30098 26392 30104 26444
rect 30156 26432 30162 26444
rect 30944 26441 30972 26472
rect 30929 26435 30987 26441
rect 30156 26404 30788 26432
rect 30156 26392 30162 26404
rect 25501 26367 25559 26373
rect 25501 26333 25513 26367
rect 25547 26364 25559 26367
rect 26786 26364 26792 26376
rect 25547 26336 26792 26364
rect 25547 26333 25559 26336
rect 25501 26327 25559 26333
rect 26786 26324 26792 26336
rect 26844 26364 26850 26376
rect 27617 26367 27675 26373
rect 27617 26364 27629 26367
rect 26844 26336 27629 26364
rect 26844 26324 26850 26336
rect 27617 26333 27629 26336
rect 27663 26364 27675 26367
rect 27706 26364 27712 26376
rect 27663 26336 27712 26364
rect 27663 26333 27675 26336
rect 27617 26327 27675 26333
rect 27706 26324 27712 26336
rect 27764 26324 27770 26376
rect 29086 26324 29092 26376
rect 29144 26364 29150 26376
rect 29733 26367 29791 26373
rect 29733 26364 29745 26367
rect 29144 26336 29745 26364
rect 29144 26324 29150 26336
rect 29733 26333 29745 26336
rect 29779 26333 29791 26367
rect 29733 26327 29791 26333
rect 30558 26324 30564 26376
rect 30616 26364 30622 26376
rect 30653 26367 30711 26373
rect 30653 26364 30665 26367
rect 30616 26336 30665 26364
rect 30616 26324 30622 26336
rect 30653 26333 30665 26336
rect 30699 26333 30711 26367
rect 30653 26327 30711 26333
rect 25768 26299 25826 26305
rect 24872 26268 25728 26296
rect 25222 26228 25228 26240
rect 24596 26200 25228 26228
rect 25222 26188 25228 26200
rect 25280 26188 25286 26240
rect 25700 26228 25728 26268
rect 25768 26265 25780 26299
rect 25814 26296 25826 26299
rect 26970 26296 26976 26308
rect 25814 26268 26976 26296
rect 25814 26265 25826 26268
rect 25768 26259 25826 26265
rect 26970 26256 26976 26268
rect 27028 26256 27034 26308
rect 27884 26299 27942 26305
rect 27884 26265 27896 26299
rect 27930 26296 27942 26299
rect 29549 26299 29607 26305
rect 29549 26296 29561 26299
rect 27930 26268 29561 26296
rect 27930 26265 27942 26268
rect 27884 26259 27942 26265
rect 29549 26265 29561 26268
rect 29595 26265 29607 26299
rect 29549 26259 29607 26265
rect 30098 26256 30104 26308
rect 30156 26296 30162 26308
rect 30469 26299 30527 26305
rect 30469 26296 30481 26299
rect 30156 26268 30481 26296
rect 30156 26256 30162 26268
rect 30469 26265 30481 26268
rect 30515 26265 30527 26299
rect 30760 26296 30788 26404
rect 30929 26401 30941 26435
rect 30975 26401 30987 26435
rect 30929 26395 30987 26401
rect 32320 26296 33120 26310
rect 30760 26268 33120 26296
rect 30469 26259 30527 26265
rect 32320 26254 33120 26268
rect 26326 26228 26332 26240
rect 25700 26200 26332 26228
rect 26326 26188 26332 26200
rect 26384 26188 26390 26240
rect 26510 26188 26516 26240
rect 26568 26228 26574 26240
rect 26881 26231 26939 26237
rect 26881 26228 26893 26231
rect 26568 26200 26893 26228
rect 26568 26188 26574 26200
rect 26881 26197 26893 26200
rect 26927 26197 26939 26231
rect 26881 26191 26939 26197
rect 28997 26231 29055 26237
rect 28997 26197 29009 26231
rect 29043 26228 29055 26231
rect 29730 26228 29736 26240
rect 29043 26200 29736 26228
rect 29043 26197 29055 26200
rect 28997 26191 29055 26197
rect 29730 26188 29736 26200
rect 29788 26188 29794 26240
rect 1104 26138 32016 26160
rect 1104 26086 7288 26138
rect 7340 26086 17592 26138
rect 17644 26086 27896 26138
rect 27948 26086 32016 26138
rect 1104 26064 32016 26086
rect 1581 26027 1639 26033
rect 1581 25993 1593 26027
rect 1627 26024 1639 26027
rect 1670 26024 1676 26036
rect 1627 25996 1676 26024
rect 1627 25993 1639 25996
rect 1581 25987 1639 25993
rect 1670 25984 1676 25996
rect 1728 25984 1734 26036
rect 2222 25984 2228 26036
rect 2280 26024 2286 26036
rect 6733 26027 6791 26033
rect 6733 26024 6745 26027
rect 2280 25996 6745 26024
rect 2280 25984 2286 25996
rect 6733 25993 6745 25996
rect 6779 25993 6791 26027
rect 9398 26024 9404 26036
rect 6733 25987 6791 25993
rect 6840 25996 9404 26024
rect 1302 25916 1308 25968
rect 1360 25956 1366 25968
rect 2240 25956 2268 25984
rect 2774 25965 2780 25968
rect 2768 25956 2780 25965
rect 1360 25928 2268 25956
rect 2735 25928 2780 25956
rect 1360 25916 1366 25928
rect 2768 25919 2780 25928
rect 2774 25916 2780 25919
rect 2832 25916 2838 25968
rect 4338 25956 4344 25968
rect 4299 25928 4344 25956
rect 4338 25916 4344 25928
rect 4396 25916 4402 25968
rect 5721 25959 5779 25965
rect 5721 25925 5733 25959
rect 5767 25956 5779 25959
rect 6840 25956 6868 25996
rect 9398 25984 9404 25996
rect 9456 25984 9462 26036
rect 12802 26024 12808 26036
rect 9683 25996 12808 26024
rect 5767 25928 6868 25956
rect 5767 25925 5779 25928
rect 5721 25919 5779 25925
rect 6914 25916 6920 25968
rect 6972 25956 6978 25968
rect 9493 25959 9551 25965
rect 9493 25956 9505 25959
rect 6972 25928 9505 25956
rect 6972 25916 6978 25928
rect 9493 25925 9505 25928
rect 9539 25956 9551 25959
rect 9582 25956 9588 25968
rect 9539 25928 9588 25956
rect 9539 25925 9551 25928
rect 9493 25919 9551 25925
rect 9582 25916 9588 25928
rect 9640 25916 9646 25968
rect 1762 25888 1768 25900
rect 1723 25860 1768 25888
rect 1762 25848 1768 25860
rect 1820 25848 1826 25900
rect 1854 25848 1860 25900
rect 1912 25888 1918 25900
rect 4525 25891 4583 25897
rect 4525 25888 4537 25891
rect 1912 25860 4537 25888
rect 1912 25848 1918 25860
rect 4525 25857 4537 25860
rect 4571 25857 4583 25891
rect 4798 25888 4804 25900
rect 4759 25860 4804 25888
rect 4525 25851 4583 25857
rect 4798 25848 4804 25860
rect 4856 25848 4862 25900
rect 4985 25891 5043 25897
rect 4985 25857 4997 25891
rect 5031 25857 5043 25891
rect 4985 25851 5043 25857
rect 5629 25891 5687 25897
rect 5629 25857 5641 25891
rect 5675 25857 5687 25891
rect 5629 25851 5687 25857
rect 5813 25891 5871 25897
rect 5813 25857 5825 25891
rect 5859 25888 5871 25891
rect 7742 25888 7748 25900
rect 5859 25860 7604 25888
rect 7655 25860 7748 25888
rect 5859 25857 5871 25860
rect 5813 25851 5871 25857
rect 1670 25780 1676 25832
rect 1728 25820 1734 25832
rect 2041 25823 2099 25829
rect 2041 25820 2053 25823
rect 1728 25792 2053 25820
rect 1728 25780 1734 25792
rect 2041 25789 2053 25792
rect 2087 25789 2099 25823
rect 2041 25783 2099 25789
rect 2501 25823 2559 25829
rect 2501 25789 2513 25823
rect 2547 25789 2559 25823
rect 5000 25820 5028 25851
rect 2501 25783 2559 25789
rect 4448 25792 5028 25820
rect 5644 25820 5672 25851
rect 6270 25820 6276 25832
rect 5644 25792 6276 25820
rect 1394 25712 1400 25764
rect 1452 25752 1458 25764
rect 2516 25752 2544 25783
rect 1452 25724 2544 25752
rect 1452 25712 1458 25724
rect 4448 25696 4476 25792
rect 6270 25780 6276 25792
rect 6328 25780 6334 25832
rect 6825 25823 6883 25829
rect 6825 25789 6837 25823
rect 6871 25789 6883 25823
rect 6825 25783 6883 25789
rect 7009 25823 7067 25829
rect 7009 25789 7021 25823
rect 7055 25820 7067 25823
rect 7576 25820 7604 25860
rect 7742 25848 7748 25860
rect 7800 25888 7806 25900
rect 9306 25888 9312 25900
rect 7800 25860 9312 25888
rect 7800 25848 7806 25860
rect 9306 25848 9312 25860
rect 9364 25848 9370 25900
rect 9683 25820 9711 25996
rect 12802 25984 12808 25996
rect 12860 25984 12866 26036
rect 12894 25984 12900 26036
rect 12952 26024 12958 26036
rect 12952 25996 13045 26024
rect 12952 25984 12958 25996
rect 14826 25984 14832 26036
rect 14884 26024 14890 26036
rect 16666 26024 16672 26036
rect 14884 25996 16672 26024
rect 14884 25984 14890 25996
rect 16666 25984 16672 25996
rect 16724 25984 16730 26036
rect 18506 26024 18512 26036
rect 16776 25996 18512 26024
rect 11054 25916 11060 25968
rect 11112 25956 11118 25968
rect 11112 25928 12296 25956
rect 11112 25916 11118 25928
rect 10505 25891 10563 25897
rect 10505 25857 10517 25891
rect 10551 25888 10563 25891
rect 10594 25888 10600 25900
rect 10551 25860 10600 25888
rect 10551 25857 10563 25860
rect 10505 25851 10563 25857
rect 10594 25848 10600 25860
rect 10652 25848 10658 25900
rect 10781 25891 10839 25897
rect 10781 25857 10793 25891
rect 10827 25857 10839 25891
rect 10781 25851 10839 25857
rect 7055 25792 7144 25820
rect 7576 25792 9711 25820
rect 7055 25789 7067 25792
rect 7009 25783 7067 25789
rect 5994 25712 6000 25764
rect 6052 25752 6058 25764
rect 6840 25752 6868 25783
rect 6052 25724 6868 25752
rect 6052 25712 6058 25724
rect 1578 25644 1584 25696
rect 1636 25684 1642 25696
rect 1949 25687 2007 25693
rect 1949 25684 1961 25687
rect 1636 25656 1961 25684
rect 1636 25644 1642 25656
rect 1949 25653 1961 25656
rect 1995 25653 2007 25687
rect 1949 25647 2007 25653
rect 3881 25687 3939 25693
rect 3881 25653 3893 25687
rect 3927 25684 3939 25687
rect 4430 25684 4436 25696
rect 3927 25656 4436 25684
rect 3927 25653 3939 25656
rect 3881 25647 3939 25653
rect 4430 25644 4436 25656
rect 4488 25644 4494 25696
rect 6365 25687 6423 25693
rect 6365 25653 6377 25687
rect 6411 25684 6423 25687
rect 6546 25684 6552 25696
rect 6411 25656 6552 25684
rect 6411 25653 6423 25656
rect 6365 25647 6423 25653
rect 6546 25644 6552 25656
rect 6604 25644 6610 25696
rect 6730 25644 6736 25696
rect 6788 25684 6794 25696
rect 7116 25684 7144 25792
rect 10318 25780 10324 25832
rect 10376 25820 10382 25832
rect 10796 25820 10824 25851
rect 10870 25848 10876 25900
rect 10928 25888 10934 25900
rect 10965 25891 11023 25897
rect 10965 25888 10977 25891
rect 10928 25860 10977 25888
rect 10928 25848 10934 25860
rect 10965 25857 10977 25860
rect 11011 25857 11023 25891
rect 11514 25888 11520 25900
rect 11475 25860 11520 25888
rect 10965 25851 11023 25857
rect 11514 25848 11520 25860
rect 11572 25848 11578 25900
rect 11606 25848 11612 25900
rect 11664 25888 11670 25900
rect 11773 25891 11831 25897
rect 11773 25888 11785 25891
rect 11664 25860 11785 25888
rect 11664 25848 11670 25860
rect 11773 25857 11785 25860
rect 11819 25857 11831 25891
rect 12268 25888 12296 25928
rect 12342 25916 12348 25968
rect 12400 25956 12406 25968
rect 12710 25956 12716 25968
rect 12400 25928 12716 25956
rect 12400 25916 12406 25928
rect 12710 25916 12716 25928
rect 12768 25916 12774 25968
rect 12912 25888 12940 25984
rect 13630 25916 13636 25968
rect 13688 25956 13694 25968
rect 16114 25956 16120 25968
rect 13688 25928 16120 25956
rect 13688 25916 13694 25928
rect 16114 25916 16120 25928
rect 16172 25916 16178 25968
rect 13538 25888 13544 25900
rect 12268 25860 12940 25888
rect 13499 25860 13544 25888
rect 11773 25851 11831 25857
rect 13538 25848 13544 25860
rect 13596 25848 13602 25900
rect 14550 25888 14556 25900
rect 14511 25860 14556 25888
rect 14550 25848 14556 25860
rect 14608 25848 14614 25900
rect 14820 25891 14878 25897
rect 14820 25857 14832 25891
rect 14866 25888 14878 25891
rect 15194 25888 15200 25900
rect 14866 25860 15200 25888
rect 14866 25857 14878 25860
rect 14820 25851 14878 25857
rect 15194 25848 15200 25860
rect 15252 25848 15258 25900
rect 16298 25848 16304 25900
rect 16356 25888 16362 25900
rect 16776 25897 16804 25996
rect 18506 25984 18512 25996
rect 18564 25984 18570 26036
rect 20070 25984 20076 26036
rect 20128 26024 20134 26036
rect 20165 26027 20223 26033
rect 20165 26024 20177 26027
rect 20128 25996 20177 26024
rect 20128 25984 20134 25996
rect 20165 25993 20177 25996
rect 20211 25993 20223 26027
rect 20165 25987 20223 25993
rect 21818 25984 21824 26036
rect 21876 26024 21882 26036
rect 23477 26027 23535 26033
rect 23477 26024 23489 26027
rect 21876 25996 23489 26024
rect 21876 25984 21882 25996
rect 23477 25993 23489 25996
rect 23523 25993 23535 26027
rect 23477 25987 23535 25993
rect 16942 25916 16948 25968
rect 17000 25956 17006 25968
rect 19337 25959 19395 25965
rect 19337 25956 19349 25959
rect 17000 25928 19349 25956
rect 17000 25916 17006 25928
rect 19337 25925 19349 25928
rect 19383 25925 19395 25959
rect 19337 25919 19395 25925
rect 19426 25916 19432 25968
rect 19484 25956 19490 25968
rect 22189 25959 22247 25965
rect 22189 25956 22201 25959
rect 19484 25928 22201 25956
rect 19484 25916 19490 25928
rect 22189 25925 22201 25928
rect 22235 25925 22247 25959
rect 22189 25919 22247 25925
rect 16761 25891 16819 25897
rect 16761 25888 16773 25891
rect 16356 25860 16773 25888
rect 16356 25848 16362 25860
rect 16761 25857 16773 25860
rect 16807 25857 16819 25891
rect 16761 25851 16819 25857
rect 17672 25891 17730 25897
rect 17672 25857 17684 25891
rect 17718 25888 17730 25891
rect 18046 25888 18052 25900
rect 17718 25860 18052 25888
rect 17718 25857 17730 25860
rect 17672 25851 17730 25857
rect 18046 25848 18052 25860
rect 18104 25848 18110 25900
rect 19518 25888 19524 25900
rect 19479 25860 19524 25888
rect 19518 25848 19524 25860
rect 19576 25848 19582 25900
rect 20349 25891 20407 25897
rect 20349 25857 20361 25891
rect 20395 25857 20407 25891
rect 20622 25888 20628 25900
rect 20583 25860 20628 25888
rect 20349 25851 20407 25857
rect 10376 25792 10824 25820
rect 10376 25780 10382 25792
rect 12802 25780 12808 25832
rect 12860 25820 12866 25832
rect 13630 25820 13636 25832
rect 12860 25792 13636 25820
rect 12860 25780 12866 25792
rect 13630 25780 13636 25792
rect 13688 25820 13694 25832
rect 13817 25823 13875 25829
rect 13817 25820 13829 25823
rect 13688 25792 13829 25820
rect 13688 25780 13694 25792
rect 13817 25789 13829 25792
rect 13863 25789 13875 25823
rect 13817 25783 13875 25789
rect 16850 25780 16856 25832
rect 16908 25820 16914 25832
rect 17310 25820 17316 25832
rect 16908 25792 17316 25820
rect 16908 25780 16914 25792
rect 17310 25780 17316 25792
rect 17368 25820 17374 25832
rect 17405 25823 17463 25829
rect 17405 25820 17417 25823
rect 17368 25792 17417 25820
rect 17368 25780 17374 25792
rect 17405 25789 17417 25792
rect 17451 25789 17463 25823
rect 17405 25783 17463 25789
rect 19426 25780 19432 25832
rect 19484 25820 19490 25832
rect 20364 25820 20392 25851
rect 20622 25848 20628 25860
rect 20680 25848 20686 25900
rect 20809 25891 20867 25897
rect 20809 25857 20821 25891
rect 20855 25888 20867 25891
rect 21174 25888 21180 25900
rect 20855 25860 21180 25888
rect 20855 25857 20867 25860
rect 20809 25851 20867 25857
rect 21174 25848 21180 25860
rect 21232 25848 21238 25900
rect 23492 25888 23520 25987
rect 24486 25984 24492 26036
rect 24544 26024 24550 26036
rect 25777 26027 25835 26033
rect 25777 26024 25789 26027
rect 24544 25996 25789 26024
rect 24544 25984 24550 25996
rect 25777 25993 25789 25996
rect 25823 25993 25835 26027
rect 25777 25987 25835 25993
rect 23750 25916 23756 25968
rect 23808 25956 23814 25968
rect 24642 25959 24700 25965
rect 24642 25956 24654 25959
rect 23808 25928 24654 25956
rect 23808 25916 23814 25928
rect 24642 25925 24654 25928
rect 24688 25925 24700 25959
rect 24642 25919 24700 25925
rect 24397 25891 24455 25897
rect 24397 25888 24409 25891
rect 23492 25860 24409 25888
rect 24397 25857 24409 25860
rect 24443 25857 24455 25891
rect 25792 25888 25820 25987
rect 29908 25959 29966 25965
rect 27724 25928 29684 25956
rect 27724 25900 27752 25928
rect 26973 25891 27031 25897
rect 26973 25888 26985 25891
rect 25792 25860 26985 25888
rect 24397 25851 24455 25857
rect 26973 25857 26985 25860
rect 27019 25857 27031 25891
rect 26973 25851 27031 25857
rect 27617 25891 27675 25897
rect 27617 25857 27629 25891
rect 27663 25888 27675 25891
rect 27706 25888 27712 25900
rect 27663 25860 27712 25888
rect 27663 25857 27675 25860
rect 27617 25851 27675 25857
rect 27706 25848 27712 25860
rect 27764 25848 27770 25900
rect 27884 25891 27942 25897
rect 27884 25857 27896 25891
rect 27930 25888 27942 25891
rect 28626 25888 28632 25900
rect 27930 25860 28632 25888
rect 27930 25857 27942 25860
rect 27884 25851 27942 25857
rect 28626 25848 28632 25860
rect 28684 25848 28690 25900
rect 29656 25897 29684 25928
rect 29908 25925 29920 25959
rect 29954 25956 29966 25959
rect 30098 25956 30104 25968
rect 29954 25928 30104 25956
rect 29954 25925 29966 25928
rect 29908 25919 29966 25925
rect 30098 25916 30104 25928
rect 30156 25916 30162 25968
rect 29641 25891 29699 25897
rect 29641 25857 29653 25891
rect 29687 25857 29699 25891
rect 29641 25851 29699 25857
rect 21634 25820 21640 25832
rect 19484 25792 21640 25820
rect 19484 25780 19490 25792
rect 21634 25780 21640 25792
rect 21692 25780 21698 25832
rect 22186 25780 22192 25832
rect 22244 25820 22250 25832
rect 23198 25820 23204 25832
rect 22244 25792 23204 25820
rect 22244 25780 22250 25792
rect 23198 25780 23204 25792
rect 23256 25780 23262 25832
rect 8202 25712 8208 25764
rect 8260 25752 8266 25764
rect 11054 25752 11060 25764
rect 8260 25724 11060 25752
rect 8260 25712 8266 25724
rect 11054 25712 11060 25724
rect 11112 25712 11118 25764
rect 9214 25684 9220 25696
rect 6788 25656 9220 25684
rect 6788 25644 6794 25656
rect 9214 25644 9220 25656
rect 9272 25644 9278 25696
rect 9306 25644 9312 25696
rect 9364 25684 9370 25696
rect 10226 25684 10232 25696
rect 9364 25656 10232 25684
rect 9364 25644 9370 25656
rect 10226 25644 10232 25656
rect 10284 25644 10290 25696
rect 10321 25687 10379 25693
rect 10321 25653 10333 25687
rect 10367 25684 10379 25687
rect 12618 25684 12624 25696
rect 10367 25656 12624 25684
rect 10367 25653 10379 25656
rect 10321 25647 10379 25653
rect 12618 25644 12624 25656
rect 12676 25644 12682 25696
rect 13078 25644 13084 25696
rect 13136 25684 13142 25696
rect 13357 25687 13415 25693
rect 13357 25684 13369 25687
rect 13136 25656 13369 25684
rect 13136 25644 13142 25656
rect 13357 25653 13369 25656
rect 13403 25653 13415 25687
rect 13357 25647 13415 25653
rect 13725 25687 13783 25693
rect 13725 25653 13737 25687
rect 13771 25684 13783 25687
rect 13906 25684 13912 25696
rect 13771 25656 13912 25684
rect 13771 25653 13783 25656
rect 13725 25647 13783 25653
rect 13906 25644 13912 25656
rect 13964 25684 13970 25696
rect 14918 25684 14924 25696
rect 13964 25656 14924 25684
rect 13964 25644 13970 25656
rect 14918 25644 14924 25656
rect 14976 25644 14982 25696
rect 15838 25644 15844 25696
rect 15896 25684 15902 25696
rect 15933 25687 15991 25693
rect 15933 25684 15945 25687
rect 15896 25656 15945 25684
rect 15896 25644 15902 25656
rect 15933 25653 15945 25656
rect 15979 25653 15991 25687
rect 15933 25647 15991 25653
rect 16853 25687 16911 25693
rect 16853 25653 16865 25687
rect 16899 25684 16911 25687
rect 17402 25684 17408 25696
rect 16899 25656 17408 25684
rect 16899 25653 16911 25656
rect 16853 25647 16911 25653
rect 17402 25644 17408 25656
rect 17460 25644 17466 25696
rect 18690 25644 18696 25696
rect 18748 25684 18754 25696
rect 18785 25687 18843 25693
rect 18785 25684 18797 25687
rect 18748 25656 18797 25684
rect 18748 25644 18754 25656
rect 18785 25653 18797 25656
rect 18831 25653 18843 25687
rect 18785 25647 18843 25653
rect 23566 25644 23572 25696
rect 23624 25684 23630 25696
rect 27065 25687 27123 25693
rect 27065 25684 27077 25687
rect 23624 25656 27077 25684
rect 23624 25644 23630 25656
rect 27065 25653 27077 25656
rect 27111 25653 27123 25687
rect 28994 25684 29000 25696
rect 28955 25656 29000 25684
rect 27065 25647 27123 25653
rect 28994 25644 29000 25656
rect 29052 25644 29058 25696
rect 31021 25687 31079 25693
rect 31021 25653 31033 25687
rect 31067 25684 31079 25687
rect 31110 25684 31116 25696
rect 31067 25656 31116 25684
rect 31067 25653 31079 25656
rect 31021 25647 31079 25653
rect 31110 25644 31116 25656
rect 31168 25644 31174 25696
rect 1104 25594 32016 25616
rect 1104 25542 2136 25594
rect 2188 25542 12440 25594
rect 12492 25542 22744 25594
rect 22796 25542 32016 25594
rect 1104 25520 32016 25542
rect 3881 25483 3939 25489
rect 3881 25449 3893 25483
rect 3927 25480 3939 25483
rect 3970 25480 3976 25492
rect 3927 25452 3976 25480
rect 3927 25449 3939 25452
rect 3881 25443 3939 25449
rect 3970 25440 3976 25452
rect 4028 25440 4034 25492
rect 6089 25483 6147 25489
rect 6089 25449 6101 25483
rect 6135 25480 6147 25483
rect 6546 25480 6552 25492
rect 6135 25452 6552 25480
rect 6135 25449 6147 25452
rect 6089 25443 6147 25449
rect 6546 25440 6552 25452
rect 6604 25440 6610 25492
rect 8297 25483 8355 25489
rect 8297 25449 8309 25483
rect 8343 25480 8355 25483
rect 11698 25480 11704 25492
rect 8343 25452 11704 25480
rect 8343 25449 8355 25452
rect 8297 25443 8355 25449
rect 11698 25440 11704 25452
rect 11756 25440 11762 25492
rect 11974 25440 11980 25492
rect 12032 25480 12038 25492
rect 12989 25483 13047 25489
rect 12989 25480 13001 25483
rect 12032 25452 13001 25480
rect 12032 25440 12038 25452
rect 12989 25449 13001 25452
rect 13035 25449 13047 25483
rect 12989 25443 13047 25449
rect 13630 25440 13636 25492
rect 13688 25480 13694 25492
rect 13909 25483 13967 25489
rect 13909 25480 13921 25483
rect 13688 25452 13921 25480
rect 13688 25440 13694 25452
rect 13909 25449 13921 25452
rect 13955 25449 13967 25483
rect 15194 25480 15200 25492
rect 15155 25452 15200 25480
rect 13909 25443 13967 25449
rect 15194 25440 15200 25452
rect 15252 25440 15258 25492
rect 18046 25480 18052 25492
rect 18007 25452 18052 25480
rect 18046 25440 18052 25452
rect 18104 25440 18110 25492
rect 19518 25440 19524 25492
rect 19576 25480 19582 25492
rect 22373 25483 22431 25489
rect 19576 25452 21036 25480
rect 19576 25440 19582 25452
rect 2317 25415 2375 25421
rect 2317 25381 2329 25415
rect 2363 25412 2375 25415
rect 2958 25412 2964 25424
rect 2363 25384 2964 25412
rect 2363 25381 2375 25384
rect 2317 25375 2375 25381
rect 2958 25372 2964 25384
rect 3016 25372 3022 25424
rect 5721 25415 5779 25421
rect 5721 25381 5733 25415
rect 5767 25412 5779 25415
rect 6181 25415 6239 25421
rect 6181 25412 6193 25415
rect 5767 25384 6193 25412
rect 5767 25381 5779 25384
rect 5721 25375 5779 25381
rect 6181 25381 6193 25384
rect 6227 25381 6239 25415
rect 7929 25415 7987 25421
rect 6181 25375 6239 25381
rect 6472 25384 7420 25412
rect 2222 25344 2228 25356
rect 1688 25316 2228 25344
rect 1397 25279 1455 25285
rect 1397 25245 1409 25279
rect 1443 25276 1455 25279
rect 1486 25276 1492 25288
rect 1443 25248 1492 25276
rect 1443 25245 1455 25248
rect 1397 25239 1455 25245
rect 1486 25236 1492 25248
rect 1544 25236 1550 25288
rect 1688 25208 1716 25316
rect 2222 25304 2228 25316
rect 2280 25304 2286 25356
rect 2866 25344 2872 25356
rect 2827 25316 2872 25344
rect 2866 25304 2872 25316
rect 2924 25304 2930 25356
rect 6472 25344 6500 25384
rect 3988 25316 6500 25344
rect 3988 25276 4016 25316
rect 6546 25304 6552 25356
rect 6604 25344 6610 25356
rect 7285 25347 7343 25353
rect 7285 25344 7297 25347
rect 6604 25316 7297 25344
rect 6604 25304 6610 25316
rect 7285 25313 7297 25316
rect 7331 25313 7343 25347
rect 7392 25344 7420 25384
rect 7929 25381 7941 25415
rect 7975 25412 7987 25415
rect 8941 25415 8999 25421
rect 8941 25412 8953 25415
rect 7975 25384 8953 25412
rect 7975 25381 7987 25384
rect 7929 25375 7987 25381
rect 8941 25381 8953 25384
rect 8987 25381 8999 25415
rect 8941 25375 8999 25381
rect 9398 25372 9404 25424
rect 9456 25412 9462 25424
rect 9456 25384 14596 25412
rect 9456 25372 9462 25384
rect 9125 25347 9183 25353
rect 9125 25344 9137 25347
rect 7392 25316 9137 25344
rect 7285 25307 7343 25313
rect 9125 25313 9137 25316
rect 9171 25313 9183 25347
rect 9125 25307 9183 25313
rect 9214 25304 9220 25356
rect 9272 25344 9278 25356
rect 9272 25316 9317 25344
rect 9272 25304 9278 25316
rect 9766 25304 9772 25356
rect 9824 25344 9830 25356
rect 10594 25344 10600 25356
rect 9824 25316 10600 25344
rect 9824 25304 9830 25316
rect 10594 25304 10600 25316
rect 10652 25344 10658 25356
rect 12710 25344 12716 25356
rect 10652 25316 11008 25344
rect 10652 25304 10658 25316
rect 1504 25180 1716 25208
rect 1780 25248 4016 25276
rect 4065 25279 4123 25285
rect 1504 25152 1532 25180
rect 1780 25152 1808 25248
rect 4065 25245 4077 25279
rect 4111 25245 4123 25279
rect 4706 25276 4712 25288
rect 4667 25248 4712 25276
rect 4065 25239 4123 25245
rect 2222 25168 2228 25220
rect 2280 25208 2286 25220
rect 2777 25211 2835 25217
rect 2777 25208 2789 25211
rect 2280 25180 2789 25208
rect 2280 25168 2286 25180
rect 2777 25177 2789 25180
rect 2823 25177 2835 25211
rect 2777 25171 2835 25177
rect 3970 25168 3976 25220
rect 4028 25208 4034 25220
rect 4080 25208 4108 25239
rect 4706 25236 4712 25248
rect 4764 25236 4770 25288
rect 4982 25276 4988 25288
rect 4943 25248 4988 25276
rect 4982 25236 4988 25248
rect 5040 25236 5046 25288
rect 5074 25236 5080 25288
rect 5132 25276 5138 25288
rect 5169 25279 5227 25285
rect 5169 25276 5181 25279
rect 5132 25248 5181 25276
rect 5132 25236 5138 25248
rect 5169 25245 5181 25248
rect 5215 25276 5227 25279
rect 5905 25279 5963 25285
rect 5905 25276 5917 25279
rect 5215 25248 5917 25276
rect 5215 25245 5227 25248
rect 5169 25239 5227 25245
rect 5905 25245 5917 25248
rect 5951 25245 5963 25279
rect 5905 25239 5963 25245
rect 5997 25279 6055 25285
rect 5997 25245 6009 25279
rect 6043 25276 6055 25279
rect 6089 25279 6147 25285
rect 6089 25276 6101 25279
rect 6043 25248 6101 25276
rect 6043 25245 6055 25248
rect 5997 25239 6055 25245
rect 6089 25245 6101 25248
rect 6135 25245 6147 25279
rect 6089 25239 6147 25245
rect 6181 25279 6239 25285
rect 6181 25245 6193 25279
rect 6227 25276 6239 25279
rect 6457 25279 6515 25285
rect 6457 25276 6469 25279
rect 6227 25248 6469 25276
rect 6227 25245 6239 25248
rect 6181 25239 6239 25245
rect 6457 25245 6469 25248
rect 6503 25245 6515 25279
rect 7190 25276 7196 25288
rect 7151 25248 7196 25276
rect 6457 25239 6515 25245
rect 7190 25236 7196 25248
rect 7248 25236 7254 25288
rect 8202 25276 8208 25288
rect 8163 25248 8208 25276
rect 8202 25236 8208 25248
rect 8260 25236 8266 25288
rect 9306 25276 9312 25288
rect 9267 25248 9312 25276
rect 9306 25236 9312 25248
rect 9364 25236 9370 25288
rect 9398 25236 9404 25288
rect 9456 25276 9462 25288
rect 9456 25248 9501 25276
rect 9456 25236 9462 25248
rect 9674 25236 9680 25288
rect 9732 25276 9738 25288
rect 10980 25285 11008 25316
rect 11072 25316 12716 25344
rect 9953 25279 10011 25285
rect 9953 25276 9965 25279
rect 9732 25248 9965 25276
rect 9732 25236 9738 25248
rect 9953 25245 9965 25248
rect 9999 25245 10011 25279
rect 9953 25239 10011 25245
rect 10965 25279 11023 25285
rect 10965 25245 10977 25279
rect 11011 25245 11023 25279
rect 10965 25239 11023 25245
rect 4028 25180 4108 25208
rect 5721 25211 5779 25217
rect 4028 25168 4034 25180
rect 5721 25177 5733 25211
rect 5767 25208 5779 25211
rect 7929 25211 7987 25217
rect 7929 25208 7941 25211
rect 5767 25180 7941 25208
rect 5767 25177 5779 25180
rect 5721 25171 5779 25177
rect 7929 25177 7941 25180
rect 7975 25177 7987 25211
rect 9324 25208 9352 25236
rect 10045 25211 10103 25217
rect 10045 25208 10057 25211
rect 9324 25180 10057 25208
rect 7929 25171 7987 25177
rect 10045 25177 10057 25180
rect 10091 25177 10103 25211
rect 11072 25208 11100 25316
rect 12710 25304 12716 25316
rect 12768 25344 12774 25356
rect 12986 25344 12992 25356
rect 12768 25316 12992 25344
rect 12768 25304 12774 25316
rect 12986 25304 12992 25316
rect 13044 25304 13050 25356
rect 13265 25347 13323 25353
rect 13265 25344 13277 25347
rect 13096 25316 13277 25344
rect 11241 25279 11299 25285
rect 11241 25245 11253 25279
rect 11287 25245 11299 25279
rect 11422 25276 11428 25288
rect 11383 25248 11428 25276
rect 11241 25239 11299 25245
rect 10045 25171 10103 25177
rect 10152 25180 11100 25208
rect 1486 25100 1492 25152
rect 1544 25100 1550 25152
rect 1581 25143 1639 25149
rect 1581 25109 1593 25143
rect 1627 25140 1639 25143
rect 1762 25140 1768 25152
rect 1627 25112 1768 25140
rect 1627 25109 1639 25112
rect 1581 25103 1639 25109
rect 1762 25100 1768 25112
rect 1820 25100 1826 25152
rect 2685 25143 2743 25149
rect 2685 25109 2697 25143
rect 2731 25140 2743 25143
rect 3786 25140 3792 25152
rect 2731 25112 3792 25140
rect 2731 25109 2743 25112
rect 2685 25103 2743 25109
rect 3786 25100 3792 25112
rect 3844 25100 3850 25152
rect 4525 25143 4583 25149
rect 4525 25109 4537 25143
rect 4571 25140 4583 25143
rect 5166 25140 5172 25152
rect 4571 25112 5172 25140
rect 4571 25109 4583 25112
rect 4525 25103 4583 25109
rect 5166 25100 5172 25112
rect 5224 25100 5230 25152
rect 6549 25143 6607 25149
rect 6549 25109 6561 25143
rect 6595 25140 6607 25143
rect 10152 25140 10180 25180
rect 6595 25112 10180 25140
rect 6595 25109 6607 25112
rect 6549 25103 6607 25109
rect 10226 25100 10232 25152
rect 10284 25140 10290 25152
rect 10594 25140 10600 25152
rect 10284 25112 10600 25140
rect 10284 25100 10290 25112
rect 10594 25100 10600 25112
rect 10652 25100 10658 25152
rect 10781 25143 10839 25149
rect 10781 25109 10793 25143
rect 10827 25140 10839 25143
rect 10962 25140 10968 25152
rect 10827 25112 10968 25140
rect 10827 25109 10839 25112
rect 10781 25103 10839 25109
rect 10962 25100 10968 25112
rect 11020 25100 11026 25152
rect 11256 25140 11284 25239
rect 11422 25236 11428 25248
rect 11480 25236 11486 25288
rect 12066 25276 12072 25288
rect 11979 25248 12072 25276
rect 12066 25236 12072 25248
rect 12124 25276 12130 25288
rect 12250 25276 12256 25288
rect 12124 25248 12256 25276
rect 12124 25236 12130 25248
rect 12250 25236 12256 25248
rect 12308 25236 12314 25288
rect 12345 25279 12403 25285
rect 12345 25245 12357 25279
rect 12391 25245 12403 25279
rect 12526 25276 12532 25288
rect 12487 25248 12532 25276
rect 12345 25239 12403 25245
rect 11330 25168 11336 25220
rect 11388 25208 11394 25220
rect 11974 25208 11980 25220
rect 11388 25180 11980 25208
rect 11388 25168 11394 25180
rect 11974 25168 11980 25180
rect 12032 25168 12038 25220
rect 12360 25208 12388 25239
rect 12526 25236 12532 25248
rect 12584 25236 12590 25288
rect 12802 25236 12808 25288
rect 12860 25276 12866 25288
rect 13096 25276 13124 25316
rect 13265 25313 13277 25316
rect 13311 25313 13323 25347
rect 13265 25307 13323 25313
rect 13449 25347 13507 25353
rect 13449 25313 13461 25347
rect 13495 25344 13507 25347
rect 14093 25347 14151 25353
rect 14093 25344 14105 25347
rect 13495 25316 14105 25344
rect 13495 25313 13507 25316
rect 13449 25307 13507 25313
rect 14093 25313 14105 25316
rect 14139 25313 14151 25347
rect 14093 25307 14151 25313
rect 14568 25285 14596 25384
rect 15102 25372 15108 25424
rect 15160 25412 15166 25424
rect 15565 25415 15623 25421
rect 15565 25412 15577 25415
rect 15160 25384 15577 25412
rect 15160 25372 15166 25384
rect 15565 25381 15577 25384
rect 15611 25412 15623 25415
rect 16022 25412 16028 25424
rect 15611 25384 16028 25412
rect 15611 25381 15623 25384
rect 15565 25375 15623 25381
rect 16022 25372 16028 25384
rect 16080 25372 16086 25424
rect 17497 25415 17555 25421
rect 17497 25381 17509 25415
rect 17543 25412 17555 25415
rect 20898 25412 20904 25424
rect 17543 25384 20904 25412
rect 17543 25381 17555 25384
rect 17497 25375 17555 25381
rect 20898 25372 20904 25384
rect 20956 25372 20962 25424
rect 21008 25412 21036 25452
rect 22373 25449 22385 25483
rect 22419 25480 22431 25483
rect 23750 25480 23756 25492
rect 22419 25452 23756 25480
rect 22419 25449 22431 25452
rect 22373 25443 22431 25449
rect 23750 25440 23756 25452
rect 23808 25440 23814 25492
rect 24486 25440 24492 25492
rect 24544 25480 24550 25492
rect 24765 25483 24823 25489
rect 24765 25480 24777 25483
rect 24544 25452 24777 25480
rect 24544 25440 24550 25452
rect 24765 25449 24777 25452
rect 24811 25449 24823 25483
rect 24765 25443 24823 25449
rect 31202 25440 31208 25492
rect 31260 25480 31266 25492
rect 31297 25483 31355 25489
rect 31297 25480 31309 25483
rect 31260 25452 31309 25480
rect 31260 25440 31266 25452
rect 31297 25449 31309 25452
rect 31343 25449 31355 25483
rect 31297 25443 31355 25449
rect 27154 25412 27160 25424
rect 21008 25384 27160 25412
rect 27154 25372 27160 25384
rect 27212 25372 27218 25424
rect 15286 25304 15292 25356
rect 15344 25344 15350 25356
rect 15657 25347 15715 25353
rect 15344 25316 15516 25344
rect 15344 25304 15350 25316
rect 12860 25248 13124 25276
rect 13173 25279 13231 25285
rect 12860 25236 12866 25248
rect 13173 25245 13185 25279
rect 13219 25245 13231 25279
rect 13173 25239 13231 25245
rect 13357 25279 13415 25285
rect 13357 25245 13369 25279
rect 13403 25276 13415 25279
rect 13909 25279 13967 25285
rect 13403 25248 13860 25276
rect 13403 25245 13415 25248
rect 13357 25239 13415 25245
rect 13188 25208 13216 25239
rect 13630 25208 13636 25220
rect 12360 25180 13032 25208
rect 13188 25180 13636 25208
rect 11606 25140 11612 25152
rect 11256 25112 11612 25140
rect 11606 25100 11612 25112
rect 11664 25100 11670 25152
rect 11885 25143 11943 25149
rect 11885 25109 11897 25143
rect 11931 25140 11943 25143
rect 12342 25140 12348 25152
rect 11931 25112 12348 25140
rect 11931 25109 11943 25112
rect 11885 25103 11943 25109
rect 12342 25100 12348 25112
rect 12400 25100 12406 25152
rect 13004 25140 13032 25180
rect 13630 25168 13636 25180
rect 13688 25168 13694 25220
rect 13170 25140 13176 25152
rect 13004 25112 13176 25140
rect 13170 25100 13176 25112
rect 13228 25100 13234 25152
rect 13832 25140 13860 25248
rect 13909 25245 13921 25279
rect 13955 25276 13967 25279
rect 14369 25279 14427 25285
rect 14369 25276 14381 25279
rect 13955 25248 14381 25276
rect 13955 25245 13967 25248
rect 13909 25239 13967 25245
rect 14369 25245 14381 25248
rect 14415 25245 14427 25279
rect 14369 25239 14427 25245
rect 14461 25279 14519 25285
rect 14461 25245 14473 25279
rect 14507 25245 14519 25279
rect 14461 25239 14519 25245
rect 14553 25279 14611 25285
rect 14553 25245 14565 25279
rect 14599 25245 14611 25279
rect 14734 25276 14740 25288
rect 14695 25248 14740 25276
rect 14553 25239 14611 25245
rect 13998 25168 14004 25220
rect 14056 25208 14062 25220
rect 14476 25208 14504 25239
rect 14734 25236 14740 25248
rect 14792 25236 14798 25288
rect 15378 25276 15384 25288
rect 15339 25248 15384 25276
rect 15378 25236 15384 25248
rect 15436 25236 15442 25288
rect 15488 25276 15516 25316
rect 15657 25313 15669 25347
rect 15703 25344 15715 25347
rect 16390 25344 16396 25356
rect 15703 25316 16396 25344
rect 15703 25313 15715 25316
rect 15657 25307 15715 25313
rect 16390 25304 16396 25316
rect 16448 25304 16454 25356
rect 19245 25347 19303 25353
rect 19245 25344 19257 25347
rect 18248 25316 19257 25344
rect 18248 25285 18276 25316
rect 19245 25313 19257 25316
rect 19291 25313 19303 25347
rect 20622 25344 20628 25356
rect 19245 25307 19303 25313
rect 19720 25316 20628 25344
rect 19720 25288 19748 25316
rect 20622 25304 20628 25316
rect 20680 25344 20686 25356
rect 22462 25344 22468 25356
rect 20680 25316 22468 25344
rect 20680 25304 20686 25316
rect 17221 25279 17279 25285
rect 17221 25276 17233 25279
rect 15488 25248 17233 25276
rect 17221 25245 17233 25248
rect 17267 25245 17279 25279
rect 17221 25239 17279 25245
rect 18233 25279 18291 25285
rect 18233 25245 18245 25279
rect 18279 25245 18291 25279
rect 18414 25276 18420 25288
rect 18375 25248 18420 25276
rect 18233 25239 18291 25245
rect 18414 25236 18420 25248
rect 18472 25236 18478 25288
rect 18509 25279 18567 25285
rect 18509 25245 18521 25279
rect 18555 25245 18567 25279
rect 19426 25276 19432 25288
rect 19387 25248 19432 25276
rect 18509 25239 18567 25245
rect 15746 25208 15752 25220
rect 14056 25180 15752 25208
rect 14056 25168 14062 25180
rect 15746 25168 15752 25180
rect 15804 25168 15810 25220
rect 16298 25208 16304 25220
rect 16259 25180 16304 25208
rect 16298 25168 16304 25180
rect 16356 25168 16362 25220
rect 16666 25208 16672 25220
rect 16408 25180 16672 25208
rect 16408 25140 16436 25180
rect 16666 25168 16672 25180
rect 16724 25168 16730 25220
rect 18322 25168 18328 25220
rect 18380 25208 18386 25220
rect 18524 25208 18552 25239
rect 19426 25236 19432 25248
rect 19484 25236 19490 25288
rect 19702 25276 19708 25288
rect 19615 25248 19708 25276
rect 19702 25236 19708 25248
rect 19760 25236 19766 25288
rect 21376 25285 21404 25316
rect 22462 25304 22468 25316
rect 22520 25304 22526 25356
rect 22741 25347 22799 25353
rect 22741 25313 22753 25347
rect 22787 25344 22799 25347
rect 24762 25344 24768 25356
rect 22787 25316 24768 25344
rect 22787 25313 22799 25316
rect 22741 25307 22799 25313
rect 24762 25304 24768 25316
rect 24820 25304 24826 25356
rect 19889 25279 19947 25285
rect 19889 25245 19901 25279
rect 19935 25245 19947 25279
rect 19889 25239 19947 25245
rect 21085 25279 21143 25285
rect 21085 25245 21097 25279
rect 21131 25245 21143 25279
rect 21085 25239 21143 25245
rect 21361 25279 21419 25285
rect 21361 25245 21373 25279
rect 21407 25245 21419 25279
rect 21361 25239 21419 25245
rect 21545 25279 21603 25285
rect 21545 25245 21557 25279
rect 21591 25276 21603 25279
rect 22094 25276 22100 25288
rect 21591 25248 22100 25276
rect 21591 25245 21603 25248
rect 21545 25239 21603 25245
rect 18380 25180 18552 25208
rect 18380 25168 18386 25180
rect 18690 25168 18696 25220
rect 18748 25208 18754 25220
rect 19904 25208 19932 25239
rect 18748 25180 19932 25208
rect 21100 25208 21128 25239
rect 22094 25236 22100 25248
rect 22152 25236 22158 25288
rect 22554 25276 22560 25288
rect 22515 25248 22560 25276
rect 22554 25236 22560 25248
rect 22612 25236 22618 25288
rect 22833 25279 22891 25285
rect 22833 25245 22845 25279
rect 22879 25276 22891 25279
rect 23382 25276 23388 25288
rect 22879 25248 23388 25276
rect 22879 25245 22891 25248
rect 22833 25239 22891 25245
rect 23382 25236 23388 25248
rect 23440 25236 23446 25288
rect 23845 25279 23903 25285
rect 23845 25245 23857 25279
rect 23891 25276 23903 25279
rect 25041 25279 25099 25285
rect 25041 25276 25053 25279
rect 23891 25248 25053 25276
rect 23891 25245 23903 25248
rect 23845 25239 23903 25245
rect 25041 25245 25053 25248
rect 25087 25245 25099 25279
rect 25041 25239 25099 25245
rect 25222 25236 25228 25288
rect 25280 25276 25286 25288
rect 25961 25279 26019 25285
rect 25961 25276 25973 25279
rect 25280 25248 25973 25276
rect 25280 25236 25286 25248
rect 25961 25245 25973 25248
rect 26007 25245 26019 25279
rect 25961 25239 26019 25245
rect 26237 25279 26295 25285
rect 26237 25245 26249 25279
rect 26283 25276 26295 25279
rect 26326 25276 26332 25288
rect 26283 25248 26332 25276
rect 26283 25245 26295 25248
rect 26237 25239 26295 25245
rect 26326 25236 26332 25248
rect 26384 25236 26390 25288
rect 26421 25279 26479 25285
rect 26421 25245 26433 25279
rect 26467 25276 26479 25279
rect 26510 25276 26516 25288
rect 26467 25248 26516 25276
rect 26467 25245 26479 25248
rect 26421 25239 26479 25245
rect 26510 25236 26516 25248
rect 26568 25236 26574 25288
rect 27157 25279 27215 25285
rect 27157 25245 27169 25279
rect 27203 25276 27215 25279
rect 28258 25276 28264 25288
rect 27203 25248 28264 25276
rect 27203 25245 27215 25248
rect 27157 25239 27215 25245
rect 28258 25236 28264 25248
rect 28316 25236 28322 25288
rect 29917 25279 29975 25285
rect 29917 25276 29929 25279
rect 28460 25248 29929 25276
rect 21634 25208 21640 25220
rect 21100 25180 21640 25208
rect 18748 25168 18754 25180
rect 21634 25168 21640 25180
rect 21692 25168 21698 25220
rect 23477 25211 23535 25217
rect 23477 25177 23489 25211
rect 23523 25208 23535 25211
rect 24118 25208 24124 25220
rect 23523 25180 24124 25208
rect 23523 25177 23535 25180
rect 23477 25171 23535 25177
rect 24118 25168 24124 25180
rect 24176 25168 24182 25220
rect 24397 25211 24455 25217
rect 24397 25208 24409 25211
rect 24228 25180 24409 25208
rect 13832 25112 16436 25140
rect 16482 25100 16488 25152
rect 16540 25140 16546 25152
rect 16577 25143 16635 25149
rect 16577 25140 16589 25143
rect 16540 25112 16589 25140
rect 16540 25100 16546 25112
rect 16577 25109 16589 25112
rect 16623 25109 16635 25143
rect 16684 25140 16712 25168
rect 20254 25140 20260 25152
rect 16684 25112 20260 25140
rect 16577 25103 16635 25109
rect 20254 25100 20260 25112
rect 20312 25100 20318 25152
rect 20901 25143 20959 25149
rect 20901 25109 20913 25143
rect 20947 25140 20959 25143
rect 20990 25140 20996 25152
rect 20947 25112 20996 25140
rect 20947 25109 20959 25112
rect 20901 25103 20959 25109
rect 20990 25100 20996 25112
rect 21048 25100 21054 25152
rect 22462 25100 22468 25152
rect 22520 25140 22526 25152
rect 23385 25143 23443 25149
rect 23385 25140 23397 25143
rect 22520 25112 23397 25140
rect 22520 25100 22526 25112
rect 23385 25109 23397 25112
rect 23431 25109 23443 25143
rect 23566 25140 23572 25152
rect 23527 25112 23572 25140
rect 23385 25103 23443 25109
rect 23566 25100 23572 25112
rect 23624 25100 23630 25152
rect 23661 25143 23719 25149
rect 23661 25109 23673 25143
rect 23707 25140 23719 25143
rect 24228 25140 24256 25180
rect 24397 25177 24409 25180
rect 24443 25208 24455 25211
rect 24946 25208 24952 25220
rect 24443 25180 24952 25208
rect 24443 25177 24455 25180
rect 24397 25171 24455 25177
rect 24946 25168 24952 25180
rect 25004 25168 25010 25220
rect 23707 25112 24256 25140
rect 23707 25109 23719 25112
rect 23661 25103 23719 25109
rect 24302 25100 24308 25152
rect 24360 25140 24366 25152
rect 24774 25143 24832 25149
rect 24774 25140 24786 25143
rect 24360 25112 24786 25140
rect 24360 25100 24366 25112
rect 24774 25109 24786 25112
rect 24820 25140 24832 25143
rect 25314 25140 25320 25152
rect 24820 25112 25320 25140
rect 24820 25109 24832 25112
rect 24774 25103 24832 25109
rect 25314 25100 25320 25112
rect 25372 25100 25378 25152
rect 25777 25143 25835 25149
rect 25777 25109 25789 25143
rect 25823 25140 25835 25143
rect 27154 25140 27160 25152
rect 25823 25112 27160 25140
rect 25823 25109 25835 25112
rect 25777 25103 25835 25109
rect 27154 25100 27160 25112
rect 27212 25100 27218 25152
rect 27798 25100 27804 25152
rect 27856 25140 27862 25152
rect 28460 25149 28488 25248
rect 29917 25245 29929 25248
rect 29963 25245 29975 25279
rect 29917 25239 29975 25245
rect 30184 25211 30242 25217
rect 30184 25177 30196 25211
rect 30230 25208 30242 25211
rect 30282 25208 30288 25220
rect 30230 25180 30288 25208
rect 30230 25177 30242 25180
rect 30184 25171 30242 25177
rect 30282 25168 30288 25180
rect 30340 25168 30346 25220
rect 28445 25143 28503 25149
rect 28445 25140 28457 25143
rect 27856 25112 28457 25140
rect 27856 25100 27862 25112
rect 28445 25109 28457 25112
rect 28491 25109 28503 25143
rect 28445 25103 28503 25109
rect 1104 25050 32016 25072
rect 1104 24998 7288 25050
rect 7340 24998 17592 25050
rect 17644 24998 27896 25050
rect 27948 24998 32016 25050
rect 1104 24976 32016 24998
rect 2133 24939 2191 24945
rect 2133 24905 2145 24939
rect 2179 24936 2191 24939
rect 2222 24936 2228 24948
rect 2179 24908 2228 24936
rect 2179 24905 2191 24908
rect 2133 24899 2191 24905
rect 2222 24896 2228 24908
rect 2280 24896 2286 24948
rect 5074 24896 5080 24948
rect 5132 24936 5138 24948
rect 5445 24939 5503 24945
rect 5445 24936 5457 24939
rect 5132 24908 5457 24936
rect 5132 24896 5138 24908
rect 5445 24905 5457 24908
rect 5491 24905 5503 24939
rect 5445 24899 5503 24905
rect 6362 24896 6368 24948
rect 6420 24896 6426 24948
rect 7190 24896 7196 24948
rect 7248 24936 7254 24948
rect 9398 24936 9404 24948
rect 7248 24908 9404 24936
rect 7248 24896 7254 24908
rect 9398 24896 9404 24908
rect 9456 24896 9462 24948
rect 9508 24908 10364 24936
rect 1670 24868 1676 24880
rect 1631 24840 1676 24868
rect 1670 24828 1676 24840
rect 1728 24828 1734 24880
rect 2590 24828 2596 24880
rect 2648 24828 2654 24880
rect 4430 24868 4436 24880
rect 3160 24840 4436 24868
rect 2222 24760 2228 24812
rect 2280 24800 2286 24812
rect 2608 24800 2636 24828
rect 2958 24800 2964 24812
rect 2280 24772 2636 24800
rect 2919 24772 2964 24800
rect 2280 24760 2286 24772
rect 2958 24760 2964 24772
rect 3016 24760 3022 24812
rect 3160 24809 3188 24840
rect 4430 24828 4436 24840
rect 4488 24828 4494 24880
rect 6380 24868 6408 24896
rect 9508 24868 9536 24908
rect 6380 24840 9536 24868
rect 9582 24828 9588 24880
rect 9640 24868 9646 24880
rect 10336 24877 10364 24908
rect 10594 24896 10600 24948
rect 10652 24936 10658 24948
rect 11790 24936 11796 24948
rect 10652 24908 11796 24936
rect 10652 24896 10658 24908
rect 11790 24896 11796 24908
rect 11848 24896 11854 24948
rect 12158 24896 12164 24948
rect 12216 24936 12222 24948
rect 16482 24936 16488 24948
rect 12216 24908 16488 24936
rect 12216 24896 12222 24908
rect 16482 24896 16488 24908
rect 16540 24896 16546 24948
rect 18046 24896 18052 24948
rect 18104 24936 18110 24948
rect 18414 24936 18420 24948
rect 18104 24908 18420 24936
rect 18104 24896 18110 24908
rect 18414 24896 18420 24908
rect 18472 24936 18478 24948
rect 19242 24936 19248 24948
rect 18472 24908 19248 24936
rect 18472 24896 18478 24908
rect 19242 24896 19248 24908
rect 19300 24896 19306 24948
rect 22186 24945 22192 24948
rect 22179 24939 22192 24945
rect 22179 24905 22191 24939
rect 22244 24936 22250 24948
rect 22244 24908 22279 24936
rect 22179 24899 22192 24905
rect 22186 24896 22192 24899
rect 22244 24896 22250 24908
rect 22554 24896 22560 24948
rect 22612 24936 22618 24948
rect 22612 24908 22876 24936
rect 22612 24896 22618 24908
rect 10321 24871 10379 24877
rect 9640 24840 10088 24868
rect 9640 24828 9646 24840
rect 3145 24803 3203 24809
rect 3145 24769 3157 24803
rect 3191 24769 3203 24803
rect 3145 24763 3203 24769
rect 4332 24803 4390 24809
rect 4332 24769 4344 24803
rect 4378 24800 4390 24803
rect 4890 24800 4896 24812
rect 4378 24772 4896 24800
rect 4378 24769 4390 24772
rect 4332 24763 4390 24769
rect 4890 24760 4896 24772
rect 4948 24760 4954 24812
rect 6362 24800 6368 24812
rect 6323 24772 6368 24800
rect 6362 24760 6368 24772
rect 6420 24760 6426 24812
rect 6549 24803 6607 24809
rect 6549 24769 6561 24803
rect 6595 24769 6607 24803
rect 6549 24763 6607 24769
rect 2590 24692 2596 24744
rect 2648 24732 2654 24744
rect 2869 24735 2927 24741
rect 2869 24732 2881 24735
rect 2648 24704 2881 24732
rect 2648 24692 2654 24704
rect 2869 24701 2881 24704
rect 2915 24701 2927 24735
rect 2869 24695 2927 24701
rect 3510 24692 3516 24744
rect 3568 24732 3574 24744
rect 3605 24735 3663 24741
rect 3605 24732 3617 24735
rect 3568 24704 3617 24732
rect 3568 24692 3574 24704
rect 3605 24701 3617 24704
rect 3651 24701 3663 24735
rect 3605 24695 3663 24701
rect 4065 24735 4123 24741
rect 4065 24701 4077 24735
rect 4111 24701 4123 24735
rect 6564 24732 6592 24763
rect 6638 24760 6644 24812
rect 6696 24800 6702 24812
rect 6696 24772 6741 24800
rect 6696 24760 6702 24772
rect 6822 24760 6828 24812
rect 6880 24800 6886 24812
rect 7101 24803 7159 24809
rect 7101 24800 7113 24803
rect 6880 24772 7113 24800
rect 6880 24760 6886 24772
rect 7101 24769 7113 24772
rect 7147 24769 7159 24803
rect 7101 24763 7159 24769
rect 7368 24803 7426 24809
rect 7368 24769 7380 24803
rect 7414 24800 7426 24803
rect 8202 24800 8208 24812
rect 7414 24772 8208 24800
rect 7414 24769 7426 24772
rect 7368 24763 7426 24769
rect 8202 24760 8208 24772
rect 8260 24760 8266 24812
rect 8662 24760 8668 24812
rect 8720 24800 8726 24812
rect 8941 24803 8999 24809
rect 8941 24800 8953 24803
rect 8720 24772 8953 24800
rect 8720 24760 8726 24772
rect 8941 24769 8953 24772
rect 8987 24769 8999 24803
rect 8941 24763 8999 24769
rect 8956 24732 8984 24763
rect 9122 24760 9128 24812
rect 9180 24800 9186 24812
rect 9309 24803 9367 24809
rect 9309 24800 9321 24803
rect 9180 24772 9321 24800
rect 9180 24760 9186 24772
rect 9309 24769 9321 24772
rect 9355 24769 9367 24803
rect 9309 24763 9367 24769
rect 9398 24760 9404 24812
rect 9456 24800 9462 24812
rect 10060 24809 10088 24840
rect 10321 24837 10333 24871
rect 10367 24837 10379 24871
rect 10321 24831 10379 24837
rect 10410 24828 10416 24880
rect 10468 24868 10474 24880
rect 10778 24868 10784 24880
rect 10468 24840 10784 24868
rect 10468 24828 10474 24840
rect 10778 24828 10784 24840
rect 10836 24828 10842 24880
rect 11514 24828 11520 24880
rect 11572 24868 11578 24880
rect 13078 24877 13084 24880
rect 13072 24868 13084 24877
rect 11572 24840 12848 24868
rect 13039 24840 13084 24868
rect 11572 24828 11578 24840
rect 9677 24803 9735 24809
rect 9677 24800 9689 24803
rect 9456 24772 9689 24800
rect 9456 24760 9462 24772
rect 9677 24769 9689 24772
rect 9723 24769 9735 24803
rect 9677 24763 9735 24769
rect 10045 24803 10103 24809
rect 10045 24769 10057 24803
rect 10091 24769 10103 24803
rect 11606 24800 11612 24812
rect 10045 24763 10103 24769
rect 10336 24772 11612 24800
rect 10336 24744 10364 24772
rect 11606 24760 11612 24772
rect 11664 24800 11670 24812
rect 11793 24803 11851 24809
rect 11793 24800 11805 24803
rect 11664 24772 11805 24800
rect 11664 24760 11670 24772
rect 11793 24769 11805 24772
rect 11839 24769 11851 24803
rect 11793 24763 11851 24769
rect 12820 24744 12848 24840
rect 13072 24831 13084 24840
rect 13078 24828 13084 24831
rect 13136 24828 13142 24880
rect 14918 24868 14924 24880
rect 14879 24840 14924 24868
rect 14918 24828 14924 24840
rect 14976 24828 14982 24880
rect 15470 24828 15476 24880
rect 15528 24868 15534 24880
rect 15654 24868 15660 24880
rect 15528 24840 15660 24868
rect 15528 24828 15534 24840
rect 15654 24828 15660 24840
rect 15712 24868 15718 24880
rect 16117 24871 16175 24877
rect 16117 24868 16129 24871
rect 15712 24840 16129 24868
rect 15712 24828 15718 24840
rect 16117 24837 16129 24840
rect 16163 24837 16175 24871
rect 16117 24831 16175 24837
rect 16206 24828 16212 24880
rect 16264 24868 16270 24880
rect 22462 24868 22468 24880
rect 16264 24840 22468 24868
rect 16264 24828 16270 24840
rect 22462 24828 22468 24840
rect 22520 24828 22526 24880
rect 22646 24868 22652 24880
rect 22607 24840 22652 24868
rect 22646 24828 22652 24840
rect 22704 24828 22710 24880
rect 13630 24760 13636 24812
rect 13688 24800 13694 24812
rect 13688 24772 13860 24800
rect 13688 24760 13694 24772
rect 6564 24704 7144 24732
rect 8956 24704 9674 24732
rect 4065 24695 4123 24701
rect 1946 24664 1952 24676
rect 1907 24636 1952 24664
rect 1946 24624 1952 24636
rect 2004 24624 2010 24676
rect 4080 24596 4108 24695
rect 6822 24664 6828 24676
rect 5000 24636 6828 24664
rect 5000 24596 5028 24636
rect 6822 24624 6828 24636
rect 6880 24624 6886 24676
rect 4080 24568 5028 24596
rect 6365 24599 6423 24605
rect 6365 24565 6377 24599
rect 6411 24596 6423 24599
rect 6546 24596 6552 24608
rect 6411 24568 6552 24596
rect 6411 24565 6423 24568
rect 6365 24559 6423 24565
rect 6546 24556 6552 24568
rect 6604 24556 6610 24608
rect 7116 24596 7144 24704
rect 9306 24664 9312 24676
rect 8404 24636 9312 24664
rect 8404 24596 8432 24636
rect 9306 24624 9312 24636
rect 9364 24624 9370 24676
rect 9646 24664 9674 24704
rect 10318 24692 10324 24744
rect 10376 24692 10382 24744
rect 10502 24692 10508 24744
rect 10560 24732 10566 24744
rect 11517 24735 11575 24741
rect 11517 24732 11529 24735
rect 10560 24704 11529 24732
rect 10560 24692 10566 24704
rect 11517 24701 11529 24704
rect 11563 24701 11575 24735
rect 12802 24732 12808 24744
rect 12763 24704 12808 24732
rect 11517 24695 11575 24701
rect 12802 24692 12808 24704
rect 12860 24692 12866 24744
rect 13832 24732 13860 24772
rect 14458 24760 14464 24812
rect 14516 24800 14522 24812
rect 14737 24803 14795 24809
rect 14737 24800 14749 24803
rect 14516 24772 14749 24800
rect 14516 24760 14522 24772
rect 14737 24769 14749 24772
rect 14783 24769 14795 24803
rect 14737 24763 14795 24769
rect 15933 24803 15991 24809
rect 15933 24769 15945 24803
rect 15979 24800 15991 24803
rect 16853 24803 16911 24809
rect 16853 24800 16865 24803
rect 15979 24772 16865 24800
rect 15979 24769 15991 24772
rect 15933 24763 15991 24769
rect 16853 24769 16865 24772
rect 16899 24800 16911 24803
rect 16942 24800 16948 24812
rect 16899 24772 16948 24800
rect 16899 24769 16911 24772
rect 16853 24763 16911 24769
rect 16942 24760 16948 24772
rect 17000 24760 17006 24812
rect 18322 24760 18328 24812
rect 18380 24800 18386 24812
rect 18509 24803 18567 24809
rect 18509 24800 18521 24803
rect 18380 24772 18521 24800
rect 18380 24760 18386 24772
rect 18509 24769 18521 24772
rect 18555 24769 18567 24803
rect 18509 24763 18567 24769
rect 18693 24803 18751 24809
rect 18693 24769 18705 24803
rect 18739 24769 18751 24803
rect 18693 24763 18751 24769
rect 18785 24803 18843 24809
rect 18785 24769 18797 24803
rect 18831 24800 18843 24803
rect 18877 24803 18935 24809
rect 18877 24800 18889 24803
rect 18831 24772 18889 24800
rect 18831 24769 18843 24772
rect 18785 24763 18843 24769
rect 18877 24769 18889 24772
rect 18923 24769 18935 24803
rect 19426 24800 19432 24812
rect 19387 24772 19432 24800
rect 18877 24763 18935 24769
rect 13832 24704 14780 24732
rect 14752 24664 14780 24704
rect 16022 24692 16028 24744
rect 16080 24732 16086 24744
rect 16209 24735 16267 24741
rect 16209 24732 16221 24735
rect 16080 24704 16221 24732
rect 16080 24692 16086 24704
rect 16209 24701 16221 24704
rect 16255 24701 16267 24735
rect 16209 24695 16267 24701
rect 17129 24735 17187 24741
rect 17129 24701 17141 24735
rect 17175 24732 17187 24735
rect 17310 24732 17316 24744
rect 17175 24704 17316 24732
rect 17175 24701 17187 24704
rect 17129 24695 17187 24701
rect 17310 24692 17316 24704
rect 17368 24692 17374 24744
rect 18708 24732 18736 24763
rect 19426 24760 19432 24772
rect 19484 24760 19490 24812
rect 19702 24800 19708 24812
rect 19663 24772 19708 24800
rect 19702 24760 19708 24772
rect 19760 24760 19766 24812
rect 19889 24803 19947 24809
rect 19889 24769 19901 24803
rect 19935 24769 19947 24803
rect 20990 24800 20996 24812
rect 20951 24772 20996 24800
rect 19889 24763 19947 24769
rect 19794 24732 19800 24744
rect 18708 24704 19800 24732
rect 19794 24692 19800 24704
rect 19852 24732 19858 24744
rect 19904 24732 19932 24763
rect 20990 24760 20996 24772
rect 21048 24760 21054 24812
rect 21082 24760 21088 24812
rect 21140 24800 21146 24812
rect 21177 24803 21235 24809
rect 21177 24800 21189 24803
rect 21140 24772 21189 24800
rect 21140 24760 21146 24772
rect 21177 24769 21189 24772
rect 21223 24769 21235 24803
rect 21177 24763 21235 24769
rect 22094 24760 22100 24812
rect 22152 24800 22158 24812
rect 22741 24803 22799 24809
rect 22741 24800 22753 24803
rect 22152 24772 22753 24800
rect 22152 24760 22158 24772
rect 22741 24769 22753 24772
rect 22787 24769 22799 24803
rect 22848 24800 22876 24908
rect 24121 24871 24179 24877
rect 24121 24837 24133 24871
rect 24167 24868 24179 24871
rect 24670 24868 24676 24880
rect 24167 24840 24676 24868
rect 24167 24837 24179 24840
rect 24121 24831 24179 24837
rect 24670 24828 24676 24840
rect 24728 24828 24734 24880
rect 26510 24868 26516 24880
rect 25608 24840 26516 24868
rect 23290 24800 23296 24812
rect 22848 24772 23296 24800
rect 22741 24763 22799 24769
rect 23290 24760 23296 24772
rect 23348 24760 23354 24812
rect 23474 24800 23480 24812
rect 23435 24772 23480 24800
rect 23474 24760 23480 24772
rect 23532 24760 23538 24812
rect 24305 24803 24363 24809
rect 24305 24769 24317 24803
rect 24351 24800 24363 24803
rect 25041 24803 25099 24809
rect 25041 24800 25053 24803
rect 24351 24772 25053 24800
rect 24351 24769 24363 24772
rect 24305 24763 24363 24769
rect 25041 24769 25053 24772
rect 25087 24769 25099 24803
rect 25222 24800 25228 24812
rect 25183 24772 25228 24800
rect 25041 24763 25099 24769
rect 25222 24760 25228 24772
rect 25280 24760 25286 24812
rect 25498 24800 25504 24812
rect 25459 24772 25504 24800
rect 25498 24760 25504 24772
rect 25556 24760 25562 24812
rect 19852 24704 19932 24732
rect 21269 24735 21327 24741
rect 19852 24692 19858 24704
rect 21269 24701 21281 24735
rect 21315 24732 21327 24735
rect 22554 24732 22560 24744
rect 21315 24704 22560 24732
rect 21315 24701 21327 24704
rect 21269 24695 21327 24701
rect 22554 24692 22560 24704
rect 22612 24692 22618 24744
rect 22649 24735 22707 24741
rect 22649 24701 22661 24735
rect 22695 24732 22707 24735
rect 22695 24704 22764 24732
rect 22695 24701 22707 24704
rect 22649 24695 22707 24701
rect 15930 24664 15936 24676
rect 9646 24636 10640 24664
rect 14752 24636 15936 24664
rect 7116 24568 8432 24596
rect 8478 24556 8484 24608
rect 8536 24596 8542 24608
rect 9122 24596 9128 24608
rect 8536 24568 9128 24596
rect 8536 24556 8542 24568
rect 9122 24556 9128 24568
rect 9180 24556 9186 24608
rect 10612 24596 10640 24636
rect 15930 24624 15936 24636
rect 15988 24664 15994 24676
rect 17862 24664 17868 24676
rect 15988 24636 17868 24664
rect 15988 24624 15994 24636
rect 17862 24624 17868 24636
rect 17920 24624 17926 24676
rect 18325 24667 18383 24673
rect 18325 24633 18337 24667
rect 18371 24664 18383 24667
rect 22002 24664 22008 24676
rect 18371 24636 22008 24664
rect 18371 24633 18383 24636
rect 18325 24627 18383 24633
rect 22002 24624 22008 24636
rect 22060 24624 22066 24676
rect 22736 24664 22764 24704
rect 23382 24692 23388 24744
rect 23440 24732 23446 24744
rect 24581 24735 24639 24741
rect 23440 24704 24532 24732
rect 23440 24692 23446 24704
rect 23661 24667 23719 24673
rect 23661 24664 23673 24667
rect 22736 24636 23673 24664
rect 23661 24633 23673 24636
rect 23707 24633 23719 24667
rect 24504 24664 24532 24704
rect 24581 24701 24593 24735
rect 24627 24732 24639 24735
rect 25608 24732 25636 24840
rect 26510 24828 26516 24840
rect 26568 24828 26574 24880
rect 29656 24840 30512 24868
rect 25685 24803 25743 24809
rect 25685 24769 25697 24803
rect 25731 24769 25743 24803
rect 25685 24763 25743 24769
rect 26237 24803 26295 24809
rect 26237 24769 26249 24803
rect 26283 24800 26295 24803
rect 26786 24800 26792 24812
rect 26283 24772 26792 24800
rect 26283 24769 26295 24772
rect 26237 24763 26295 24769
rect 24627 24704 25636 24732
rect 24627 24701 24639 24704
rect 24581 24695 24639 24701
rect 25700 24664 25728 24763
rect 26786 24760 26792 24772
rect 26844 24760 26850 24812
rect 26970 24800 26976 24812
rect 26931 24772 26976 24800
rect 26970 24760 26976 24772
rect 27028 24760 27034 24812
rect 27154 24800 27160 24812
rect 27115 24772 27160 24800
rect 27154 24760 27160 24772
rect 27212 24760 27218 24812
rect 27430 24800 27436 24812
rect 27391 24772 27436 24800
rect 27430 24760 27436 24772
rect 27488 24760 27494 24812
rect 28077 24803 28135 24809
rect 28077 24769 28089 24803
rect 28123 24800 28135 24803
rect 28166 24800 28172 24812
rect 28123 24772 28172 24800
rect 28123 24769 28135 24772
rect 28077 24763 28135 24769
rect 28166 24760 28172 24772
rect 28224 24760 28230 24812
rect 29086 24800 29092 24812
rect 29047 24772 29092 24800
rect 29086 24760 29092 24772
rect 29144 24760 29150 24812
rect 29273 24803 29331 24809
rect 29273 24769 29285 24803
rect 29319 24769 29331 24803
rect 29273 24763 29331 24769
rect 29549 24803 29607 24809
rect 29549 24769 29561 24803
rect 29595 24800 29607 24803
rect 29656 24800 29684 24840
rect 29595 24772 29684 24800
rect 29595 24769 29607 24772
rect 29549 24763 29607 24769
rect 26421 24735 26479 24741
rect 26421 24701 26433 24735
rect 26467 24732 26479 24735
rect 27341 24735 27399 24741
rect 27341 24732 27353 24735
rect 26467 24704 27353 24732
rect 26467 24701 26479 24704
rect 26421 24695 26479 24701
rect 27341 24701 27353 24704
rect 27387 24701 27399 24735
rect 27341 24695 27399 24701
rect 25866 24664 25872 24676
rect 24504 24636 25872 24664
rect 23661 24627 23719 24633
rect 25866 24624 25872 24636
rect 25924 24624 25930 24676
rect 14090 24596 14096 24608
rect 10612 24568 14096 24596
rect 14090 24556 14096 24568
rect 14148 24556 14154 24608
rect 14182 24556 14188 24608
rect 14240 24596 14246 24608
rect 14240 24568 14285 24596
rect 14240 24556 14246 24568
rect 14918 24556 14924 24608
rect 14976 24596 14982 24608
rect 18506 24596 18512 24608
rect 14976 24568 18512 24596
rect 14976 24556 14982 24568
rect 18506 24556 18512 24568
rect 18564 24596 18570 24608
rect 18877 24599 18935 24605
rect 18877 24596 18889 24599
rect 18564 24568 18889 24596
rect 18564 24556 18570 24568
rect 18877 24565 18889 24568
rect 18923 24565 18935 24599
rect 18877 24559 18935 24565
rect 19150 24556 19156 24608
rect 19208 24596 19214 24608
rect 19245 24599 19303 24605
rect 19245 24596 19257 24599
rect 19208 24568 19257 24596
rect 19208 24556 19214 24568
rect 19245 24565 19257 24568
rect 19291 24565 19303 24599
rect 19245 24559 19303 24565
rect 20809 24599 20867 24605
rect 20809 24565 20821 24599
rect 20855 24596 20867 24599
rect 20898 24596 20904 24608
rect 20855 24568 20904 24596
rect 20855 24565 20867 24568
rect 20809 24559 20867 24565
rect 20898 24556 20904 24568
rect 20956 24556 20962 24608
rect 24489 24599 24547 24605
rect 24489 24565 24501 24599
rect 24535 24596 24547 24599
rect 24762 24596 24768 24608
rect 24535 24568 24768 24596
rect 24535 24565 24547 24568
rect 24489 24559 24547 24565
rect 24762 24556 24768 24568
rect 24820 24596 24826 24608
rect 26436 24596 26464 24695
rect 27706 24692 27712 24744
rect 27764 24732 27770 24744
rect 28353 24735 28411 24741
rect 28353 24732 28365 24735
rect 27764 24704 28365 24732
rect 27764 24692 27770 24704
rect 28353 24701 28365 24704
rect 28399 24701 28411 24735
rect 29288 24732 29316 24763
rect 29730 24760 29736 24812
rect 29788 24800 29794 24812
rect 29788 24772 29833 24800
rect 29788 24760 29794 24772
rect 30006 24760 30012 24812
rect 30064 24800 30070 24812
rect 30377 24803 30435 24809
rect 30377 24800 30389 24803
rect 30064 24772 30389 24800
rect 30064 24760 30070 24772
rect 30377 24769 30389 24772
rect 30423 24769 30435 24803
rect 30484 24800 30512 24840
rect 30650 24800 30656 24812
rect 30484 24772 30656 24800
rect 30377 24763 30435 24769
rect 30650 24760 30656 24772
rect 30708 24760 30714 24812
rect 30837 24803 30895 24809
rect 30837 24769 30849 24803
rect 30883 24800 30895 24803
rect 31110 24800 31116 24812
rect 30883 24772 31116 24800
rect 30883 24769 30895 24772
rect 30837 24763 30895 24769
rect 31110 24760 31116 24772
rect 31168 24760 31174 24812
rect 30024 24732 30052 24760
rect 29288 24704 30052 24732
rect 30193 24735 30251 24741
rect 28353 24695 28411 24701
rect 30193 24701 30205 24735
rect 30239 24732 30251 24735
rect 30558 24732 30564 24744
rect 30239 24704 30564 24732
rect 30239 24701 30251 24704
rect 30193 24695 30251 24701
rect 30558 24692 30564 24704
rect 30616 24692 30622 24744
rect 24820 24568 26464 24596
rect 24820 24556 24826 24568
rect 27430 24556 27436 24608
rect 27488 24596 27494 24608
rect 27893 24599 27951 24605
rect 27893 24596 27905 24599
rect 27488 24568 27905 24596
rect 27488 24556 27494 24568
rect 27893 24565 27905 24568
rect 27939 24565 27951 24599
rect 27893 24559 27951 24565
rect 28261 24599 28319 24605
rect 28261 24565 28273 24599
rect 28307 24596 28319 24599
rect 28442 24596 28448 24608
rect 28307 24568 28448 24596
rect 28307 24565 28319 24568
rect 28261 24559 28319 24565
rect 28442 24556 28448 24568
rect 28500 24556 28506 24608
rect 1104 24506 32016 24528
rect 0 24460 800 24474
rect 0 24432 888 24460
rect 1104 24454 2136 24506
rect 2188 24454 12440 24506
rect 12492 24454 22744 24506
rect 22796 24454 32016 24506
rect 32320 24460 33120 24474
rect 1104 24432 32016 24454
rect 32232 24432 33120 24460
rect 0 24418 800 24432
rect 860 24188 888 24432
rect 2317 24395 2375 24401
rect 2317 24361 2329 24395
rect 2363 24392 2375 24395
rect 2682 24392 2688 24404
rect 2363 24364 2688 24392
rect 2363 24361 2375 24364
rect 2317 24355 2375 24361
rect 2682 24352 2688 24364
rect 2740 24352 2746 24404
rect 3786 24392 3792 24404
rect 3747 24364 3792 24392
rect 3786 24352 3792 24364
rect 3844 24352 3850 24404
rect 4890 24352 4896 24404
rect 4948 24392 4954 24404
rect 4985 24395 5043 24401
rect 4985 24392 4997 24395
rect 4948 24364 4997 24392
rect 4948 24352 4954 24364
rect 4985 24361 4997 24364
rect 5031 24361 5043 24395
rect 5350 24392 5356 24404
rect 5311 24364 5356 24392
rect 4985 24355 5043 24361
rect 5350 24352 5356 24364
rect 5408 24352 5414 24404
rect 5534 24352 5540 24404
rect 5592 24392 5598 24404
rect 6457 24395 6515 24401
rect 6457 24392 6469 24395
rect 5592 24364 6469 24392
rect 5592 24352 5598 24364
rect 6457 24361 6469 24364
rect 6503 24361 6515 24395
rect 6457 24355 6515 24361
rect 8113 24395 8171 24401
rect 8113 24361 8125 24395
rect 8159 24392 8171 24395
rect 8754 24392 8760 24404
rect 8159 24364 8760 24392
rect 8159 24361 8171 24364
rect 8113 24355 8171 24361
rect 8754 24352 8760 24364
rect 8812 24352 8818 24404
rect 9125 24395 9183 24401
rect 9125 24361 9137 24395
rect 9171 24392 9183 24395
rect 9398 24392 9404 24404
rect 9171 24364 9404 24392
rect 9171 24361 9183 24364
rect 9125 24355 9183 24361
rect 9398 24352 9404 24364
rect 9456 24352 9462 24404
rect 9582 24352 9588 24404
rect 9640 24392 9646 24404
rect 9677 24395 9735 24401
rect 9677 24392 9689 24395
rect 9640 24364 9689 24392
rect 9640 24352 9646 24364
rect 9677 24361 9689 24364
rect 9723 24361 9735 24395
rect 11422 24392 11428 24404
rect 9677 24355 9735 24361
rect 10428 24364 11428 24392
rect 6362 24284 6368 24336
rect 6420 24324 6426 24336
rect 6641 24327 6699 24333
rect 6641 24324 6653 24327
rect 6420 24296 6653 24324
rect 6420 24284 6426 24296
rect 6641 24293 6653 24296
rect 6687 24293 6699 24327
rect 6641 24287 6699 24293
rect 1670 24216 1676 24268
rect 1728 24256 1734 24268
rect 2409 24259 2467 24265
rect 1728 24228 2360 24256
rect 1728 24216 1734 24228
rect 1765 24191 1823 24197
rect 1765 24188 1777 24191
rect 860 24160 1777 24188
rect 1765 24157 1777 24160
rect 1811 24157 1823 24191
rect 2332 24188 2360 24228
rect 2409 24225 2421 24259
rect 2455 24256 2467 24259
rect 2774 24256 2780 24268
rect 2455 24228 2780 24256
rect 2455 24225 2467 24228
rect 2409 24219 2467 24225
rect 2774 24216 2780 24228
rect 2832 24256 2838 24268
rect 4341 24259 4399 24265
rect 4341 24256 4353 24259
rect 2832 24228 4353 24256
rect 2832 24216 2838 24228
rect 4341 24225 4353 24228
rect 4387 24225 4399 24259
rect 4341 24219 4399 24225
rect 4522 24216 4528 24268
rect 4580 24256 4586 24268
rect 5445 24259 5503 24265
rect 4580 24228 5396 24256
rect 4580 24216 4586 24228
rect 2682 24188 2688 24200
rect 2332 24160 2688 24188
rect 1765 24151 1823 24157
rect 2682 24148 2688 24160
rect 2740 24148 2746 24200
rect 5166 24188 5172 24200
rect 3344 24160 4292 24188
rect 5127 24160 5172 24188
rect 2317 24123 2375 24129
rect 2317 24089 2329 24123
rect 2363 24120 2375 24123
rect 3344 24120 3372 24160
rect 4157 24123 4215 24129
rect 4157 24120 4169 24123
rect 2363 24092 3372 24120
rect 3436 24092 4169 24120
rect 2363 24089 2375 24092
rect 2317 24083 2375 24089
rect 1578 24012 1584 24064
rect 1636 24052 1642 24064
rect 1857 24055 1915 24061
rect 1857 24052 1869 24055
rect 1636 24024 1869 24052
rect 1636 24012 1642 24024
rect 1857 24021 1869 24024
rect 1903 24052 1915 24055
rect 3436 24052 3464 24092
rect 4157 24089 4169 24092
rect 4203 24089 4215 24123
rect 4157 24083 4215 24089
rect 4264 24061 4292 24160
rect 5166 24148 5172 24160
rect 5224 24148 5230 24200
rect 5368 24188 5396 24228
rect 5445 24225 5457 24259
rect 5491 24256 5503 24259
rect 6089 24259 6147 24265
rect 6089 24256 6101 24259
rect 5491 24228 6101 24256
rect 5491 24225 5503 24228
rect 5445 24219 5503 24225
rect 6089 24225 6101 24228
rect 6135 24256 6147 24259
rect 6730 24256 6736 24268
rect 6135 24228 6736 24256
rect 6135 24225 6147 24228
rect 6089 24219 6147 24225
rect 6730 24216 6736 24228
rect 6788 24216 6794 24268
rect 10060 24228 10272 24256
rect 6914 24188 6920 24200
rect 5368 24160 6920 24188
rect 6914 24148 6920 24160
rect 6972 24148 6978 24200
rect 7650 24148 7656 24200
rect 7708 24188 7714 24200
rect 7745 24191 7803 24197
rect 7745 24188 7757 24191
rect 7708 24160 7757 24188
rect 7708 24148 7714 24160
rect 7745 24157 7757 24160
rect 7791 24157 7803 24191
rect 7745 24151 7803 24157
rect 8113 24191 8171 24197
rect 8113 24157 8125 24191
rect 8159 24188 8171 24191
rect 8205 24191 8263 24197
rect 8205 24188 8217 24191
rect 8159 24160 8217 24188
rect 8159 24157 8171 24160
rect 8113 24151 8171 24157
rect 8205 24157 8217 24160
rect 8251 24157 8263 24191
rect 8205 24151 8263 24157
rect 8389 24191 8447 24197
rect 8389 24157 8401 24191
rect 8435 24188 8447 24191
rect 8478 24188 8484 24200
rect 8435 24160 8484 24188
rect 8435 24157 8447 24160
rect 8389 24151 8447 24157
rect 8478 24148 8484 24160
rect 8536 24148 8542 24200
rect 8938 24148 8944 24200
rect 8996 24188 9002 24200
rect 9033 24191 9091 24197
rect 9033 24188 9045 24191
rect 8996 24160 9045 24188
rect 8996 24148 9002 24160
rect 9033 24157 9045 24160
rect 9079 24157 9091 24191
rect 9033 24151 9091 24157
rect 9122 24148 9128 24200
rect 9180 24188 9186 24200
rect 9674 24188 9680 24200
rect 9180 24160 9680 24188
rect 9180 24148 9186 24160
rect 9674 24148 9680 24160
rect 9732 24188 9738 24200
rect 10060 24197 10088 24228
rect 9953 24191 10011 24197
rect 9953 24188 9965 24191
rect 9732 24160 9965 24188
rect 9732 24148 9738 24160
rect 9953 24157 9965 24160
rect 9999 24157 10011 24191
rect 9953 24151 10011 24157
rect 10045 24191 10103 24197
rect 10045 24157 10057 24191
rect 10091 24157 10103 24191
rect 10045 24151 10103 24157
rect 10137 24191 10195 24197
rect 10137 24157 10149 24191
rect 10183 24157 10195 24191
rect 10137 24151 10195 24157
rect 6086 24080 6092 24132
rect 6144 24120 6150 24132
rect 7190 24120 7196 24132
rect 6144 24092 7196 24120
rect 6144 24080 6150 24092
rect 7190 24080 7196 24092
rect 7248 24080 7254 24132
rect 8297 24123 8355 24129
rect 8297 24089 8309 24123
rect 8343 24120 8355 24123
rect 8343 24092 9996 24120
rect 8343 24089 8355 24092
rect 8297 24083 8355 24089
rect 1903 24024 3464 24052
rect 4249 24055 4307 24061
rect 1903 24021 1915 24024
rect 1857 24015 1915 24021
rect 4249 24021 4261 24055
rect 4295 24052 4307 24055
rect 4522 24052 4528 24064
rect 4295 24024 4528 24052
rect 4295 24021 4307 24024
rect 4249 24015 4307 24021
rect 4522 24012 4528 24024
rect 4580 24012 4586 24064
rect 5074 24012 5080 24064
rect 5132 24052 5138 24064
rect 6457 24055 6515 24061
rect 6457 24052 6469 24055
rect 5132 24024 6469 24052
rect 5132 24012 5138 24024
rect 6457 24021 6469 24024
rect 6503 24021 6515 24055
rect 6457 24015 6515 24021
rect 7561 24055 7619 24061
rect 7561 24021 7573 24055
rect 7607 24052 7619 24055
rect 9858 24052 9864 24064
rect 7607 24024 9864 24052
rect 7607 24021 7619 24024
rect 7561 24015 7619 24021
rect 9858 24012 9864 24024
rect 9916 24012 9922 24064
rect 9968 24052 9996 24092
rect 10152 24052 10180 24151
rect 10244 24120 10272 24228
rect 10321 24191 10379 24197
rect 10321 24157 10333 24191
rect 10367 24188 10379 24191
rect 10428 24188 10456 24364
rect 11422 24352 11428 24364
rect 11480 24352 11486 24404
rect 12618 24352 12624 24404
rect 12676 24392 12682 24404
rect 13630 24392 13636 24404
rect 12676 24364 13636 24392
rect 12676 24352 12682 24364
rect 13630 24352 13636 24364
rect 13688 24352 13694 24404
rect 13725 24395 13783 24401
rect 13725 24361 13737 24395
rect 13771 24392 13783 24395
rect 13771 24364 14044 24392
rect 13771 24361 13783 24364
rect 13725 24355 13783 24361
rect 11149 24327 11207 24333
rect 11149 24293 11161 24327
rect 11195 24324 11207 24327
rect 13814 24324 13820 24336
rect 11195 24296 13820 24324
rect 11195 24293 11207 24296
rect 11149 24287 11207 24293
rect 13814 24284 13820 24296
rect 13872 24284 13878 24336
rect 14016 24324 14044 24364
rect 14090 24352 14096 24404
rect 14148 24392 14154 24404
rect 14148 24364 19647 24392
rect 14148 24352 14154 24364
rect 15102 24324 15108 24336
rect 14016 24296 15108 24324
rect 15102 24284 15108 24296
rect 15160 24324 15166 24336
rect 15289 24327 15347 24333
rect 15289 24324 15301 24327
rect 15160 24296 15301 24324
rect 15160 24284 15166 24296
rect 15289 24293 15301 24296
rect 15335 24324 15347 24327
rect 15654 24324 15660 24336
rect 15335 24296 15660 24324
rect 15335 24293 15347 24296
rect 15289 24287 15347 24293
rect 15654 24284 15660 24296
rect 15712 24284 15718 24336
rect 19150 24284 19156 24336
rect 19208 24284 19214 24336
rect 19242 24284 19248 24336
rect 19300 24324 19306 24336
rect 19619 24324 19647 24364
rect 20088 24364 22140 24392
rect 20088 24324 20116 24364
rect 20254 24324 20260 24336
rect 19300 24296 19544 24324
rect 19619 24296 20116 24324
rect 20215 24296 20260 24324
rect 19300 24284 19306 24296
rect 10502 24216 10508 24268
rect 10560 24256 10566 24268
rect 11241 24259 11299 24265
rect 11241 24256 11253 24259
rect 10560 24228 11253 24256
rect 10560 24216 10566 24228
rect 11241 24225 11253 24228
rect 11287 24225 11299 24259
rect 11241 24219 11299 24225
rect 13078 24216 13084 24268
rect 13136 24256 13142 24268
rect 13998 24256 14004 24268
rect 13136 24228 14004 24256
rect 13136 24216 13142 24228
rect 13998 24216 14004 24228
rect 14056 24216 14062 24268
rect 14182 24216 14188 24268
rect 14240 24256 14246 24268
rect 14734 24256 14740 24268
rect 14240 24228 14740 24256
rect 14240 24216 14246 24228
rect 14734 24216 14740 24228
rect 14792 24256 14798 24268
rect 16850 24256 16856 24268
rect 14792 24228 16160 24256
rect 16811 24228 16856 24256
rect 14792 24216 14798 24228
rect 10594 24188 10600 24200
rect 10367 24160 10600 24188
rect 10367 24157 10379 24160
rect 10321 24151 10379 24157
rect 10594 24148 10600 24160
rect 10652 24148 10658 24200
rect 10962 24188 10968 24200
rect 10923 24160 10968 24188
rect 10962 24148 10968 24160
rect 11020 24148 11026 24200
rect 11330 24148 11336 24200
rect 11388 24188 11394 24200
rect 13633 24191 13691 24197
rect 13633 24188 13645 24191
rect 11388 24160 13645 24188
rect 11388 24148 11394 24160
rect 13633 24157 13645 24160
rect 13679 24157 13691 24191
rect 13633 24151 13691 24157
rect 13722 24148 13728 24200
rect 13780 24188 13786 24200
rect 14093 24191 14151 24197
rect 14093 24188 14105 24191
rect 13780 24160 14105 24188
rect 13780 24148 13786 24160
rect 14093 24157 14105 24160
rect 14139 24157 14151 24191
rect 14093 24151 14151 24157
rect 14277 24191 14335 24197
rect 14277 24157 14289 24191
rect 14323 24188 14335 24191
rect 14918 24188 14924 24200
rect 14323 24160 14924 24188
rect 14323 24157 14335 24160
rect 14277 24151 14335 24157
rect 14918 24148 14924 24160
rect 14976 24148 14982 24200
rect 15102 24188 15108 24200
rect 15063 24160 15108 24188
rect 15102 24148 15108 24160
rect 15160 24148 15166 24200
rect 15381 24191 15439 24197
rect 15381 24157 15393 24191
rect 15427 24188 15439 24191
rect 15838 24188 15844 24200
rect 15427 24160 15844 24188
rect 15427 24157 15439 24160
rect 15381 24151 15439 24157
rect 15838 24148 15844 24160
rect 15896 24148 15902 24200
rect 15930 24148 15936 24200
rect 15988 24188 15994 24200
rect 16025 24191 16083 24197
rect 16025 24188 16037 24191
rect 15988 24160 16037 24188
rect 15988 24148 15994 24160
rect 16025 24157 16037 24160
rect 16071 24157 16083 24191
rect 16132 24188 16160 24228
rect 16850 24216 16856 24228
rect 16908 24216 16914 24268
rect 19168 24256 19196 24284
rect 19516 24256 19544 24296
rect 20254 24284 20260 24296
rect 20312 24284 20318 24336
rect 19613 24259 19671 24265
rect 19613 24256 19625 24259
rect 19168 24228 19472 24256
rect 19516 24228 19625 24256
rect 19444 24197 19472 24228
rect 19613 24225 19625 24228
rect 19659 24225 19671 24259
rect 20806 24256 20812 24268
rect 20767 24228 20812 24256
rect 19613 24219 19671 24225
rect 20806 24216 20812 24228
rect 20864 24216 20870 24268
rect 22112 24256 22140 24364
rect 22186 24352 22192 24404
rect 22244 24392 22250 24404
rect 25866 24392 25872 24404
rect 22244 24364 22289 24392
rect 25827 24364 25872 24392
rect 22244 24352 22250 24364
rect 25866 24352 25872 24364
rect 25924 24352 25930 24404
rect 28169 24395 28227 24401
rect 28169 24361 28181 24395
rect 28215 24392 28227 24395
rect 29178 24392 29184 24404
rect 28215 24364 29184 24392
rect 28215 24361 28227 24364
rect 28169 24355 28227 24361
rect 29178 24352 29184 24364
rect 29236 24352 29242 24404
rect 22646 24284 22652 24336
rect 22704 24324 22710 24336
rect 22704 24296 22749 24324
rect 22704 24284 22710 24296
rect 27614 24284 27620 24336
rect 27672 24324 27678 24336
rect 27709 24327 27767 24333
rect 27709 24324 27721 24327
rect 27672 24296 27721 24324
rect 27672 24284 27678 24296
rect 27709 24293 27721 24296
rect 27755 24324 27767 24327
rect 28534 24324 28540 24336
rect 27755 24296 28540 24324
rect 27755 24293 27767 24296
rect 27709 24287 27767 24293
rect 28534 24284 28540 24296
rect 28592 24284 28598 24336
rect 32232 24324 32260 24432
rect 32320 24418 33120 24432
rect 32232 24296 32352 24324
rect 23290 24256 23296 24268
rect 22112 24228 23060 24256
rect 23251 24228 23296 24256
rect 19429 24191 19487 24197
rect 16132 24160 17632 24188
rect 16025 24151 16083 24157
rect 11422 24120 11428 24132
rect 10244 24092 11428 24120
rect 11422 24080 11428 24092
rect 11480 24080 11486 24132
rect 11790 24120 11796 24132
rect 11751 24092 11796 24120
rect 11790 24080 11796 24092
rect 11848 24080 11854 24132
rect 12158 24080 12164 24132
rect 12216 24120 12222 24132
rect 14461 24123 14519 24129
rect 14461 24120 14473 24123
rect 12216 24092 14473 24120
rect 12216 24080 12222 24092
rect 14461 24089 14473 24092
rect 14507 24089 14519 24123
rect 17120 24123 17178 24129
rect 14461 24083 14519 24089
rect 14568 24092 16344 24120
rect 10778 24052 10784 24064
rect 9968 24024 10180 24052
rect 10739 24024 10784 24052
rect 10778 24012 10784 24024
rect 10836 24012 10842 24064
rect 12802 24012 12808 24064
rect 12860 24052 12866 24064
rect 13081 24055 13139 24061
rect 13081 24052 13093 24055
rect 12860 24024 13093 24052
rect 12860 24012 12866 24024
rect 13081 24021 13093 24024
rect 13127 24021 13139 24055
rect 13081 24015 13139 24021
rect 13998 24012 14004 24064
rect 14056 24052 14062 24064
rect 14568 24052 14596 24092
rect 14918 24052 14924 24064
rect 14056 24024 14596 24052
rect 14879 24024 14924 24052
rect 14056 24012 14062 24024
rect 14918 24012 14924 24024
rect 14976 24012 14982 24064
rect 16206 24052 16212 24064
rect 16167 24024 16212 24052
rect 16206 24012 16212 24024
rect 16264 24012 16270 24064
rect 16316 24052 16344 24092
rect 17120 24089 17132 24123
rect 17166 24120 17178 24123
rect 17494 24120 17500 24132
rect 17166 24092 17500 24120
rect 17166 24089 17178 24092
rect 17120 24083 17178 24089
rect 17494 24080 17500 24092
rect 17552 24080 17558 24132
rect 17604 24120 17632 24160
rect 19429 24157 19441 24191
rect 19475 24157 19487 24191
rect 19429 24151 19487 24157
rect 19705 24191 19763 24197
rect 19705 24157 19717 24191
rect 19751 24188 19763 24191
rect 20070 24188 20076 24200
rect 19751 24160 20076 24188
rect 19751 24157 19763 24160
rect 19705 24151 19763 24157
rect 20070 24148 20076 24160
rect 20128 24148 20134 24200
rect 20165 24191 20223 24197
rect 20165 24157 20177 24191
rect 20211 24157 20223 24191
rect 20165 24151 20223 24157
rect 20180 24120 20208 24151
rect 20898 24148 20904 24200
rect 20956 24188 20962 24200
rect 21065 24191 21123 24197
rect 21065 24188 21077 24191
rect 20956 24160 21077 24188
rect 20956 24148 20962 24160
rect 21065 24157 21077 24160
rect 21111 24157 21123 24191
rect 21065 24151 21123 24157
rect 22646 24148 22652 24200
rect 22704 24188 22710 24200
rect 22830 24188 22836 24200
rect 22704 24160 22836 24188
rect 22704 24148 22710 24160
rect 22830 24148 22836 24160
rect 22888 24148 22894 24200
rect 23032 24197 23060 24228
rect 23290 24216 23296 24228
rect 23348 24216 23354 24268
rect 27338 24216 27344 24268
rect 27396 24256 27402 24268
rect 27396 24228 28396 24256
rect 27396 24216 27402 24228
rect 23017 24191 23075 24197
rect 23017 24157 23029 24191
rect 23063 24188 23075 24191
rect 23198 24188 23204 24200
rect 23063 24160 23204 24188
rect 23063 24157 23075 24160
rect 23017 24151 23075 24157
rect 23198 24148 23204 24160
rect 23256 24148 23262 24200
rect 24210 24148 24216 24200
rect 24268 24188 24274 24200
rect 28368 24197 28396 24228
rect 24489 24191 24547 24197
rect 24489 24188 24501 24191
rect 24268 24160 24501 24188
rect 24268 24148 24274 24160
rect 24489 24157 24501 24160
rect 24535 24157 24547 24191
rect 24489 24151 24547 24157
rect 24756 24191 24814 24197
rect 24756 24157 24768 24191
rect 24802 24157 24814 24191
rect 24756 24151 24814 24157
rect 26329 24191 26387 24197
rect 26329 24157 26341 24191
rect 26375 24157 26387 24191
rect 26329 24151 26387 24157
rect 28353 24191 28411 24197
rect 28353 24157 28365 24191
rect 28399 24157 28411 24191
rect 28353 24151 28411 24157
rect 28629 24191 28687 24197
rect 28629 24157 28641 24191
rect 28675 24157 28687 24191
rect 28629 24151 28687 24157
rect 17604 24092 19472 24120
rect 17954 24052 17960 24064
rect 16316 24024 17960 24052
rect 17954 24012 17960 24024
rect 18012 24012 18018 24064
rect 18233 24055 18291 24061
rect 18233 24021 18245 24055
rect 18279 24052 18291 24055
rect 18322 24052 18328 24064
rect 18279 24024 18328 24052
rect 18279 24021 18291 24024
rect 18233 24015 18291 24021
rect 18322 24012 18328 24024
rect 18380 24012 18386 24064
rect 19245 24055 19303 24061
rect 19245 24021 19257 24055
rect 19291 24052 19303 24055
rect 19334 24052 19340 24064
rect 19291 24024 19340 24052
rect 19291 24021 19303 24024
rect 19245 24015 19303 24021
rect 19334 24012 19340 24024
rect 19392 24012 19398 24064
rect 19444 24052 19472 24092
rect 19619 24092 20208 24120
rect 19619 24052 19647 24092
rect 20254 24080 20260 24132
rect 20312 24120 20318 24132
rect 21542 24120 21548 24132
rect 20312 24092 21548 24120
rect 20312 24080 20318 24092
rect 21542 24080 21548 24092
rect 21600 24080 21606 24132
rect 23106 24052 23112 24064
rect 19444 24024 19647 24052
rect 23067 24024 23112 24052
rect 23106 24012 23112 24024
rect 23164 24012 23170 24064
rect 24504 24052 24532 24151
rect 24670 24080 24676 24132
rect 24728 24120 24734 24132
rect 24780 24120 24808 24151
rect 24728 24092 24808 24120
rect 24728 24080 24734 24092
rect 26344 24052 26372 24151
rect 26596 24123 26654 24129
rect 26596 24089 26608 24123
rect 26642 24120 26654 24123
rect 27430 24120 27436 24132
rect 26642 24092 27436 24120
rect 26642 24089 26654 24092
rect 26596 24083 26654 24089
rect 27430 24080 27436 24092
rect 27488 24080 27494 24132
rect 27522 24080 27528 24132
rect 27580 24120 27586 24132
rect 28644 24120 28672 24151
rect 28718 24148 28724 24200
rect 28776 24188 28782 24200
rect 28813 24191 28871 24197
rect 28813 24188 28825 24191
rect 28776 24160 28825 24188
rect 28776 24148 28782 24160
rect 28813 24157 28825 24160
rect 28859 24188 28871 24191
rect 28994 24188 29000 24200
rect 28859 24160 29000 24188
rect 28859 24157 28871 24160
rect 28813 24151 28871 24157
rect 28994 24148 29000 24160
rect 29052 24148 29058 24200
rect 30006 24148 30012 24200
rect 30064 24188 30070 24200
rect 30285 24191 30343 24197
rect 30285 24188 30297 24191
rect 30064 24160 30297 24188
rect 30064 24148 30070 24160
rect 30285 24157 30297 24160
rect 30331 24157 30343 24191
rect 30285 24151 30343 24157
rect 30374 24148 30380 24200
rect 30432 24188 30438 24200
rect 30561 24191 30619 24197
rect 30561 24188 30573 24191
rect 30432 24160 30573 24188
rect 30432 24148 30438 24160
rect 30561 24157 30573 24160
rect 30607 24188 30619 24191
rect 30650 24188 30656 24200
rect 30607 24160 30656 24188
rect 30607 24157 30619 24160
rect 30561 24151 30619 24157
rect 30650 24148 30656 24160
rect 30708 24148 30714 24200
rect 30745 24191 30803 24197
rect 30745 24157 30757 24191
rect 30791 24188 30803 24191
rect 31202 24188 31208 24200
rect 30791 24160 31208 24188
rect 30791 24157 30803 24160
rect 30745 24151 30803 24157
rect 27580 24092 28672 24120
rect 27580 24080 27586 24092
rect 30466 24080 30472 24132
rect 30524 24120 30530 24132
rect 30760 24120 30788 24151
rect 31202 24148 31208 24160
rect 31260 24148 31266 24200
rect 30524 24092 30788 24120
rect 30524 24080 30530 24092
rect 27798 24052 27804 24064
rect 24504 24024 27804 24052
rect 27798 24012 27804 24024
rect 27856 24012 27862 24064
rect 30101 24055 30159 24061
rect 30101 24021 30113 24055
rect 30147 24052 30159 24055
rect 30834 24052 30840 24064
rect 30147 24024 30840 24052
rect 30147 24021 30159 24024
rect 30101 24015 30159 24021
rect 30834 24012 30840 24024
rect 30892 24012 30898 24064
rect 1104 23962 32016 23984
rect 1104 23910 7288 23962
rect 7340 23910 17592 23962
rect 17644 23910 27896 23962
rect 27948 23910 32016 23962
rect 1104 23888 32016 23910
rect 1302 23808 1308 23860
rect 1360 23848 1366 23860
rect 1486 23848 1492 23860
rect 1360 23820 1492 23848
rect 1360 23808 1366 23820
rect 1486 23808 1492 23820
rect 1544 23808 1550 23860
rect 2774 23808 2780 23860
rect 2832 23848 2838 23860
rect 5534 23848 5540 23860
rect 2832 23820 2877 23848
rect 3988 23820 5540 23848
rect 2832 23808 2838 23820
rect 3605 23783 3663 23789
rect 3605 23749 3617 23783
rect 3651 23780 3663 23783
rect 3694 23780 3700 23792
rect 3651 23752 3700 23780
rect 3651 23749 3663 23752
rect 3605 23743 3663 23749
rect 3694 23740 3700 23752
rect 3752 23740 3758 23792
rect 1394 23712 1400 23724
rect 1355 23684 1400 23712
rect 1394 23672 1400 23684
rect 1452 23672 1458 23724
rect 1486 23672 1492 23724
rect 1544 23712 1550 23724
rect 1653 23715 1711 23721
rect 1653 23712 1665 23715
rect 1544 23684 1665 23712
rect 1544 23672 1550 23684
rect 1653 23681 1665 23684
rect 1699 23681 1711 23715
rect 1653 23675 1711 23681
rect 2222 23672 2228 23724
rect 2280 23712 2286 23724
rect 3988 23712 4016 23820
rect 5534 23808 5540 23820
rect 5592 23808 5598 23860
rect 5718 23808 5724 23860
rect 5776 23808 5782 23860
rect 6365 23851 6423 23857
rect 6365 23817 6377 23851
rect 6411 23848 6423 23851
rect 6638 23848 6644 23860
rect 6411 23820 6644 23848
rect 6411 23817 6423 23820
rect 6365 23811 6423 23817
rect 6638 23808 6644 23820
rect 6696 23808 6702 23860
rect 6733 23851 6791 23857
rect 6733 23817 6745 23851
rect 6779 23848 6791 23851
rect 6914 23848 6920 23860
rect 6779 23820 6920 23848
rect 6779 23817 6791 23820
rect 6733 23811 6791 23817
rect 6914 23808 6920 23820
rect 6972 23808 6978 23860
rect 8938 23848 8944 23860
rect 8851 23820 8944 23848
rect 8938 23808 8944 23820
rect 8996 23848 9002 23860
rect 9582 23848 9588 23860
rect 8996 23820 9588 23848
rect 8996 23808 9002 23820
rect 9582 23808 9588 23820
rect 9640 23848 9646 23860
rect 10594 23848 10600 23860
rect 9640 23820 10600 23848
rect 9640 23808 9646 23820
rect 10594 23808 10600 23820
rect 10652 23808 10658 23860
rect 11054 23808 11060 23860
rect 11112 23848 11118 23860
rect 11793 23851 11851 23857
rect 11793 23848 11805 23851
rect 11112 23820 11805 23848
rect 11112 23808 11118 23820
rect 11793 23817 11805 23820
rect 11839 23817 11851 23851
rect 12158 23848 12164 23860
rect 12119 23820 12164 23848
rect 11793 23811 11851 23817
rect 12158 23808 12164 23820
rect 12216 23808 12222 23860
rect 12253 23851 12311 23857
rect 12253 23817 12265 23851
rect 12299 23848 12311 23851
rect 13173 23851 13231 23857
rect 13173 23848 13185 23851
rect 12299 23820 13185 23848
rect 12299 23817 12311 23820
rect 12253 23811 12311 23817
rect 13173 23817 13185 23820
rect 13219 23817 13231 23851
rect 13173 23811 13231 23817
rect 13541 23851 13599 23857
rect 13541 23817 13553 23851
rect 13587 23848 13599 23851
rect 15378 23848 15384 23860
rect 13587 23820 15384 23848
rect 13587 23817 13599 23820
rect 13541 23811 13599 23817
rect 15378 23808 15384 23820
rect 15436 23848 15442 23860
rect 16758 23848 16764 23860
rect 15436 23820 16764 23848
rect 15436 23808 15442 23820
rect 16758 23808 16764 23820
rect 16816 23808 16822 23860
rect 17129 23851 17187 23857
rect 17129 23817 17141 23851
rect 17175 23848 17187 23851
rect 19518 23848 19524 23860
rect 17175 23820 19524 23848
rect 17175 23817 17187 23820
rect 17129 23811 17187 23817
rect 19518 23808 19524 23820
rect 19576 23808 19582 23860
rect 28350 23848 28356 23860
rect 19996 23820 28356 23848
rect 4062 23740 4068 23792
rect 4120 23780 4126 23792
rect 5736 23780 5764 23808
rect 7828 23783 7886 23789
rect 4120 23752 4936 23780
rect 5736 23752 7788 23780
rect 4120 23740 4126 23752
rect 4908 23721 4936 23752
rect 2280 23684 4016 23712
rect 4433 23715 4491 23721
rect 2280 23672 2286 23684
rect 4433 23681 4445 23715
rect 4479 23681 4491 23715
rect 4433 23675 4491 23681
rect 4709 23715 4767 23721
rect 4709 23681 4721 23715
rect 4755 23712 4767 23715
rect 4893 23715 4951 23721
rect 4755 23684 4844 23712
rect 4755 23681 4767 23684
rect 4709 23675 4767 23681
rect 4448 23644 4476 23675
rect 4816 23644 4844 23684
rect 4893 23681 4905 23715
rect 4939 23681 4951 23715
rect 4893 23675 4951 23681
rect 5445 23715 5503 23721
rect 5445 23681 5457 23715
rect 5491 23712 5503 23715
rect 5718 23712 5724 23724
rect 5491 23684 5724 23712
rect 5491 23681 5503 23684
rect 5445 23675 5503 23681
rect 5718 23672 5724 23684
rect 5776 23672 5782 23724
rect 6178 23672 6184 23724
rect 6236 23712 6242 23724
rect 6362 23712 6368 23724
rect 6236 23684 6368 23712
rect 6236 23672 6242 23684
rect 6362 23672 6368 23684
rect 6420 23672 6426 23724
rect 7561 23715 7619 23721
rect 7561 23681 7573 23715
rect 7607 23681 7619 23715
rect 7760 23712 7788 23752
rect 7828 23749 7840 23783
rect 7874 23780 7886 23783
rect 8294 23780 8300 23792
rect 7874 23752 8300 23780
rect 7874 23749 7886 23752
rect 7828 23743 7886 23749
rect 8294 23740 8300 23752
rect 8352 23740 8358 23792
rect 9674 23740 9680 23792
rect 9732 23780 9738 23792
rect 9732 23752 10456 23780
rect 9732 23740 9738 23752
rect 7760 23684 9720 23712
rect 7561 23675 7619 23681
rect 4982 23644 4988 23656
rect 4448 23616 4752 23644
rect 4816 23616 4988 23644
rect 4724 23588 4752 23616
rect 4982 23604 4988 23616
rect 5040 23644 5046 23656
rect 5258 23644 5264 23656
rect 5040 23616 5264 23644
rect 5040 23604 5046 23616
rect 5258 23604 5264 23616
rect 5316 23604 5322 23656
rect 6546 23644 6552 23656
rect 5460 23616 6552 23644
rect 5460 23588 5488 23616
rect 6546 23604 6552 23616
rect 6604 23644 6610 23656
rect 6825 23647 6883 23653
rect 6825 23644 6837 23647
rect 6604 23616 6837 23644
rect 6604 23604 6610 23616
rect 6825 23613 6837 23616
rect 6871 23613 6883 23647
rect 6825 23607 6883 23613
rect 6917 23647 6975 23653
rect 6917 23613 6929 23647
rect 6963 23613 6975 23647
rect 6917 23607 6975 23613
rect 2958 23536 2964 23588
rect 3016 23576 3022 23588
rect 3237 23579 3295 23585
rect 3237 23576 3249 23579
rect 3016 23548 3249 23576
rect 3016 23536 3022 23548
rect 3237 23545 3249 23548
rect 3283 23545 3295 23579
rect 3237 23539 3295 23545
rect 4706 23536 4712 23588
rect 4764 23536 4770 23588
rect 5442 23536 5448 23588
rect 5500 23536 5506 23588
rect 6638 23536 6644 23588
rect 6696 23576 6702 23588
rect 6932 23576 6960 23607
rect 6696 23548 6960 23576
rect 6696 23536 6702 23548
rect 2682 23468 2688 23520
rect 2740 23508 2746 23520
rect 3605 23511 3663 23517
rect 3605 23508 3617 23511
rect 2740 23480 3617 23508
rect 2740 23468 2746 23480
rect 3605 23477 3617 23480
rect 3651 23477 3663 23511
rect 3786 23508 3792 23520
rect 3747 23480 3792 23508
rect 3605 23471 3663 23477
rect 3786 23468 3792 23480
rect 3844 23468 3850 23520
rect 4154 23468 4160 23520
rect 4212 23508 4218 23520
rect 4249 23511 4307 23517
rect 4249 23508 4261 23511
rect 4212 23480 4261 23508
rect 4212 23468 4218 23480
rect 4249 23477 4261 23480
rect 4295 23477 4307 23511
rect 4249 23471 4307 23477
rect 4798 23468 4804 23520
rect 4856 23508 4862 23520
rect 5166 23508 5172 23520
rect 4856 23480 5172 23508
rect 4856 23468 4862 23480
rect 5166 23468 5172 23480
rect 5224 23508 5230 23520
rect 5537 23511 5595 23517
rect 5537 23508 5549 23511
rect 5224 23480 5549 23508
rect 5224 23468 5230 23480
rect 5537 23477 5549 23480
rect 5583 23477 5595 23511
rect 5537 23471 5595 23477
rect 6822 23468 6828 23520
rect 6880 23508 6886 23520
rect 7576 23508 7604 23675
rect 9692 23644 9720 23684
rect 9858 23672 9864 23724
rect 9916 23712 9922 23724
rect 10045 23715 10103 23721
rect 10045 23712 10057 23715
rect 9916 23684 10057 23712
rect 9916 23672 9922 23684
rect 10045 23681 10057 23684
rect 10091 23681 10103 23715
rect 10318 23712 10324 23724
rect 10279 23684 10324 23712
rect 10045 23675 10103 23681
rect 10318 23672 10324 23684
rect 10376 23672 10382 23724
rect 10428 23712 10456 23752
rect 11422 23740 11428 23792
rect 11480 23780 11486 23792
rect 13998 23780 14004 23792
rect 11480 23752 14004 23780
rect 11480 23740 11486 23752
rect 13998 23740 14004 23752
rect 14056 23740 14062 23792
rect 14636 23783 14694 23789
rect 14636 23749 14648 23783
rect 14682 23780 14694 23783
rect 14918 23780 14924 23792
rect 14682 23752 14924 23780
rect 14682 23749 14694 23752
rect 14636 23743 14694 23749
rect 14918 23740 14924 23752
rect 14976 23740 14982 23792
rect 15746 23740 15752 23792
rect 15804 23780 15810 23792
rect 17037 23783 17095 23789
rect 17037 23780 17049 23783
rect 15804 23752 17049 23780
rect 15804 23740 15810 23752
rect 17037 23749 17049 23752
rect 17083 23780 17095 23783
rect 17083 23752 17356 23780
rect 17083 23749 17095 23752
rect 17037 23743 17095 23749
rect 10502 23712 10508 23724
rect 10428 23684 10508 23712
rect 10502 23672 10508 23684
rect 10560 23712 10566 23724
rect 13633 23715 13691 23721
rect 10560 23684 10653 23712
rect 10560 23672 10566 23684
rect 13633 23681 13645 23715
rect 13679 23712 13691 23715
rect 13679 23684 14136 23712
rect 13679 23681 13691 23684
rect 13633 23675 13691 23681
rect 12345 23647 12403 23653
rect 9692 23616 9996 23644
rect 9968 23576 9996 23616
rect 12345 23613 12357 23647
rect 12391 23644 12403 23647
rect 12526 23644 12532 23656
rect 12391 23616 12532 23644
rect 12391 23613 12403 23616
rect 12345 23607 12403 23613
rect 12526 23604 12532 23616
rect 12584 23604 12590 23656
rect 12894 23604 12900 23656
rect 12952 23644 12958 23656
rect 13725 23647 13783 23653
rect 13725 23644 13737 23647
rect 12952 23616 13737 23644
rect 12952 23604 12958 23616
rect 13725 23613 13737 23616
rect 13771 23613 13783 23647
rect 14108 23644 14136 23684
rect 15838 23672 15844 23724
rect 15896 23712 15902 23724
rect 17328 23712 17356 23752
rect 17862 23740 17868 23792
rect 17920 23780 17926 23792
rect 19886 23780 19892 23792
rect 17920 23752 19892 23780
rect 17920 23740 17926 23752
rect 19886 23740 19892 23752
rect 19944 23740 19950 23792
rect 19996 23789 20024 23820
rect 28350 23808 28356 23820
rect 28408 23808 28414 23860
rect 30282 23808 30288 23860
rect 30340 23848 30346 23860
rect 30653 23851 30711 23857
rect 30653 23848 30665 23851
rect 30340 23820 30665 23848
rect 30340 23808 30346 23820
rect 30653 23817 30665 23820
rect 30699 23817 30711 23851
rect 30653 23811 30711 23817
rect 19981 23783 20039 23789
rect 19981 23749 19993 23783
rect 20027 23749 20039 23783
rect 20714 23780 20720 23792
rect 19981 23743 20039 23749
rect 20456 23752 20720 23780
rect 18049 23715 18107 23721
rect 18049 23712 18061 23715
rect 15896 23684 17264 23712
rect 17328 23684 18061 23712
rect 15896 23672 15902 23684
rect 14274 23644 14280 23656
rect 14108 23616 14280 23644
rect 13725 23607 13783 23613
rect 14274 23604 14280 23616
rect 14332 23604 14338 23656
rect 17236 23653 17264 23684
rect 18049 23681 18061 23684
rect 18095 23681 18107 23715
rect 18049 23675 18107 23681
rect 18233 23715 18291 23721
rect 18233 23681 18245 23715
rect 18279 23702 18291 23715
rect 18340 23702 18552 23718
rect 18279 23690 18552 23702
rect 18279 23681 18368 23690
rect 18233 23675 18368 23681
rect 18239 23674 18368 23675
rect 14369 23647 14427 23653
rect 14369 23613 14381 23647
rect 14415 23613 14427 23647
rect 14369 23607 14427 23613
rect 17221 23647 17279 23653
rect 17221 23613 17233 23647
rect 17267 23613 17279 23647
rect 18524 23644 18552 23690
rect 18598 23672 18604 23724
rect 18656 23712 18662 23724
rect 20254 23712 20260 23724
rect 18656 23684 20260 23712
rect 18656 23672 18662 23684
rect 20254 23672 20260 23684
rect 20312 23672 20318 23724
rect 20456 23644 20484 23752
rect 20714 23740 20720 23752
rect 20772 23740 20778 23792
rect 21266 23740 21272 23792
rect 21324 23780 21330 23792
rect 21821 23783 21879 23789
rect 21821 23780 21833 23783
rect 21324 23752 21833 23780
rect 21324 23740 21330 23752
rect 21821 23749 21833 23752
rect 21867 23749 21879 23783
rect 21821 23743 21879 23749
rect 21910 23740 21916 23792
rect 21968 23780 21974 23792
rect 22021 23783 22079 23789
rect 22021 23780 22033 23783
rect 21968 23752 22033 23780
rect 21968 23740 21974 23752
rect 22021 23749 22033 23752
rect 22067 23749 22079 23783
rect 32324 23780 32352 24296
rect 22021 23743 22079 23749
rect 22112 23752 32352 23780
rect 20622 23712 20628 23724
rect 20583 23684 20628 23712
rect 20622 23672 20628 23684
rect 20680 23672 20686 23724
rect 22112 23712 22140 23752
rect 20732 23684 22140 23712
rect 23100 23715 23158 23721
rect 18524 23616 20484 23644
rect 17221 23607 17279 23613
rect 9968 23548 10364 23576
rect 6880 23480 7604 23508
rect 9861 23511 9919 23517
rect 6880 23468 6886 23480
rect 9861 23477 9873 23511
rect 9907 23508 9919 23511
rect 10226 23508 10232 23520
rect 9907 23480 10232 23508
rect 9907 23477 9919 23480
rect 9861 23471 9919 23477
rect 10226 23468 10232 23480
rect 10284 23468 10290 23520
rect 10336 23508 10364 23548
rect 12802 23536 12808 23588
rect 12860 23576 12866 23588
rect 14384 23576 14412 23607
rect 20732 23576 20760 23684
rect 23100 23681 23112 23715
rect 23146 23712 23158 23715
rect 23658 23712 23664 23724
rect 23146 23684 23664 23712
rect 23146 23681 23158 23684
rect 23100 23675 23158 23681
rect 23658 23672 23664 23684
rect 23716 23672 23722 23724
rect 25222 23712 25228 23724
rect 25135 23684 25228 23712
rect 25222 23672 25228 23684
rect 25280 23712 25286 23724
rect 25498 23712 25504 23724
rect 25280 23684 25360 23712
rect 25411 23684 25504 23712
rect 25280 23672 25286 23684
rect 20901 23647 20959 23653
rect 20901 23613 20913 23647
rect 20947 23644 20959 23647
rect 22462 23644 22468 23656
rect 20947 23616 22468 23644
rect 20947 23613 20959 23616
rect 20901 23607 20959 23613
rect 22462 23604 22468 23616
rect 22520 23604 22526 23656
rect 22830 23644 22836 23656
rect 22791 23616 22836 23644
rect 22830 23604 22836 23616
rect 22888 23604 22894 23656
rect 22094 23576 22100 23588
rect 12860 23548 14412 23576
rect 15580 23548 20760 23576
rect 20824 23548 22100 23576
rect 12860 23536 12866 23548
rect 15580 23508 15608 23548
rect 15746 23508 15752 23520
rect 10336 23480 15608 23508
rect 15707 23480 15752 23508
rect 15746 23468 15752 23480
rect 15804 23468 15810 23520
rect 15838 23468 15844 23520
rect 15896 23508 15902 23520
rect 16669 23511 16727 23517
rect 16669 23508 16681 23511
rect 15896 23480 16681 23508
rect 15896 23468 15902 23480
rect 16669 23477 16681 23480
rect 16715 23477 16727 23511
rect 16669 23471 16727 23477
rect 16942 23468 16948 23520
rect 17000 23508 17006 23520
rect 17402 23508 17408 23520
rect 17000 23480 17408 23508
rect 17000 23468 17006 23480
rect 17402 23468 17408 23480
rect 17460 23468 17466 23520
rect 18049 23511 18107 23517
rect 18049 23477 18061 23511
rect 18095 23508 18107 23511
rect 18598 23508 18604 23520
rect 18095 23480 18604 23508
rect 18095 23477 18107 23480
rect 18049 23471 18107 23477
rect 18598 23468 18604 23480
rect 18656 23468 18662 23520
rect 20438 23508 20444 23520
rect 20399 23480 20444 23508
rect 20438 23468 20444 23480
rect 20496 23468 20502 23520
rect 20824 23517 20852 23548
rect 22094 23536 22100 23548
rect 22152 23536 22158 23588
rect 24118 23536 24124 23588
rect 24176 23576 24182 23588
rect 24213 23579 24271 23585
rect 24213 23576 24225 23579
rect 24176 23548 24225 23576
rect 24176 23536 24182 23548
rect 24213 23545 24225 23548
rect 24259 23545 24271 23579
rect 25130 23576 25136 23588
rect 24213 23539 24271 23545
rect 24688 23548 25136 23576
rect 20809 23511 20867 23517
rect 20809 23477 20821 23511
rect 20855 23477 20867 23511
rect 22002 23508 22008 23520
rect 21963 23480 22008 23508
rect 20809 23471 20867 23477
rect 22002 23468 22008 23480
rect 22060 23468 22066 23520
rect 22189 23511 22247 23517
rect 22189 23477 22201 23511
rect 22235 23508 22247 23511
rect 24688 23508 24716 23548
rect 25130 23536 25136 23548
rect 25188 23536 25194 23588
rect 25332 23576 25360 23684
rect 25498 23672 25504 23684
rect 25556 23672 25562 23724
rect 25590 23672 25596 23724
rect 25648 23712 25654 23724
rect 25685 23715 25743 23721
rect 25685 23712 25697 23715
rect 25648 23684 25697 23712
rect 25648 23672 25654 23684
rect 25685 23681 25697 23684
rect 25731 23681 25743 23715
rect 26234 23712 26240 23724
rect 26195 23684 26240 23712
rect 25685 23675 25743 23681
rect 26234 23672 26240 23684
rect 26292 23672 26298 23724
rect 27154 23712 27160 23724
rect 27115 23684 27160 23712
rect 27154 23672 27160 23684
rect 27212 23672 27218 23724
rect 27430 23712 27436 23724
rect 27391 23684 27436 23712
rect 27430 23672 27436 23684
rect 27488 23672 27494 23724
rect 27614 23712 27620 23724
rect 27575 23684 27620 23712
rect 27614 23672 27620 23684
rect 27672 23672 27678 23724
rect 28077 23715 28135 23721
rect 28077 23681 28089 23715
rect 28123 23712 28135 23715
rect 28258 23712 28264 23724
rect 28123 23684 28264 23712
rect 28123 23681 28135 23684
rect 28077 23675 28135 23681
rect 28258 23672 28264 23684
rect 28316 23712 28322 23724
rect 28902 23712 28908 23724
rect 28316 23684 28908 23712
rect 28316 23672 28322 23684
rect 28902 23672 28908 23684
rect 28960 23712 28966 23724
rect 29365 23715 29423 23721
rect 29365 23712 29377 23715
rect 28960 23684 29377 23712
rect 28960 23672 28966 23684
rect 29365 23681 29377 23684
rect 29411 23681 29423 23715
rect 30834 23712 30840 23724
rect 30795 23684 30840 23712
rect 29365 23675 29423 23681
rect 30834 23672 30840 23684
rect 30892 23672 30898 23724
rect 30926 23672 30932 23724
rect 30984 23712 30990 23724
rect 31021 23715 31079 23721
rect 31021 23712 31033 23715
rect 30984 23684 31033 23712
rect 30984 23672 30990 23684
rect 31021 23681 31033 23684
rect 31067 23681 31079 23715
rect 31021 23675 31079 23681
rect 25516 23644 25544 23672
rect 26418 23644 26424 23656
rect 25516 23616 26424 23644
rect 26418 23604 26424 23616
rect 26476 23604 26482 23656
rect 26973 23647 27031 23653
rect 26973 23613 26985 23647
rect 27019 23644 27031 23647
rect 28166 23644 28172 23656
rect 27019 23616 28172 23644
rect 27019 23613 27031 23616
rect 26973 23607 27031 23613
rect 28166 23604 28172 23616
rect 28224 23604 28230 23656
rect 28353 23647 28411 23653
rect 28353 23613 28365 23647
rect 28399 23613 28411 23647
rect 28353 23607 28411 23613
rect 29641 23647 29699 23653
rect 29641 23613 29653 23647
rect 29687 23644 29699 23647
rect 30374 23644 30380 23656
rect 29687 23616 30380 23644
rect 29687 23613 29699 23616
rect 29641 23607 29699 23613
rect 25866 23576 25872 23588
rect 25332 23548 25872 23576
rect 25866 23536 25872 23548
rect 25924 23536 25930 23588
rect 27430 23536 27436 23588
rect 27488 23576 27494 23588
rect 28368 23576 28396 23607
rect 30374 23604 30380 23616
rect 30432 23604 30438 23656
rect 31110 23644 31116 23656
rect 31071 23616 31116 23644
rect 31110 23604 31116 23616
rect 31168 23604 31174 23656
rect 27488 23548 28396 23576
rect 27488 23536 27494 23548
rect 22235 23480 24716 23508
rect 22235 23477 22247 23480
rect 22189 23471 22247 23477
rect 24762 23468 24768 23520
rect 24820 23508 24826 23520
rect 25041 23511 25099 23517
rect 25041 23508 25053 23511
rect 24820 23480 25053 23508
rect 24820 23468 24826 23480
rect 25041 23477 25053 23480
rect 25087 23477 25099 23511
rect 25041 23471 25099 23477
rect 26234 23468 26240 23520
rect 26292 23508 26298 23520
rect 26329 23511 26387 23517
rect 26329 23508 26341 23511
rect 26292 23480 26341 23508
rect 26292 23468 26298 23480
rect 26329 23477 26341 23480
rect 26375 23477 26387 23511
rect 26329 23471 26387 23477
rect 1104 23418 32016 23440
rect 1104 23366 2136 23418
rect 2188 23366 12440 23418
rect 12492 23366 22744 23418
rect 22796 23366 32016 23418
rect 1104 23344 32016 23366
rect 2590 23304 2596 23316
rect 2551 23276 2596 23304
rect 2590 23264 2596 23276
rect 2648 23264 2654 23316
rect 4341 23307 4399 23313
rect 4341 23273 4353 23307
rect 4387 23304 4399 23307
rect 4798 23304 4804 23316
rect 4387 23276 4804 23304
rect 4387 23273 4399 23276
rect 4341 23267 4399 23273
rect 4798 23264 4804 23276
rect 4856 23304 4862 23316
rect 5350 23304 5356 23316
rect 4856 23276 5356 23304
rect 4856 23264 4862 23276
rect 5350 23264 5356 23276
rect 5408 23264 5414 23316
rect 8018 23304 8024 23316
rect 7979 23276 8024 23304
rect 8018 23264 8024 23276
rect 8076 23264 8082 23316
rect 8202 23264 8208 23316
rect 8260 23304 8266 23316
rect 10045 23307 10103 23313
rect 10045 23304 10057 23307
rect 8260 23276 10057 23304
rect 8260 23264 8266 23276
rect 10045 23273 10057 23276
rect 10091 23273 10103 23307
rect 10045 23267 10103 23273
rect 12437 23307 12495 23313
rect 12437 23273 12449 23307
rect 12483 23304 12495 23307
rect 12526 23304 12532 23316
rect 12483 23276 12532 23304
rect 12483 23273 12495 23276
rect 12437 23267 12495 23273
rect 12526 23264 12532 23276
rect 12584 23264 12590 23316
rect 13354 23264 13360 23316
rect 13412 23304 13418 23316
rect 14918 23304 14924 23316
rect 13412 23276 14924 23304
rect 13412 23264 13418 23276
rect 14918 23264 14924 23276
rect 14976 23264 14982 23316
rect 17678 23304 17684 23316
rect 15120 23276 17684 23304
rect 3970 23196 3976 23248
rect 4028 23236 4034 23248
rect 8036 23236 8064 23264
rect 4028 23208 8064 23236
rect 4028 23196 4034 23208
rect 8294 23196 8300 23248
rect 8352 23236 8358 23248
rect 10778 23236 10784 23248
rect 8352 23208 10784 23236
rect 8352 23196 8358 23208
rect 10778 23196 10784 23208
rect 10836 23196 10842 23248
rect 13538 23196 13544 23248
rect 13596 23236 13602 23248
rect 13596 23208 14412 23236
rect 13596 23196 13602 23208
rect 3786 23168 3792 23180
rect 2792 23140 3792 23168
rect 2792 23109 2820 23140
rect 3786 23128 3792 23140
rect 3844 23128 3850 23180
rect 4430 23168 4436 23180
rect 4391 23140 4436 23168
rect 4430 23128 4436 23140
rect 4488 23128 4494 23180
rect 5258 23128 5264 23180
rect 5316 23168 5322 23180
rect 6730 23168 6736 23180
rect 5316 23140 6040 23168
rect 5316 23128 5322 23140
rect 2777 23103 2835 23109
rect 2777 23069 2789 23103
rect 2823 23069 2835 23103
rect 3050 23100 3056 23112
rect 3011 23072 3056 23100
rect 2777 23063 2835 23069
rect 3050 23060 3056 23072
rect 3108 23060 3114 23112
rect 4154 23100 4160 23112
rect 4115 23072 4160 23100
rect 4154 23060 4160 23072
rect 4212 23060 4218 23112
rect 5077 23103 5135 23109
rect 5077 23069 5089 23103
rect 5123 23100 5135 23103
rect 5350 23100 5356 23112
rect 5123 23072 5356 23100
rect 5123 23069 5135 23072
rect 5077 23063 5135 23069
rect 5350 23060 5356 23072
rect 5408 23060 5414 23112
rect 5721 23103 5779 23109
rect 5721 23069 5733 23103
rect 5767 23100 5779 23103
rect 5810 23100 5816 23112
rect 5767 23072 5816 23100
rect 5767 23069 5779 23072
rect 5721 23063 5779 23069
rect 5810 23060 5816 23072
rect 5868 23060 5874 23112
rect 6012 23109 6040 23140
rect 6196 23140 6736 23168
rect 6196 23109 6224 23140
rect 6730 23128 6736 23140
rect 6788 23168 6794 23180
rect 6917 23171 6975 23177
rect 6917 23168 6929 23171
rect 6788 23140 6929 23168
rect 6788 23128 6794 23140
rect 6917 23137 6929 23140
rect 6963 23137 6975 23171
rect 6917 23131 6975 23137
rect 9493 23171 9551 23177
rect 9493 23137 9505 23171
rect 9539 23168 9551 23171
rect 10505 23171 10563 23177
rect 9539 23140 10456 23168
rect 9539 23137 9551 23140
rect 9493 23131 9551 23137
rect 5997 23103 6055 23109
rect 5997 23069 6009 23103
rect 6043 23069 6055 23103
rect 5997 23063 6055 23069
rect 6181 23103 6239 23109
rect 6181 23069 6193 23103
rect 6227 23069 6239 23103
rect 6638 23100 6644 23112
rect 6599 23072 6644 23100
rect 6181 23063 6239 23069
rect 6638 23060 6644 23072
rect 6696 23060 6702 23112
rect 7926 23100 7932 23112
rect 7887 23072 7932 23100
rect 7926 23060 7932 23072
rect 7984 23060 7990 23112
rect 9306 23100 9312 23112
rect 9267 23072 9312 23100
rect 9306 23060 9312 23072
rect 9364 23060 9370 23112
rect 9582 23100 9588 23112
rect 9543 23072 9588 23100
rect 9582 23060 9588 23072
rect 9640 23060 9646 23112
rect 10226 23100 10232 23112
rect 10187 23072 10232 23100
rect 10226 23060 10232 23072
rect 10284 23060 10290 23112
rect 10428 23109 10456 23140
rect 10505 23137 10517 23171
rect 10551 23168 10563 23171
rect 10870 23168 10876 23180
rect 10551 23140 10876 23168
rect 10551 23137 10563 23140
rect 10505 23131 10563 23137
rect 10870 23128 10876 23140
rect 10928 23128 10934 23180
rect 12897 23171 12955 23177
rect 12897 23137 12909 23171
rect 12943 23168 12955 23171
rect 14384 23168 14412 23208
rect 14642 23196 14648 23248
rect 14700 23236 14706 23248
rect 15120 23236 15148 23276
rect 17678 23264 17684 23276
rect 17736 23264 17742 23316
rect 19426 23304 19432 23316
rect 19260 23276 19432 23304
rect 14700 23208 15148 23236
rect 14700 23196 14706 23208
rect 15194 23196 15200 23248
rect 15252 23236 15258 23248
rect 15381 23239 15439 23245
rect 15381 23236 15393 23239
rect 15252 23208 15393 23236
rect 15252 23196 15258 23208
rect 15381 23205 15393 23208
rect 15427 23205 15439 23239
rect 16485 23239 16543 23245
rect 16485 23236 16497 23239
rect 15381 23199 15439 23205
rect 15488 23208 16497 23236
rect 15488 23168 15516 23208
rect 16485 23205 16497 23208
rect 16531 23205 16543 23239
rect 16485 23199 16543 23205
rect 17310 23196 17316 23248
rect 17368 23236 17374 23248
rect 19260 23236 19288 23276
rect 19426 23264 19432 23276
rect 19484 23264 19490 23316
rect 19886 23264 19892 23316
rect 19944 23304 19950 23316
rect 23474 23304 23480 23316
rect 19944 23276 23480 23304
rect 19944 23264 19950 23276
rect 23474 23264 23480 23276
rect 23532 23264 23538 23316
rect 23661 23307 23719 23313
rect 23661 23273 23673 23307
rect 23707 23304 23719 23307
rect 24670 23304 24676 23316
rect 23707 23276 24676 23304
rect 23707 23273 23719 23276
rect 23661 23267 23719 23273
rect 24670 23264 24676 23276
rect 24728 23264 24734 23316
rect 24946 23264 24952 23316
rect 25004 23304 25010 23316
rect 25041 23307 25099 23313
rect 25041 23304 25053 23307
rect 25004 23276 25053 23304
rect 25004 23264 25010 23276
rect 25041 23273 25053 23276
rect 25087 23273 25099 23307
rect 27982 23304 27988 23316
rect 27943 23276 27988 23304
rect 25041 23267 25099 23273
rect 27982 23264 27988 23276
rect 28040 23264 28046 23316
rect 17368 23208 19288 23236
rect 25225 23239 25283 23245
rect 17368 23196 17374 23208
rect 25225 23205 25237 23239
rect 25271 23236 25283 23239
rect 29178 23236 29184 23248
rect 25271 23208 29184 23236
rect 25271 23205 25283 23208
rect 25225 23199 25283 23205
rect 29178 23196 29184 23208
rect 29236 23196 29242 23248
rect 12943 23140 14320 23168
rect 14384 23140 15516 23168
rect 15841 23171 15899 23177
rect 12943 23137 12955 23140
rect 12897 23131 12955 23137
rect 10413 23103 10471 23109
rect 10413 23069 10425 23103
rect 10459 23100 10471 23103
rect 10778 23100 10784 23112
rect 10459 23072 10784 23100
rect 10459 23069 10471 23072
rect 10413 23063 10471 23069
rect 10778 23060 10784 23072
rect 10836 23060 10842 23112
rect 11057 23103 11115 23109
rect 11057 23069 11069 23103
rect 11103 23100 11115 23103
rect 12802 23100 12808 23112
rect 11103 23072 12808 23100
rect 11103 23069 11115 23072
rect 11057 23063 11115 23069
rect 12802 23060 12808 23072
rect 12860 23060 12866 23112
rect 13081 23103 13139 23109
rect 13081 23069 13093 23103
rect 13127 23069 13139 23103
rect 13081 23063 13139 23069
rect 1857 23035 1915 23041
rect 1857 23032 1869 23035
rect 768 23004 1869 23032
rect 768 22828 796 23004
rect 1857 23001 1869 23004
rect 1903 23001 1915 23035
rect 1857 22995 1915 23001
rect 2041 23035 2099 23041
rect 2041 23001 2053 23035
rect 2087 23032 2099 23035
rect 2222 23032 2228 23044
rect 2087 23004 2228 23032
rect 2087 23001 2099 23004
rect 2041 22995 2099 23001
rect 2222 22992 2228 23004
rect 2280 22992 2286 23044
rect 2958 23032 2964 23044
rect 2919 23004 2964 23032
rect 2958 22992 2964 23004
rect 3016 22992 3022 23044
rect 10962 23032 10968 23044
rect 4908 23004 10968 23032
rect 3973 22967 4031 22973
rect 3973 22933 3985 22967
rect 4019 22964 4031 22967
rect 4154 22964 4160 22976
rect 4019 22936 4160 22964
rect 4019 22933 4031 22936
rect 3973 22927 4031 22933
rect 4154 22924 4160 22936
rect 4212 22924 4218 22976
rect 4908 22973 4936 23004
rect 10962 22992 10968 23004
rect 11020 22992 11026 23044
rect 11324 23035 11382 23041
rect 11324 23001 11336 23035
rect 11370 23032 11382 23035
rect 12158 23032 12164 23044
rect 11370 23004 12164 23032
rect 11370 23001 11382 23004
rect 11324 22995 11382 23001
rect 12158 22992 12164 23004
rect 12216 22992 12222 23044
rect 12250 22992 12256 23044
rect 12308 23032 12314 23044
rect 13096 23032 13124 23063
rect 13170 23060 13176 23112
rect 13228 23100 13234 23112
rect 13357 23103 13415 23109
rect 13357 23100 13369 23103
rect 13228 23072 13369 23100
rect 13228 23060 13234 23072
rect 13357 23069 13369 23072
rect 13403 23069 13415 23103
rect 13357 23063 13415 23069
rect 13541 23103 13599 23109
rect 13541 23069 13553 23103
rect 13587 23100 13599 23103
rect 13722 23100 13728 23112
rect 13587 23072 13728 23100
rect 13587 23069 13599 23072
rect 13541 23063 13599 23069
rect 12308 23004 13124 23032
rect 12308 22992 12314 23004
rect 13556 22976 13584 23063
rect 13722 23060 13728 23072
rect 13780 23060 13786 23112
rect 14292 23109 14320 23140
rect 15841 23137 15853 23171
rect 15887 23168 15899 23171
rect 16206 23168 16212 23180
rect 15887 23140 16212 23168
rect 15887 23137 15899 23140
rect 15841 23131 15899 23137
rect 16206 23128 16212 23140
rect 16264 23128 16270 23180
rect 18230 23168 18236 23180
rect 16776 23140 18236 23168
rect 14277 23103 14335 23109
rect 14277 23069 14289 23103
rect 14323 23069 14335 23103
rect 14277 23063 14335 23069
rect 14461 23103 14519 23109
rect 14461 23069 14473 23103
rect 14507 23069 14519 23103
rect 14461 23063 14519 23069
rect 14553 23103 14611 23109
rect 14553 23069 14565 23103
rect 14599 23100 14611 23103
rect 14734 23100 14740 23112
rect 14599 23072 14740 23100
rect 14599 23069 14611 23072
rect 14553 23063 14611 23069
rect 13814 22992 13820 23044
rect 13872 23032 13878 23044
rect 14476 23032 14504 23063
rect 14734 23060 14740 23072
rect 14792 23060 14798 23112
rect 16485 23103 16543 23109
rect 16485 23100 16497 23103
rect 14835 23072 16497 23100
rect 14835 23032 14863 23072
rect 16485 23069 16497 23072
rect 16531 23069 16543 23103
rect 16666 23100 16672 23112
rect 16627 23072 16672 23100
rect 16485 23063 16543 23069
rect 16666 23060 16672 23072
rect 16724 23060 16730 23112
rect 16776 23109 16804 23140
rect 18230 23128 18236 23140
rect 18288 23128 18294 23180
rect 20898 23128 20904 23180
rect 20956 23168 20962 23180
rect 21082 23168 21088 23180
rect 20956 23140 21088 23168
rect 20956 23128 20962 23140
rect 21082 23128 21088 23140
rect 21140 23128 21146 23180
rect 24118 23128 24124 23180
rect 24176 23168 24182 23180
rect 25961 23171 26019 23177
rect 25961 23168 25973 23171
rect 24176 23140 25973 23168
rect 24176 23128 24182 23140
rect 25961 23137 25973 23140
rect 26007 23137 26019 23171
rect 25961 23131 26019 23137
rect 27154 23128 27160 23180
rect 27212 23168 27218 23180
rect 27212 23140 27568 23168
rect 27212 23128 27218 23140
rect 16761 23103 16819 23109
rect 16761 23069 16773 23103
rect 16807 23069 16819 23103
rect 16761 23063 16819 23069
rect 17034 23060 17040 23112
rect 17092 23100 17098 23112
rect 17865 23103 17923 23109
rect 17865 23100 17877 23103
rect 17092 23072 17877 23100
rect 17092 23060 17098 23072
rect 17865 23069 17877 23072
rect 17911 23069 17923 23103
rect 18138 23100 18144 23112
rect 18099 23072 18144 23100
rect 17865 23063 17923 23069
rect 18138 23060 18144 23072
rect 18196 23060 18202 23112
rect 18322 23100 18328 23112
rect 18283 23072 18328 23100
rect 18322 23060 18328 23072
rect 18380 23060 18386 23112
rect 19242 23100 19248 23112
rect 19203 23072 19248 23100
rect 19242 23060 19248 23072
rect 19300 23060 19306 23112
rect 19334 23060 19340 23112
rect 19392 23100 19398 23112
rect 19501 23103 19559 23109
rect 19501 23100 19513 23103
rect 19392 23072 19513 23100
rect 19392 23060 19398 23072
rect 19501 23069 19513 23072
rect 19547 23069 19559 23103
rect 19501 23063 19559 23069
rect 25130 23060 25136 23112
rect 25188 23060 25194 23112
rect 26789 23103 26847 23109
rect 26789 23069 26801 23103
rect 26835 23069 26847 23103
rect 26789 23063 26847 23069
rect 27065 23103 27123 23109
rect 27065 23069 27077 23103
rect 27111 23069 27123 23103
rect 27246 23100 27252 23112
rect 27207 23072 27252 23100
rect 27065 23063 27123 23069
rect 13872 23004 14504 23032
rect 14568 23004 14863 23032
rect 13872 22992 13878 23004
rect 4893 22967 4951 22973
rect 4893 22933 4905 22967
rect 4939 22933 4951 22967
rect 4893 22927 4951 22933
rect 5442 22924 5448 22976
rect 5500 22964 5506 22976
rect 5537 22967 5595 22973
rect 5537 22964 5549 22967
rect 5500 22936 5549 22964
rect 5500 22924 5506 22936
rect 5537 22933 5549 22936
rect 5583 22933 5595 22967
rect 5537 22927 5595 22933
rect 6454 22924 6460 22976
rect 6512 22964 6518 22976
rect 7098 22964 7104 22976
rect 6512 22936 7104 22964
rect 6512 22924 6518 22936
rect 7098 22924 7104 22936
rect 7156 22924 7162 22976
rect 7834 22924 7840 22976
rect 7892 22964 7898 22976
rect 8389 22967 8447 22973
rect 8389 22964 8401 22967
rect 7892 22936 8401 22964
rect 7892 22924 7898 22936
rect 8389 22933 8401 22936
rect 8435 22933 8447 22967
rect 9122 22964 9128 22976
rect 9083 22936 9128 22964
rect 8389 22927 8447 22933
rect 9122 22924 9128 22936
rect 9180 22924 9186 22976
rect 12894 22924 12900 22976
rect 12952 22964 12958 22976
rect 13538 22964 13544 22976
rect 12952 22936 13544 22964
rect 12952 22924 12958 22936
rect 13538 22924 13544 22936
rect 13596 22924 13602 22976
rect 14090 22964 14096 22976
rect 14051 22936 14096 22964
rect 14090 22924 14096 22936
rect 14148 22924 14154 22976
rect 14366 22924 14372 22976
rect 14424 22964 14430 22976
rect 14568 22964 14596 23004
rect 15746 22992 15752 23044
rect 15804 23032 15810 23044
rect 15933 23035 15991 23041
rect 15933 23032 15945 23035
rect 15804 23004 15945 23032
rect 15804 22992 15810 23004
rect 15933 23001 15945 23004
rect 15979 23001 15991 23035
rect 19978 23032 19984 23044
rect 15933 22995 15991 23001
rect 16684 23004 19984 23032
rect 16684 22976 16712 23004
rect 19978 22992 19984 23004
rect 20036 22992 20042 23044
rect 20714 22992 20720 23044
rect 20772 23032 20778 23044
rect 21330 23035 21388 23041
rect 21330 23032 21342 23035
rect 20772 23004 21342 23032
rect 20772 22992 20778 23004
rect 21330 23001 21342 23004
rect 21376 23001 21388 23035
rect 21330 22995 21388 23001
rect 23382 22992 23388 23044
rect 23440 23032 23446 23044
rect 23477 23035 23535 23041
rect 23477 23032 23489 23035
rect 23440 23004 23489 23032
rect 23440 22992 23446 23004
rect 23477 23001 23489 23004
rect 23523 23001 23535 23035
rect 23477 22995 23535 23001
rect 23693 23035 23751 23041
rect 23693 23001 23705 23035
rect 23739 23032 23751 23035
rect 24302 23032 24308 23044
rect 23739 23004 24308 23032
rect 23739 23001 23751 23004
rect 23693 22995 23751 23001
rect 24302 22992 24308 23004
rect 24360 22992 24366 23044
rect 24857 23035 24915 23041
rect 24857 23001 24869 23035
rect 24903 23032 24915 23035
rect 25148 23032 25176 23060
rect 25774 23032 25780 23044
rect 24903 23004 25176 23032
rect 25735 23004 25780 23032
rect 24903 23001 24915 23004
rect 24857 22995 24915 23001
rect 25774 22992 25780 23004
rect 25832 22992 25838 23044
rect 15838 22964 15844 22976
rect 14424 22936 14596 22964
rect 15799 22936 15844 22964
rect 14424 22924 14430 22936
rect 15838 22924 15844 22936
rect 15896 22924 15902 22976
rect 16666 22924 16672 22976
rect 16724 22924 16730 22976
rect 17681 22967 17739 22973
rect 17681 22933 17693 22967
rect 17727 22964 17739 22967
rect 17862 22964 17868 22976
rect 17727 22936 17868 22964
rect 17727 22933 17739 22936
rect 17681 22927 17739 22933
rect 17862 22924 17868 22936
rect 17920 22924 17926 22976
rect 18230 22924 18236 22976
rect 18288 22964 18294 22976
rect 19794 22964 19800 22976
rect 18288 22936 19800 22964
rect 18288 22924 18294 22936
rect 19794 22924 19800 22936
rect 19852 22964 19858 22976
rect 20625 22967 20683 22973
rect 20625 22964 20637 22967
rect 19852 22936 20637 22964
rect 19852 22924 19858 22936
rect 20625 22933 20637 22936
rect 20671 22933 20683 22967
rect 22462 22964 22468 22976
rect 22423 22936 22468 22964
rect 20625 22927 20683 22933
rect 22462 22924 22468 22936
rect 22520 22924 22526 22976
rect 23845 22967 23903 22973
rect 23845 22933 23857 22967
rect 23891 22964 23903 22967
rect 23934 22964 23940 22976
rect 23891 22936 23940 22964
rect 23891 22933 23903 22936
rect 23845 22927 23903 22933
rect 23934 22924 23940 22936
rect 23992 22924 23998 22976
rect 25038 22924 25044 22976
rect 25096 22973 25102 22976
rect 25096 22967 25115 22973
rect 25103 22933 25115 22967
rect 25096 22927 25115 22933
rect 25096 22924 25102 22927
rect 26142 22924 26148 22976
rect 26200 22964 26206 22976
rect 26605 22967 26663 22973
rect 26605 22964 26617 22967
rect 26200 22936 26617 22964
rect 26200 22924 26206 22936
rect 26605 22933 26617 22936
rect 26651 22933 26663 22967
rect 26804 22964 26832 23063
rect 27080 23032 27108 23063
rect 27246 23060 27252 23072
rect 27304 23060 27310 23112
rect 27540 23100 27568 23140
rect 27798 23128 27804 23180
rect 27856 23168 27862 23180
rect 29917 23171 29975 23177
rect 29917 23168 29929 23171
rect 27856 23140 29929 23168
rect 27856 23128 27862 23140
rect 29917 23137 29929 23140
rect 29963 23137 29975 23171
rect 29917 23131 29975 23137
rect 28169 23103 28227 23109
rect 28169 23100 28181 23103
rect 27540 23072 28181 23100
rect 28169 23069 28181 23072
rect 28215 23069 28227 23103
rect 28169 23063 28227 23069
rect 28445 23103 28503 23109
rect 28445 23069 28457 23103
rect 28491 23069 28503 23103
rect 28445 23063 28503 23069
rect 28629 23103 28687 23109
rect 28629 23069 28641 23103
rect 28675 23100 28687 23103
rect 29454 23100 29460 23112
rect 28675 23072 29460 23100
rect 28675 23069 28687 23072
rect 28629 23063 28687 23069
rect 27430 23032 27436 23044
rect 27080 23004 27436 23032
rect 27430 22992 27436 23004
rect 27488 23032 27494 23044
rect 28460 23032 28488 23063
rect 29454 23060 29460 23072
rect 29512 23060 29518 23112
rect 27488 23004 28488 23032
rect 27488 22992 27494 23004
rect 29270 22992 29276 23044
rect 29328 23032 29334 23044
rect 30162 23035 30220 23041
rect 30162 23032 30174 23035
rect 29328 23004 30174 23032
rect 29328 22992 29334 23004
rect 30162 23001 30174 23004
rect 30208 23001 30220 23035
rect 30162 22995 30220 23001
rect 27154 22964 27160 22976
rect 26804 22936 27160 22964
rect 26605 22927 26663 22933
rect 27154 22924 27160 22936
rect 27212 22924 27218 22976
rect 30558 22924 30564 22976
rect 30616 22964 30622 22976
rect 31294 22964 31300 22976
rect 30616 22936 31300 22964
rect 30616 22924 30622 22936
rect 31294 22924 31300 22936
rect 31352 22924 31358 22976
rect 1104 22874 32016 22896
rect 768 22800 888 22828
rect 1104 22822 7288 22874
rect 7340 22822 17592 22874
rect 17644 22822 27896 22874
rect 27948 22822 32016 22874
rect 1104 22800 32016 22822
rect 0 22692 800 22706
rect 860 22692 888 22800
rect 1486 22760 1492 22772
rect 1447 22732 1492 22760
rect 1486 22720 1492 22732
rect 1544 22720 1550 22772
rect 1670 22720 1676 22772
rect 1728 22720 1734 22772
rect 2409 22763 2467 22769
rect 2409 22729 2421 22763
rect 2455 22760 2467 22763
rect 3050 22760 3056 22772
rect 2455 22732 3056 22760
rect 2455 22729 2467 22732
rect 2409 22723 2467 22729
rect 3050 22720 3056 22732
rect 3108 22720 3114 22772
rect 6638 22720 6644 22772
rect 6696 22760 6702 22772
rect 7745 22763 7803 22769
rect 7745 22760 7757 22763
rect 6696 22732 7757 22760
rect 6696 22720 6702 22732
rect 7745 22729 7757 22732
rect 7791 22729 7803 22763
rect 7745 22723 7803 22729
rect 8266 22732 9260 22760
rect 0 22664 888 22692
rect 1688 22692 1716 22720
rect 2777 22695 2835 22701
rect 1688 22664 1900 22692
rect 0 22650 800 22664
rect 1670 22624 1676 22636
rect 1631 22596 1676 22624
rect 1670 22584 1676 22596
rect 1728 22584 1734 22636
rect 1872 22633 1900 22664
rect 2777 22661 2789 22695
rect 2823 22692 2835 22695
rect 4798 22692 4804 22704
rect 2823 22664 2912 22692
rect 4759 22664 4804 22692
rect 2823 22661 2835 22664
rect 2777 22655 2835 22661
rect 1857 22627 1915 22633
rect 1857 22593 1869 22627
rect 1903 22593 1915 22627
rect 2884 22624 2912 22664
rect 4798 22652 4804 22664
rect 4856 22692 4862 22704
rect 6822 22692 6828 22704
rect 4856 22664 5672 22692
rect 4856 22652 4862 22664
rect 3418 22624 3424 22636
rect 2884 22596 3424 22624
rect 1857 22587 1915 22593
rect 1872 22420 1900 22587
rect 3418 22584 3424 22596
rect 3476 22584 3482 22636
rect 3786 22624 3792 22636
rect 3747 22596 3792 22624
rect 3786 22584 3792 22596
rect 3844 22584 3850 22636
rect 4062 22624 4068 22636
rect 4023 22596 4068 22624
rect 4062 22584 4068 22596
rect 4120 22584 4126 22636
rect 4614 22624 4620 22636
rect 4575 22596 4620 22624
rect 4614 22584 4620 22596
rect 4672 22584 4678 22636
rect 5442 22624 5448 22636
rect 5403 22596 5448 22624
rect 5442 22584 5448 22596
rect 5500 22584 5506 22636
rect 5644 22633 5672 22664
rect 6380 22664 6828 22692
rect 6380 22633 6408 22664
rect 6822 22652 6828 22664
rect 6880 22652 6886 22704
rect 7650 22652 7656 22704
rect 7708 22692 7714 22704
rect 8266 22692 8294 22732
rect 7708 22664 8294 22692
rect 8472 22695 8530 22701
rect 7708 22652 7714 22664
rect 8472 22661 8484 22695
rect 8518 22692 8530 22695
rect 9122 22692 9128 22704
rect 8518 22664 9128 22692
rect 8518 22661 8530 22664
rect 8472 22655 8530 22661
rect 9122 22652 9128 22664
rect 9180 22652 9186 22704
rect 9232 22692 9260 22732
rect 9306 22720 9312 22772
rect 9364 22760 9370 22772
rect 10045 22763 10103 22769
rect 10045 22760 10057 22763
rect 9364 22732 10057 22760
rect 9364 22720 9370 22732
rect 10045 22729 10057 22732
rect 10091 22729 10103 22763
rect 10045 22723 10103 22729
rect 10134 22720 10140 22772
rect 10192 22760 10198 22772
rect 11333 22763 11391 22769
rect 11333 22760 11345 22763
rect 10192 22732 11345 22760
rect 10192 22720 10198 22732
rect 11333 22729 11345 22732
rect 11379 22729 11391 22763
rect 11333 22723 11391 22729
rect 12066 22720 12072 22772
rect 12124 22760 12130 22772
rect 13446 22760 13452 22772
rect 12124 22732 13452 22760
rect 12124 22720 12130 22732
rect 13446 22720 13452 22732
rect 13504 22720 13510 22772
rect 13538 22720 13544 22772
rect 13596 22760 13602 22772
rect 14185 22763 14243 22769
rect 14185 22760 14197 22763
rect 13596 22732 14197 22760
rect 13596 22720 13602 22732
rect 14185 22729 14197 22732
rect 14231 22729 14243 22763
rect 15102 22760 15108 22772
rect 15063 22732 15108 22760
rect 14185 22723 14243 22729
rect 15102 22720 15108 22732
rect 15160 22720 15166 22772
rect 16574 22720 16580 22772
rect 16632 22760 16638 22772
rect 17126 22760 17132 22772
rect 16632 22732 17132 22760
rect 16632 22720 16638 22732
rect 17126 22720 17132 22732
rect 17184 22720 17190 22772
rect 17494 22720 17500 22772
rect 17552 22760 17558 22772
rect 17681 22763 17739 22769
rect 17681 22760 17693 22763
rect 17552 22732 17693 22760
rect 17552 22720 17558 22732
rect 17681 22729 17693 22732
rect 17727 22729 17739 22763
rect 18782 22760 18788 22772
rect 18743 22732 18788 22760
rect 17681 22723 17739 22729
rect 18782 22720 18788 22732
rect 18840 22720 18846 22772
rect 19886 22760 19892 22772
rect 18892 22732 19892 22760
rect 13072 22695 13130 22701
rect 9232 22664 10824 22692
rect 5629 22627 5687 22633
rect 5629 22593 5641 22627
rect 5675 22593 5687 22627
rect 5629 22587 5687 22593
rect 6365 22627 6423 22633
rect 6365 22593 6377 22627
rect 6411 22593 6423 22627
rect 6621 22627 6679 22633
rect 6621 22624 6633 22627
rect 6365 22587 6423 22593
rect 6472 22596 6633 22624
rect 1949 22559 2007 22565
rect 1949 22525 1961 22559
rect 1995 22556 2007 22559
rect 2590 22556 2596 22568
rect 1995 22528 2596 22556
rect 1995 22525 2007 22528
rect 1949 22519 2007 22525
rect 2590 22516 2596 22528
rect 2648 22516 2654 22568
rect 2869 22559 2927 22565
rect 2869 22525 2881 22559
rect 2915 22525 2927 22559
rect 2869 22519 2927 22525
rect 2222 22448 2228 22500
rect 2280 22488 2286 22500
rect 2884 22488 2912 22519
rect 3050 22516 3056 22568
rect 3108 22556 3114 22568
rect 4246 22556 4252 22568
rect 3108 22528 3153 22556
rect 3252 22528 4252 22556
rect 3108 22516 3114 22528
rect 3252 22488 3280 22528
rect 4246 22516 4252 22528
rect 4304 22516 4310 22568
rect 5721 22559 5779 22565
rect 5721 22525 5733 22559
rect 5767 22556 5779 22559
rect 5902 22556 5908 22568
rect 5767 22528 5908 22556
rect 5767 22525 5779 22528
rect 5721 22519 5779 22525
rect 5902 22516 5908 22528
rect 5960 22516 5966 22568
rect 6472 22556 6500 22596
rect 6621 22593 6633 22596
rect 6667 22593 6679 22627
rect 6621 22587 6679 22593
rect 8110 22584 8116 22636
rect 8168 22624 8174 22636
rect 8205 22627 8263 22633
rect 8205 22624 8217 22627
rect 8168 22596 8217 22624
rect 8168 22584 8174 22596
rect 8205 22593 8217 22596
rect 8251 22593 8263 22627
rect 8205 22587 8263 22593
rect 9766 22584 9772 22636
rect 9824 22624 9830 22636
rect 9950 22624 9956 22636
rect 9824 22596 9956 22624
rect 9824 22584 9830 22596
rect 9950 22584 9956 22596
rect 10008 22624 10014 22636
rect 10229 22627 10287 22633
rect 10229 22624 10241 22627
rect 10008 22596 10241 22624
rect 10008 22584 10014 22596
rect 10229 22593 10241 22596
rect 10275 22593 10287 22627
rect 10229 22587 10287 22593
rect 10318 22584 10324 22636
rect 10376 22624 10382 22636
rect 10505 22627 10563 22633
rect 10505 22624 10517 22627
rect 10376 22596 10517 22624
rect 10376 22584 10382 22596
rect 10505 22593 10517 22596
rect 10551 22593 10563 22627
rect 10505 22587 10563 22593
rect 10689 22627 10747 22633
rect 10689 22593 10701 22627
rect 10735 22593 10747 22627
rect 10689 22587 10747 22593
rect 6380 22528 6500 22556
rect 3973 22491 4031 22497
rect 3973 22488 3985 22491
rect 2280 22460 3280 22488
rect 3436 22460 3985 22488
rect 2280 22448 2286 22460
rect 3436 22420 3464 22460
rect 3973 22457 3985 22460
rect 4019 22488 4031 22491
rect 4982 22488 4988 22500
rect 4019 22460 4988 22488
rect 4019 22457 4031 22460
rect 3973 22451 4031 22457
rect 4982 22448 4988 22460
rect 5040 22448 5046 22500
rect 5261 22491 5319 22497
rect 5261 22457 5273 22491
rect 5307 22488 5319 22491
rect 6380 22488 6408 22528
rect 5307 22460 6408 22488
rect 9585 22491 9643 22497
rect 5307 22457 5319 22460
rect 5261 22451 5319 22457
rect 9585 22457 9597 22491
rect 9631 22488 9643 22491
rect 9674 22488 9680 22500
rect 9631 22460 9680 22488
rect 9631 22457 9643 22460
rect 9585 22451 9643 22457
rect 9674 22448 9680 22460
rect 9732 22488 9738 22500
rect 10704 22488 10732 22587
rect 10796 22556 10824 22664
rect 13072 22661 13084 22695
rect 13118 22692 13130 22695
rect 14090 22692 14096 22704
rect 13118 22664 14096 22692
rect 13118 22661 13130 22664
rect 13072 22655 13130 22661
rect 14090 22652 14096 22664
rect 14148 22652 14154 22704
rect 14274 22652 14280 22704
rect 14332 22692 14338 22704
rect 17770 22692 17776 22704
rect 14332 22664 17776 22692
rect 14332 22652 14338 22664
rect 17770 22652 17776 22664
rect 17828 22652 17834 22704
rect 18892 22692 18920 22732
rect 19886 22720 19892 22732
rect 19944 22720 19950 22772
rect 20714 22760 20720 22772
rect 20675 22732 20720 22760
rect 20714 22720 20720 22732
rect 20772 22720 20778 22772
rect 21174 22720 21180 22772
rect 21232 22760 21238 22772
rect 21450 22760 21456 22772
rect 21232 22732 21456 22760
rect 21232 22720 21238 22732
rect 21450 22720 21456 22732
rect 21508 22720 21514 22772
rect 21910 22720 21916 22772
rect 21968 22720 21974 22772
rect 24302 22720 24308 22772
rect 24360 22760 24366 22772
rect 24578 22760 24584 22772
rect 24360 22732 24584 22760
rect 24360 22720 24366 22732
rect 24578 22720 24584 22732
rect 24636 22720 24642 22772
rect 26418 22720 26424 22772
rect 26476 22760 26482 22772
rect 27157 22763 27215 22769
rect 27157 22760 27169 22763
rect 26476 22732 27169 22760
rect 26476 22720 26482 22732
rect 27157 22729 27169 22732
rect 27203 22729 27215 22763
rect 27157 22723 27215 22729
rect 29181 22763 29239 22769
rect 29181 22729 29193 22763
rect 29227 22760 29239 22763
rect 29454 22760 29460 22772
rect 29227 22732 29460 22760
rect 29227 22729 29239 22732
rect 29181 22723 29239 22729
rect 29454 22720 29460 22732
rect 29512 22720 29518 22772
rect 29822 22720 29828 22772
rect 29880 22760 29886 22772
rect 29917 22763 29975 22769
rect 29917 22760 29929 22763
rect 29880 22732 29929 22760
rect 29880 22720 29886 22732
rect 29917 22729 29929 22732
rect 29963 22729 29975 22763
rect 29917 22723 29975 22729
rect 18616 22664 18920 22692
rect 19245 22695 19303 22701
rect 10962 22584 10968 22636
rect 11020 22624 11026 22636
rect 15286 22624 15292 22636
rect 11020 22596 15194 22624
rect 15247 22596 15292 22624
rect 11020 22584 11026 22596
rect 11146 22556 11152 22568
rect 10796 22528 11152 22556
rect 11146 22516 11152 22528
rect 11204 22556 11210 22568
rect 11517 22559 11575 22565
rect 11517 22556 11529 22559
rect 11204 22528 11529 22556
rect 11204 22516 11210 22528
rect 11517 22525 11529 22528
rect 11563 22525 11575 22559
rect 11517 22519 11575 22525
rect 11793 22559 11851 22565
rect 11793 22525 11805 22559
rect 11839 22556 11851 22559
rect 12250 22556 12256 22568
rect 11839 22528 12256 22556
rect 11839 22525 11851 22528
rect 11793 22519 11851 22525
rect 12250 22516 12256 22528
rect 12308 22516 12314 22568
rect 12802 22556 12808 22568
rect 12763 22528 12808 22556
rect 12802 22516 12808 22528
rect 12860 22516 12866 22568
rect 15166 22556 15194 22596
rect 15286 22584 15292 22596
rect 15344 22584 15350 22636
rect 15470 22584 15476 22636
rect 15528 22624 15534 22636
rect 15565 22627 15623 22633
rect 15565 22624 15577 22627
rect 15528 22596 15577 22624
rect 15528 22584 15534 22596
rect 15565 22593 15577 22596
rect 15611 22593 15623 22627
rect 15746 22624 15752 22636
rect 15707 22596 15752 22624
rect 15565 22587 15623 22593
rect 15746 22584 15752 22596
rect 15804 22584 15810 22636
rect 16758 22624 16764 22636
rect 16719 22596 16764 22624
rect 16758 22584 16764 22596
rect 16816 22584 16822 22636
rect 16942 22624 16948 22636
rect 16903 22596 16948 22624
rect 16942 22584 16948 22596
rect 17000 22584 17006 22636
rect 17129 22627 17187 22633
rect 17129 22593 17141 22627
rect 17175 22624 17187 22627
rect 17862 22624 17868 22636
rect 17175 22596 17724 22624
rect 17823 22596 17868 22624
rect 17175 22593 17187 22596
rect 17129 22587 17187 22593
rect 17034 22556 17040 22568
rect 15166 22528 17040 22556
rect 17034 22516 17040 22528
rect 17092 22516 17098 22568
rect 11238 22488 11244 22500
rect 9732 22460 11244 22488
rect 9732 22448 9738 22460
rect 11238 22448 11244 22460
rect 11296 22448 11302 22500
rect 11333 22491 11391 22497
rect 11333 22457 11345 22491
rect 11379 22488 11391 22491
rect 11379 22460 12848 22488
rect 11379 22457 11391 22460
rect 11333 22451 11391 22457
rect 3602 22420 3608 22432
rect 1872 22392 3464 22420
rect 3563 22392 3608 22420
rect 3602 22380 3608 22392
rect 3660 22380 3666 22432
rect 5810 22380 5816 22432
rect 5868 22420 5874 22432
rect 6730 22420 6736 22432
rect 5868 22392 6736 22420
rect 5868 22380 5874 22392
rect 6730 22380 6736 22392
rect 6788 22380 6794 22432
rect 10502 22380 10508 22432
rect 10560 22420 10566 22432
rect 12618 22420 12624 22432
rect 10560 22392 12624 22420
rect 10560 22380 10566 22392
rect 12618 22380 12624 22392
rect 12676 22380 12682 22432
rect 12820 22420 12848 22460
rect 14090 22448 14096 22500
rect 14148 22488 14154 22500
rect 17144 22488 17172 22587
rect 17221 22559 17279 22565
rect 17221 22525 17233 22559
rect 17267 22525 17279 22559
rect 17696 22556 17724 22596
rect 17862 22584 17868 22596
rect 17920 22584 17926 22636
rect 18141 22627 18199 22633
rect 18141 22593 18153 22627
rect 18187 22624 18199 22627
rect 18230 22624 18236 22636
rect 18187 22596 18236 22624
rect 18187 22593 18199 22596
rect 18141 22587 18199 22593
rect 18230 22584 18236 22596
rect 18288 22584 18294 22636
rect 18414 22584 18420 22636
rect 18472 22624 18478 22636
rect 18616 22633 18644 22664
rect 19245 22661 19257 22695
rect 19291 22692 19303 22695
rect 21928 22692 21956 22720
rect 19291 22664 21956 22692
rect 19291 22661 19303 22664
rect 19245 22655 19303 22661
rect 22370 22652 22376 22704
rect 22428 22692 22434 22704
rect 23382 22692 23388 22704
rect 22428 22664 23388 22692
rect 22428 22652 22434 22664
rect 23382 22652 23388 22664
rect 23440 22652 23446 22704
rect 24670 22652 24676 22704
rect 24728 22692 24734 22704
rect 28074 22701 28080 22704
rect 26329 22695 26387 22701
rect 26329 22692 26341 22695
rect 24728 22664 26341 22692
rect 24728 22652 24734 22664
rect 26329 22661 26341 22664
rect 26375 22661 26387 22695
rect 26329 22655 26387 22661
rect 27065 22695 27123 22701
rect 27065 22661 27077 22695
rect 27111 22692 27123 22695
rect 28068 22692 28080 22701
rect 27111 22664 27936 22692
rect 28035 22664 28080 22692
rect 27111 22661 27123 22664
rect 27065 22655 27123 22661
rect 18601 22627 18659 22633
rect 18601 22624 18613 22627
rect 18472 22596 18613 22624
rect 18472 22584 18478 22596
rect 18601 22593 18613 22596
rect 18647 22593 18659 22627
rect 18601 22587 18659 22593
rect 18782 22584 18788 22636
rect 18840 22624 18846 22636
rect 19426 22624 19432 22636
rect 18840 22596 18885 22624
rect 19387 22596 19432 22624
rect 18840 22584 18846 22596
rect 19426 22584 19432 22596
rect 19484 22584 19490 22636
rect 19518 22584 19524 22636
rect 19576 22624 19582 22636
rect 19794 22624 19800 22636
rect 19576 22596 19669 22624
rect 19755 22596 19800 22624
rect 19576 22584 19582 22596
rect 19794 22584 19800 22596
rect 19852 22584 19858 22636
rect 20898 22624 20904 22636
rect 20859 22596 20904 22624
rect 20898 22584 20904 22596
rect 20956 22584 20962 22636
rect 21082 22584 21088 22636
rect 21140 22624 21146 22636
rect 21913 22627 21971 22633
rect 21913 22624 21925 22627
rect 21140 22596 21925 22624
rect 21140 22584 21146 22596
rect 21913 22593 21925 22596
rect 21959 22593 21971 22627
rect 21913 22587 21971 22593
rect 22002 22584 22008 22636
rect 22060 22624 22066 22636
rect 22169 22627 22227 22633
rect 22169 22624 22181 22627
rect 22060 22596 22181 22624
rect 22060 22584 22066 22596
rect 22169 22593 22181 22596
rect 22215 22593 22227 22627
rect 24210 22624 24216 22636
rect 24171 22596 24216 22624
rect 22169 22587 22227 22593
rect 24210 22584 24216 22596
rect 24268 22584 24274 22636
rect 24486 22633 24492 22636
rect 24480 22587 24492 22633
rect 24544 22624 24550 22636
rect 24544 22596 24580 22624
rect 24486 22584 24492 22587
rect 24544 22584 24550 22596
rect 25774 22584 25780 22636
rect 25832 22624 25838 22636
rect 26145 22627 26203 22633
rect 26145 22624 26157 22627
rect 25832 22596 26157 22624
rect 25832 22584 25838 22596
rect 26145 22593 26157 22596
rect 26191 22593 26203 22627
rect 27798 22624 27804 22636
rect 27759 22596 27804 22624
rect 26145 22587 26203 22593
rect 27798 22584 27804 22596
rect 27856 22584 27862 22636
rect 27908 22624 27936 22664
rect 28068 22655 28080 22664
rect 28074 22652 28080 22655
rect 28132 22652 28138 22704
rect 28902 22652 28908 22704
rect 28960 22692 28966 22704
rect 31113 22695 31171 22701
rect 31113 22692 31125 22695
rect 28960 22664 31125 22692
rect 28960 22652 28966 22664
rect 31113 22661 31125 22664
rect 31159 22661 31171 22695
rect 32320 22692 33120 22706
rect 31113 22655 31171 22661
rect 32232 22664 33120 22692
rect 28920 22624 28948 22652
rect 27908 22596 28948 22624
rect 30006 22584 30012 22636
rect 30064 22624 30070 22636
rect 30101 22627 30159 22633
rect 30101 22624 30113 22627
rect 30064 22596 30113 22624
rect 30064 22584 30070 22596
rect 30101 22593 30113 22596
rect 30147 22593 30159 22627
rect 30374 22624 30380 22636
rect 30335 22596 30380 22624
rect 30101 22587 30159 22593
rect 30374 22584 30380 22596
rect 30432 22584 30438 22636
rect 30558 22624 30564 22636
rect 30519 22596 30564 22624
rect 30558 22584 30564 22596
rect 30616 22584 30622 22636
rect 17696 22528 18719 22556
rect 17221 22519 17279 22525
rect 14148 22460 17172 22488
rect 17236 22488 17264 22519
rect 18691 22488 18719 22528
rect 19334 22516 19340 22568
rect 19392 22556 19398 22568
rect 19536 22556 19564 22584
rect 19702 22556 19708 22568
rect 19392 22528 19564 22556
rect 19615 22528 19708 22556
rect 19392 22516 19398 22528
rect 19702 22516 19708 22528
rect 19760 22556 19766 22568
rect 20530 22556 20536 22568
rect 19760 22528 20536 22556
rect 19760 22516 19766 22528
rect 20530 22516 20536 22528
rect 20588 22516 20594 22568
rect 21177 22559 21235 22565
rect 21177 22525 21189 22559
rect 21223 22525 21235 22559
rect 32232 22556 32260 22664
rect 32320 22650 33120 22664
rect 32232 22528 32352 22556
rect 21177 22519 21235 22525
rect 17236 22460 18184 22488
rect 18691 22460 19656 22488
rect 14148 22448 14154 22460
rect 15102 22420 15108 22432
rect 12820 22392 15108 22420
rect 15102 22380 15108 22392
rect 15160 22420 15166 22432
rect 15286 22420 15292 22432
rect 15160 22392 15292 22420
rect 15160 22380 15166 22392
rect 15286 22380 15292 22392
rect 15344 22380 15350 22432
rect 15562 22380 15568 22432
rect 15620 22420 15626 22432
rect 17126 22420 17132 22432
rect 15620 22392 17132 22420
rect 15620 22380 15626 22392
rect 17126 22380 17132 22392
rect 17184 22380 17190 22432
rect 17402 22380 17408 22432
rect 17460 22420 17466 22432
rect 18046 22420 18052 22432
rect 17460 22392 18052 22420
rect 17460 22380 17466 22392
rect 18046 22380 18052 22392
rect 18104 22380 18110 22432
rect 18156 22420 18184 22460
rect 19628 22432 19656 22460
rect 18690 22420 18696 22432
rect 18156 22392 18696 22420
rect 18690 22380 18696 22392
rect 18748 22380 18754 22432
rect 18874 22380 18880 22432
rect 18932 22420 18938 22432
rect 19518 22420 19524 22432
rect 18932 22392 19524 22420
rect 18932 22380 18938 22392
rect 19518 22380 19524 22392
rect 19576 22380 19582 22432
rect 19610 22380 19616 22432
rect 19668 22420 19674 22432
rect 21085 22423 21143 22429
rect 21085 22420 21097 22423
rect 19668 22392 21097 22420
rect 19668 22380 19674 22392
rect 21085 22389 21097 22392
rect 21131 22389 21143 22423
rect 21192 22420 21220 22519
rect 23293 22423 23351 22429
rect 23293 22420 23305 22423
rect 21192 22392 23305 22420
rect 21085 22383 21143 22389
rect 23293 22389 23305 22392
rect 23339 22420 23351 22423
rect 23750 22420 23756 22432
rect 23339 22392 23756 22420
rect 23339 22389 23351 22392
rect 23293 22383 23351 22389
rect 23750 22380 23756 22392
rect 23808 22380 23814 22432
rect 25590 22420 25596 22432
rect 25551 22392 25596 22420
rect 25590 22380 25596 22392
rect 25648 22380 25654 22432
rect 30650 22380 30656 22432
rect 30708 22420 30714 22432
rect 31205 22423 31263 22429
rect 31205 22420 31217 22423
rect 30708 22392 31217 22420
rect 30708 22380 30714 22392
rect 31205 22389 31217 22392
rect 31251 22389 31263 22423
rect 31205 22383 31263 22389
rect 1104 22330 32016 22352
rect 1104 22278 2136 22330
rect 2188 22278 12440 22330
rect 12492 22278 22744 22330
rect 22796 22278 32016 22330
rect 1104 22256 32016 22278
rect 1670 22176 1676 22228
rect 1728 22216 1734 22228
rect 1949 22219 2007 22225
rect 1949 22216 1961 22219
rect 1728 22188 1961 22216
rect 1728 22176 1734 22188
rect 1949 22185 1961 22188
rect 1995 22185 2007 22219
rect 3786 22216 3792 22228
rect 3747 22188 3792 22216
rect 1949 22179 2007 22185
rect 3786 22176 3792 22188
rect 3844 22176 3850 22228
rect 3878 22176 3884 22228
rect 3936 22216 3942 22228
rect 3936 22188 5672 22216
rect 3936 22176 3942 22188
rect 4890 22148 4896 22160
rect 4851 22120 4896 22148
rect 4890 22108 4896 22120
rect 4948 22108 4954 22160
rect 5258 22108 5264 22160
rect 5316 22148 5322 22160
rect 5644 22148 5672 22188
rect 5718 22176 5724 22228
rect 5776 22216 5782 22228
rect 5905 22219 5963 22225
rect 5905 22216 5917 22219
rect 5776 22188 5917 22216
rect 5776 22176 5782 22188
rect 5905 22185 5917 22188
rect 5951 22185 5963 22219
rect 5905 22179 5963 22185
rect 7469 22219 7527 22225
rect 7469 22185 7481 22219
rect 7515 22216 7527 22219
rect 7926 22216 7932 22228
rect 7515 22188 7932 22216
rect 7515 22185 7527 22188
rect 7469 22179 7527 22185
rect 7926 22176 7932 22188
rect 7984 22216 7990 22228
rect 8205 22219 8263 22225
rect 8205 22216 8217 22219
rect 7984 22188 8217 22216
rect 7984 22176 7990 22188
rect 8205 22185 8217 22188
rect 8251 22216 8263 22219
rect 9674 22216 9680 22228
rect 8251 22188 9680 22216
rect 8251 22185 8263 22188
rect 8205 22179 8263 22185
rect 9674 22176 9680 22188
rect 9732 22176 9738 22228
rect 9766 22176 9772 22228
rect 9824 22216 9830 22228
rect 12158 22216 12164 22228
rect 9824 22188 11928 22216
rect 12119 22188 12164 22216
rect 9824 22176 9830 22188
rect 9398 22148 9404 22160
rect 5316 22120 5488 22148
rect 5644 22120 9404 22148
rect 5316 22108 5322 22120
rect 5166 22080 5172 22092
rect 3896 22052 5172 22080
rect 1854 21972 1860 22024
rect 1912 22012 1918 22024
rect 2133 22015 2191 22021
rect 2133 22012 2145 22015
rect 1912 21984 2145 22012
rect 1912 21972 1918 21984
rect 2133 21981 2145 21984
rect 2179 22012 2191 22015
rect 2222 22012 2228 22024
rect 2179 21984 2228 22012
rect 2179 21981 2191 21984
rect 2133 21975 2191 21981
rect 2222 21972 2228 21984
rect 2280 21972 2286 22024
rect 2409 22015 2467 22021
rect 2409 21981 2421 22015
rect 2455 21981 2467 22015
rect 2409 21975 2467 21981
rect 2593 22015 2651 22021
rect 2593 21981 2605 22015
rect 2639 22012 2651 22015
rect 2682 22012 2688 22024
rect 2639 21984 2688 22012
rect 2639 21981 2651 21984
rect 2593 21975 2651 21981
rect 2424 21944 2452 21975
rect 2682 21972 2688 21984
rect 2740 21972 2746 22024
rect 3237 22015 3295 22021
rect 3237 21981 3249 22015
rect 3283 22012 3295 22015
rect 3786 22012 3792 22024
rect 3283 21984 3792 22012
rect 3283 21981 3295 21984
rect 3237 21975 3295 21981
rect 3786 21972 3792 21984
rect 3844 21972 3850 22024
rect 3896 21944 3924 22052
rect 4264 22021 4292 22052
rect 5166 22040 5172 22052
rect 5224 22080 5230 22092
rect 5460 22080 5488 22120
rect 9398 22108 9404 22120
rect 9456 22108 9462 22160
rect 11793 22151 11851 22157
rect 11793 22148 11805 22151
rect 10704 22120 11805 22148
rect 6273 22083 6331 22089
rect 6273 22080 6285 22083
rect 5224 22052 5396 22080
rect 5460 22052 6285 22080
rect 5224 22040 5230 22052
rect 3973 22015 4031 22021
rect 3973 21981 3985 22015
rect 4019 21981 4031 22015
rect 3973 21975 4031 21981
rect 4249 22015 4307 22021
rect 4249 21981 4261 22015
rect 4295 21981 4307 22015
rect 4430 22012 4436 22024
rect 4391 21984 4436 22012
rect 4249 21975 4307 21981
rect 2424 21916 3924 21944
rect 3988 21944 4016 21975
rect 4430 21972 4436 21984
rect 4488 21972 4494 22024
rect 4706 21972 4712 22024
rect 4764 22012 4770 22024
rect 5074 22012 5080 22024
rect 4764 21984 5080 22012
rect 4764 21972 4770 21984
rect 5074 21972 5080 21984
rect 5132 21972 5138 22024
rect 5368 22021 5396 22052
rect 6273 22049 6285 22052
rect 6319 22049 6331 22083
rect 7469 22083 7527 22089
rect 7469 22080 7481 22083
rect 6273 22043 6331 22049
rect 7116 22052 7481 22080
rect 5353 22015 5411 22021
rect 5353 21981 5365 22015
rect 5399 21981 5411 22015
rect 5353 21975 5411 21981
rect 5537 22015 5595 22021
rect 5537 21981 5549 22015
rect 5583 22012 5595 22015
rect 5718 22012 5724 22024
rect 5583 21984 5724 22012
rect 5583 21981 5595 21984
rect 5537 21975 5595 21981
rect 5718 21972 5724 21984
rect 5776 21972 5782 22024
rect 7116 22021 7144 22052
rect 7469 22049 7481 22052
rect 7515 22049 7527 22083
rect 7469 22043 7527 22049
rect 9030 22040 9036 22092
rect 9088 22080 9094 22092
rect 9088 22052 9536 22080
rect 9088 22040 9094 22052
rect 7101 22015 7159 22021
rect 6104 21984 7052 22012
rect 4724 21944 4752 21972
rect 6104 21953 6132 21984
rect 3988 21916 4752 21944
rect 5905 21947 5963 21953
rect 5905 21913 5917 21947
rect 5951 21944 5963 21947
rect 6089 21947 6147 21953
rect 6089 21944 6101 21947
rect 5951 21916 6101 21944
rect 5951 21913 5963 21916
rect 5905 21907 5963 21913
rect 6089 21913 6101 21916
rect 6135 21913 6147 21947
rect 6914 21944 6920 21956
rect 6875 21916 6920 21944
rect 6089 21907 6147 21913
rect 6914 21904 6920 21916
rect 6972 21904 6978 21956
rect 7024 21944 7052 21984
rect 7101 21981 7113 22015
rect 7147 21981 7159 22015
rect 7101 21975 7159 21981
rect 7377 22015 7435 22021
rect 7377 21981 7389 22015
rect 7423 22012 7435 22015
rect 7742 22012 7748 22024
rect 7423 21984 7748 22012
rect 7423 21981 7435 21984
rect 7377 21975 7435 21981
rect 7742 21972 7748 21984
rect 7800 21972 7806 22024
rect 7837 22015 7895 22021
rect 7837 21981 7849 22015
rect 7883 22012 7895 22015
rect 8018 22012 8024 22024
rect 7883 21984 8024 22012
rect 7883 21981 7895 21984
rect 7837 21975 7895 21981
rect 8018 21972 8024 21984
rect 8076 21972 8082 22024
rect 8294 22012 8300 22024
rect 8128 21984 8300 22012
rect 8128 21944 8156 21984
rect 8294 21972 8300 21984
rect 8352 21972 8358 22024
rect 8938 21972 8944 22024
rect 8996 22012 9002 22024
rect 9401 22015 9459 22021
rect 9401 22012 9413 22015
rect 8996 21984 9413 22012
rect 8996 21972 9002 21984
rect 9401 21981 9413 21984
rect 9447 21981 9459 22015
rect 9508 22012 9536 22052
rect 10704 22012 10732 22120
rect 11793 22117 11805 22120
rect 11839 22117 11851 22151
rect 11900 22148 11928 22188
rect 12158 22176 12164 22188
rect 12216 22176 12222 22228
rect 12268 22188 15516 22216
rect 12268 22148 12296 22188
rect 12710 22148 12716 22160
rect 11900 22120 12296 22148
rect 12360 22120 12716 22148
rect 11793 22111 11851 22117
rect 11238 22040 11244 22092
rect 11296 22080 11302 22092
rect 11701 22083 11759 22089
rect 11701 22080 11713 22083
rect 11296 22052 11713 22080
rect 11296 22040 11302 22052
rect 11701 22049 11713 22052
rect 11747 22049 11759 22083
rect 11701 22043 11759 22049
rect 12158 22040 12164 22092
rect 12216 22080 12222 22092
rect 12360 22080 12388 22120
rect 12710 22108 12716 22120
rect 12768 22108 12774 22160
rect 13357 22151 13415 22157
rect 13357 22117 13369 22151
rect 13403 22148 13415 22151
rect 13630 22148 13636 22160
rect 13403 22120 13636 22148
rect 13403 22117 13415 22120
rect 13357 22111 13415 22117
rect 13630 22108 13636 22120
rect 13688 22148 13694 22160
rect 14366 22148 14372 22160
rect 13688 22120 14372 22148
rect 13688 22108 13694 22120
rect 14366 22108 14372 22120
rect 14424 22108 14430 22160
rect 14918 22108 14924 22160
rect 14976 22148 14982 22160
rect 15286 22148 15292 22160
rect 14976 22120 15292 22148
rect 14976 22108 14982 22120
rect 15286 22108 15292 22120
rect 15344 22108 15350 22160
rect 15488 22148 15516 22188
rect 15562 22176 15568 22228
rect 15620 22216 15626 22228
rect 15657 22219 15715 22225
rect 15657 22216 15669 22219
rect 15620 22188 15669 22216
rect 15620 22176 15626 22188
rect 15657 22185 15669 22188
rect 15703 22185 15715 22219
rect 15657 22179 15715 22185
rect 15930 22176 15936 22228
rect 15988 22216 15994 22228
rect 17402 22216 17408 22228
rect 15988 22188 17408 22216
rect 15988 22176 15994 22188
rect 17402 22176 17408 22188
rect 17460 22176 17466 22228
rect 17788 22188 19380 22216
rect 17788 22148 17816 22188
rect 15488 22120 17816 22148
rect 18230 22108 18236 22160
rect 18288 22148 18294 22160
rect 19245 22151 19303 22157
rect 19245 22148 19257 22151
rect 18288 22120 19257 22148
rect 18288 22108 18294 22120
rect 19245 22117 19257 22120
rect 19291 22117 19303 22151
rect 19352 22148 19380 22188
rect 19426 22176 19432 22228
rect 19484 22216 19490 22228
rect 20257 22219 20315 22225
rect 20257 22216 20269 22219
rect 19484 22188 20269 22216
rect 19484 22176 19490 22188
rect 20257 22185 20269 22188
rect 20303 22185 20315 22219
rect 32324 22216 32352 22528
rect 20257 22179 20315 22185
rect 22066 22188 32352 22216
rect 22066 22148 22094 22188
rect 19352 22120 22094 22148
rect 19245 22111 19303 22117
rect 22554 22108 22560 22160
rect 22612 22148 22618 22160
rect 23109 22151 23167 22157
rect 23109 22148 23121 22151
rect 22612 22120 23121 22148
rect 22612 22108 22618 22120
rect 23109 22117 23121 22120
rect 23155 22117 23167 22151
rect 23109 22111 23167 22117
rect 26973 22151 27031 22157
rect 26973 22117 26985 22151
rect 27019 22148 27031 22151
rect 27246 22148 27252 22160
rect 27019 22120 27252 22148
rect 27019 22117 27031 22120
rect 26973 22111 27031 22117
rect 27246 22108 27252 22120
rect 27304 22108 27310 22160
rect 12526 22080 12532 22092
rect 12216 22052 12388 22080
rect 12487 22052 12532 22080
rect 12216 22040 12222 22052
rect 12526 22040 12532 22052
rect 12584 22040 12590 22092
rect 12621 22083 12679 22089
rect 12621 22049 12633 22083
rect 12667 22080 12679 22083
rect 12894 22080 12900 22092
rect 12667 22052 12900 22080
rect 12667 22049 12679 22052
rect 12621 22043 12679 22049
rect 12894 22040 12900 22052
rect 12952 22040 12958 22092
rect 13004 22052 13308 22080
rect 9508 21984 10732 22012
rect 9401 21975 9459 21981
rect 10870 21972 10876 22024
rect 10928 22012 10934 22024
rect 11425 22015 11483 22021
rect 11425 22012 11437 22015
rect 10928 21984 11437 22012
rect 10928 21972 10934 21984
rect 11425 21981 11437 21984
rect 11471 21981 11483 22015
rect 11609 22015 11667 22021
rect 11609 22012 11621 22015
rect 11425 21975 11483 21981
rect 11532 21984 11621 22012
rect 9668 21947 9726 21953
rect 7024 21916 8156 21944
rect 8220 21916 9628 21944
rect 3053 21879 3111 21885
rect 3053 21845 3065 21879
rect 3099 21876 3111 21879
rect 3142 21876 3148 21888
rect 3099 21848 3148 21876
rect 3099 21845 3111 21848
rect 3053 21839 3111 21845
rect 3142 21836 3148 21848
rect 3200 21836 3206 21888
rect 4246 21836 4252 21888
rect 4304 21876 4310 21888
rect 6270 21876 6276 21888
rect 4304 21848 6276 21876
rect 4304 21836 4310 21848
rect 6270 21836 6276 21848
rect 6328 21836 6334 21888
rect 7285 21879 7343 21885
rect 7285 21845 7297 21879
rect 7331 21876 7343 21879
rect 7466 21876 7472 21888
rect 7331 21848 7472 21876
rect 7331 21845 7343 21848
rect 7285 21839 7343 21845
rect 7466 21836 7472 21848
rect 7524 21836 7530 21888
rect 7926 21836 7932 21888
rect 7984 21876 7990 21888
rect 8220 21885 8248 21916
rect 8205 21879 8263 21885
rect 8205 21876 8217 21879
rect 7984 21848 8217 21876
rect 7984 21836 7990 21848
rect 8205 21845 8217 21848
rect 8251 21845 8263 21879
rect 8386 21876 8392 21888
rect 8347 21848 8392 21876
rect 8205 21839 8263 21845
rect 8386 21836 8392 21848
rect 8444 21836 8450 21888
rect 9600 21876 9628 21916
rect 9668 21913 9680 21947
rect 9714 21944 9726 21947
rect 11241 21947 11299 21953
rect 11241 21944 11253 21947
rect 9714 21916 11253 21944
rect 9714 21913 9726 21916
rect 9668 21907 9726 21913
rect 11241 21913 11253 21916
rect 11287 21913 11299 21947
rect 11241 21907 11299 21913
rect 10502 21876 10508 21888
rect 9600 21848 10508 21876
rect 10502 21836 10508 21848
rect 10560 21836 10566 21888
rect 10778 21876 10784 21888
rect 10739 21848 10784 21876
rect 10778 21836 10784 21848
rect 10836 21836 10842 21888
rect 10962 21836 10968 21888
rect 11020 21876 11026 21888
rect 11532 21876 11560 21984
rect 11609 21981 11621 21984
rect 11655 21981 11667 22015
rect 12342 22012 12348 22024
rect 12303 21984 12348 22012
rect 11609 21975 11667 21981
rect 12342 21972 12348 21984
rect 12400 21972 12406 22024
rect 13004 22012 13032 22052
rect 12452 21984 13032 22012
rect 12452 21944 12480 21984
rect 13078 21972 13084 22024
rect 13136 22012 13142 22024
rect 13173 22015 13231 22021
rect 13173 22012 13185 22015
rect 13136 21984 13185 22012
rect 13136 21972 13142 21984
rect 13173 21981 13185 21984
rect 13219 21981 13231 22015
rect 13280 22012 13308 22052
rect 13446 22040 13452 22092
rect 13504 22080 13510 22092
rect 15657 22083 15715 22089
rect 15657 22080 15669 22083
rect 13504 22052 15669 22080
rect 13504 22040 13510 22052
rect 15657 22049 15669 22052
rect 15703 22049 15715 22083
rect 15657 22043 15715 22049
rect 16114 22040 16120 22092
rect 16172 22080 16178 22092
rect 17402 22080 17408 22092
rect 16172 22052 17408 22080
rect 16172 22040 16178 22052
rect 17402 22040 17408 22052
rect 17460 22040 17466 22092
rect 18874 22080 18880 22092
rect 17984 22052 18880 22080
rect 14093 22015 14151 22021
rect 13280 21984 14044 22012
rect 13173 21975 13231 21981
rect 11624 21916 12480 21944
rect 11624 21888 11652 21916
rect 12526 21904 12532 21956
rect 12584 21944 12590 21956
rect 13814 21944 13820 21956
rect 12584 21916 13820 21944
rect 12584 21904 12590 21916
rect 13814 21904 13820 21916
rect 13872 21904 13878 21956
rect 14016 21944 14044 21984
rect 14093 21981 14105 22015
rect 14139 22012 14151 22015
rect 14550 22012 14556 22024
rect 14139 21984 14556 22012
rect 14139 21981 14151 21984
rect 14093 21975 14151 21981
rect 14550 21972 14556 21984
rect 14608 21972 14614 22024
rect 15102 22012 15108 22024
rect 15063 21984 15108 22012
rect 15102 21972 15108 21984
rect 15160 21972 15166 22024
rect 15381 22015 15439 22021
rect 15381 21981 15393 22015
rect 15427 22012 15439 22015
rect 15470 22012 15476 22024
rect 15427 21984 15476 22012
rect 15427 21981 15439 21984
rect 15381 21975 15439 21981
rect 15470 21972 15476 21984
rect 15528 21972 15534 22024
rect 15562 21972 15568 22024
rect 15620 22012 15626 22024
rect 16224 22012 16436 22014
rect 15620 21984 15665 22012
rect 16132 21986 16436 22012
rect 16132 21984 16252 21986
rect 15620 21972 15626 21984
rect 16132 21956 16160 21984
rect 14642 21944 14648 21956
rect 14016 21916 14648 21944
rect 14642 21904 14648 21916
rect 14700 21904 14706 21956
rect 15286 21904 15292 21956
rect 15344 21944 15350 21956
rect 16025 21947 16083 21953
rect 16025 21944 16037 21947
rect 15344 21916 16037 21944
rect 15344 21904 15350 21916
rect 16025 21913 16037 21916
rect 16071 21913 16083 21947
rect 16025 21907 16083 21913
rect 16114 21904 16120 21956
rect 16172 21904 16178 21956
rect 16408 21953 16436 21986
rect 17126 21972 17132 22024
rect 17184 22012 17190 22024
rect 17984 22012 18012 22052
rect 18874 22040 18880 22052
rect 18932 22040 18938 22092
rect 19610 22080 19616 22092
rect 19571 22052 19616 22080
rect 19610 22040 19616 22052
rect 19668 22040 19674 22092
rect 19705 22083 19763 22089
rect 19705 22049 19717 22083
rect 19751 22080 19763 22083
rect 20990 22080 20996 22092
rect 19751 22052 20996 22080
rect 19751 22049 19763 22052
rect 19705 22043 19763 22049
rect 20990 22040 20996 22052
rect 21048 22080 21054 22092
rect 21361 22083 21419 22089
rect 21361 22080 21373 22083
rect 21048 22052 21373 22080
rect 21048 22040 21054 22052
rect 21361 22049 21373 22052
rect 21407 22049 21419 22083
rect 22922 22080 22928 22092
rect 21361 22043 21419 22049
rect 22204 22052 22928 22080
rect 17184 21984 18012 22012
rect 17184 21972 17190 21984
rect 18046 21972 18052 22024
rect 18104 22012 18110 22024
rect 19429 22015 19487 22021
rect 19429 22012 19441 22015
rect 18104 21984 19441 22012
rect 18104 21972 18110 21984
rect 19429 21981 19441 21984
rect 19475 21981 19487 22015
rect 19429 21975 19487 21981
rect 19794 21972 19800 22024
rect 19852 22012 19858 22024
rect 20165 22015 20223 22021
rect 20165 22012 20177 22015
rect 19852 21984 20177 22012
rect 19852 21972 19858 21984
rect 20165 21981 20177 21984
rect 20211 21981 20223 22015
rect 20165 21975 20223 21981
rect 20349 22015 20407 22021
rect 20349 21981 20361 22015
rect 20395 21981 20407 22015
rect 20349 21975 20407 21981
rect 16301 21947 16359 21953
rect 16301 21913 16313 21947
rect 16347 21913 16359 21947
rect 16301 21907 16359 21913
rect 16395 21947 16453 21953
rect 16395 21913 16407 21947
rect 16441 21913 16453 21947
rect 17957 21947 18015 21953
rect 17957 21944 17969 21947
rect 16395 21907 16453 21913
rect 16546 21916 17969 21944
rect 11020 21848 11560 21876
rect 11020 21836 11026 21848
rect 11606 21836 11612 21888
rect 11664 21836 11670 21888
rect 11793 21879 11851 21885
rect 11793 21845 11805 21879
rect 11839 21876 11851 21879
rect 14277 21879 14335 21885
rect 14277 21876 14289 21879
rect 11839 21848 14289 21876
rect 11839 21845 11851 21848
rect 11793 21839 11851 21845
rect 14277 21845 14289 21848
rect 14323 21845 14335 21879
rect 14277 21839 14335 21845
rect 14366 21836 14372 21888
rect 14424 21876 14430 21888
rect 14921 21879 14979 21885
rect 14921 21876 14933 21879
rect 14424 21848 14933 21876
rect 14424 21836 14430 21848
rect 14921 21845 14933 21848
rect 14967 21845 14979 21879
rect 14921 21839 14979 21845
rect 15470 21836 15476 21888
rect 15528 21876 15534 21888
rect 15657 21879 15715 21885
rect 15657 21876 15669 21879
rect 15528 21848 15669 21876
rect 15528 21836 15534 21848
rect 15657 21845 15669 21848
rect 15703 21845 15715 21879
rect 16316 21876 16344 21907
rect 16546 21876 16574 21916
rect 17957 21913 17969 21916
rect 18003 21913 18015 21947
rect 17957 21907 18015 21913
rect 18322 21904 18328 21956
rect 18380 21944 18386 21956
rect 20364 21944 20392 21975
rect 20898 21972 20904 22024
rect 20956 22012 20962 22024
rect 22005 22015 22063 22021
rect 22005 22012 22017 22015
rect 20956 21984 22017 22012
rect 20956 21972 20962 21984
rect 22005 21981 22017 21984
rect 22051 21981 22063 22015
rect 22005 21975 22063 21981
rect 22094 21972 22100 22024
rect 22152 22012 22158 22024
rect 22204 22021 22232 22052
rect 22922 22040 22928 22052
rect 22980 22040 22986 22092
rect 27706 22080 27712 22092
rect 23768 22052 24808 22080
rect 27619 22052 27712 22080
rect 23768 22024 23796 22052
rect 22189 22015 22247 22021
rect 22189 22012 22201 22015
rect 22152 21984 22201 22012
rect 22152 21972 22158 21984
rect 22189 21981 22201 21984
rect 22235 21981 22247 22015
rect 22189 21975 22247 21981
rect 22370 21972 22376 22024
rect 22428 22012 22434 22024
rect 22465 22015 22523 22021
rect 22465 22012 22477 22015
rect 22428 21984 22477 22012
rect 22428 21972 22434 21984
rect 22465 21981 22477 21984
rect 22511 21981 22523 22015
rect 22465 21975 22523 21981
rect 22649 22015 22707 22021
rect 22649 21981 22661 22015
rect 22695 21981 22707 22015
rect 22649 21975 22707 21981
rect 23293 22015 23351 22021
rect 23293 21981 23305 22015
rect 23339 21981 23351 22015
rect 23293 21975 23351 21981
rect 18380 21916 20392 21944
rect 18380 21904 18386 21916
rect 21910 21904 21916 21956
rect 21968 21944 21974 21956
rect 22480 21944 22508 21975
rect 21968 21916 22508 21944
rect 21968 21904 21974 21916
rect 16316 21848 16574 21876
rect 15657 21839 15715 21845
rect 17678 21836 17684 21888
rect 17736 21876 17742 21888
rect 18782 21876 18788 21888
rect 17736 21848 18788 21876
rect 17736 21836 17742 21848
rect 18782 21836 18788 21848
rect 18840 21836 18846 21888
rect 19150 21836 19156 21888
rect 19208 21876 19214 21888
rect 20162 21876 20168 21888
rect 19208 21848 20168 21876
rect 19208 21836 19214 21848
rect 20162 21836 20168 21848
rect 20220 21836 20226 21888
rect 20809 21879 20867 21885
rect 20809 21845 20821 21879
rect 20855 21876 20867 21879
rect 20898 21876 20904 21888
rect 20855 21848 20904 21876
rect 20855 21845 20867 21848
rect 20809 21839 20867 21845
rect 20898 21836 20904 21848
rect 20956 21836 20962 21888
rect 21174 21876 21180 21888
rect 21135 21848 21180 21876
rect 21174 21836 21180 21848
rect 21232 21836 21238 21888
rect 21269 21879 21327 21885
rect 21269 21845 21281 21879
rect 21315 21876 21327 21879
rect 22370 21876 22376 21888
rect 21315 21848 22376 21876
rect 21315 21845 21327 21848
rect 21269 21839 21327 21845
rect 22370 21836 22376 21848
rect 22428 21836 22434 21888
rect 22462 21836 22468 21888
rect 22520 21876 22526 21888
rect 22664 21876 22692 21975
rect 22922 21904 22928 21956
rect 22980 21944 22986 21956
rect 23308 21944 23336 21975
rect 23382 21972 23388 22024
rect 23440 22012 23446 22024
rect 23569 22015 23627 22021
rect 23569 22012 23581 22015
rect 23440 21984 23581 22012
rect 23440 21972 23446 21984
rect 23569 21981 23581 21984
rect 23615 21981 23627 22015
rect 23750 22012 23756 22024
rect 23711 21984 23756 22012
rect 23569 21975 23627 21981
rect 23750 21972 23756 21984
rect 23808 21972 23814 22024
rect 24578 22012 24584 22024
rect 24539 21984 24584 22012
rect 24578 21972 24584 21984
rect 24636 21972 24642 22024
rect 24780 22021 24808 22052
rect 27706 22040 27712 22052
rect 27764 22080 27770 22092
rect 28442 22080 28448 22092
rect 27764 22052 28448 22080
rect 27764 22040 27770 22052
rect 28442 22040 28448 22052
rect 28500 22040 28506 22092
rect 24765 22015 24823 22021
rect 24765 21981 24777 22015
rect 24811 21981 24823 22015
rect 24765 21975 24823 21981
rect 24854 21972 24860 22024
rect 24912 22012 24918 22024
rect 25593 22015 25651 22021
rect 24912 21984 24957 22012
rect 24912 21972 24918 21984
rect 25593 21981 25605 22015
rect 25639 22012 25651 22015
rect 25682 22012 25688 22024
rect 25639 21984 25688 22012
rect 25639 21981 25651 21984
rect 25593 21975 25651 21981
rect 25682 21972 25688 21984
rect 25740 21972 25746 22024
rect 26786 21972 26792 22024
rect 26844 22012 26850 22024
rect 27433 22015 27491 22021
rect 27433 22012 27445 22015
rect 26844 21984 27445 22012
rect 26844 21972 26850 21984
rect 27433 21981 27445 21984
rect 27479 22012 27491 22015
rect 28813 22015 28871 22021
rect 28813 22012 28825 22015
rect 27479 21984 28825 22012
rect 27479 21981 27491 21984
rect 27433 21975 27491 21981
rect 28813 21981 28825 21984
rect 28859 22012 28871 22015
rect 29270 22012 29276 22024
rect 28859 21984 29276 22012
rect 28859 21981 28871 21984
rect 28813 21975 28871 21981
rect 29270 21972 29276 21984
rect 29328 21972 29334 22024
rect 29914 22012 29920 22024
rect 29875 21984 29920 22012
rect 29914 21972 29920 21984
rect 29972 21972 29978 22024
rect 30926 22012 30932 22024
rect 30024 21984 30932 22012
rect 22980 21916 23336 21944
rect 25860 21947 25918 21953
rect 22980 21904 22986 21916
rect 25860 21913 25872 21947
rect 25906 21944 25918 21947
rect 25958 21944 25964 21956
rect 25906 21916 25964 21944
rect 25906 21913 25918 21916
rect 25860 21907 25918 21913
rect 25958 21904 25964 21916
rect 26016 21904 26022 21956
rect 28997 21947 29055 21953
rect 28997 21913 29009 21947
rect 29043 21944 29055 21947
rect 30024 21944 30052 21984
rect 30926 21972 30932 21984
rect 30984 21972 30990 22024
rect 29043 21916 30052 21944
rect 30184 21947 30242 21953
rect 29043 21913 29055 21916
rect 28997 21907 29055 21913
rect 30184 21913 30196 21947
rect 30230 21944 30242 21947
rect 30742 21944 30748 21956
rect 30230 21916 30748 21944
rect 30230 21913 30242 21916
rect 30184 21907 30242 21913
rect 30742 21904 30748 21916
rect 30800 21904 30806 21956
rect 22520 21848 22692 21876
rect 24397 21879 24455 21885
rect 22520 21836 22526 21848
rect 24397 21845 24409 21879
rect 24443 21876 24455 21879
rect 24946 21876 24952 21888
rect 24443 21848 24952 21876
rect 24443 21845 24455 21848
rect 24397 21839 24455 21845
rect 24946 21836 24952 21848
rect 25004 21836 25010 21888
rect 30558 21836 30564 21888
rect 30616 21876 30622 21888
rect 31297 21879 31355 21885
rect 31297 21876 31309 21879
rect 30616 21848 31309 21876
rect 30616 21836 30622 21848
rect 31297 21845 31309 21848
rect 31343 21845 31355 21879
rect 31297 21839 31355 21845
rect 1104 21786 32016 21808
rect 1104 21734 7288 21786
rect 7340 21734 17592 21786
rect 17644 21734 27896 21786
rect 27948 21734 32016 21786
rect 1104 21712 32016 21734
rect 1394 21632 1400 21684
rect 1452 21672 1458 21684
rect 2314 21672 2320 21684
rect 1452 21644 2320 21672
rect 1452 21632 1458 21644
rect 2314 21632 2320 21644
rect 2372 21632 2378 21684
rect 5074 21632 5080 21684
rect 5132 21672 5138 21684
rect 5629 21675 5687 21681
rect 5629 21672 5641 21675
rect 5132 21644 5641 21672
rect 5132 21632 5138 21644
rect 5629 21641 5641 21644
rect 5675 21641 5687 21675
rect 5629 21635 5687 21641
rect 6454 21632 6460 21684
rect 6512 21672 6518 21684
rect 7653 21675 7711 21681
rect 7653 21672 7665 21675
rect 6512 21644 7665 21672
rect 6512 21632 6518 21644
rect 7653 21641 7665 21644
rect 7699 21641 7711 21675
rect 7653 21635 7711 21641
rect 9861 21675 9919 21681
rect 9861 21641 9873 21675
rect 9907 21672 9919 21675
rect 10870 21672 10876 21684
rect 9907 21644 10876 21672
rect 9907 21641 9919 21644
rect 9861 21635 9919 21641
rect 10870 21632 10876 21644
rect 10928 21632 10934 21684
rect 11977 21675 12035 21681
rect 11977 21641 11989 21675
rect 12023 21672 12035 21675
rect 12023 21644 13400 21672
rect 12023 21641 12035 21644
rect 11977 21635 12035 21641
rect 3136 21607 3194 21613
rect 3136 21573 3148 21607
rect 3182 21604 3194 21607
rect 3602 21604 3608 21616
rect 3182 21576 3608 21604
rect 3182 21573 3194 21576
rect 3136 21567 3194 21573
rect 3602 21564 3608 21576
rect 3660 21564 3666 21616
rect 3786 21564 3792 21616
rect 3844 21604 3850 21616
rect 9401 21607 9459 21613
rect 3844 21576 9352 21604
rect 3844 21564 3850 21576
rect 1397 21539 1455 21545
rect 1397 21505 1409 21539
rect 1443 21505 1455 21539
rect 1397 21499 1455 21505
rect 2409 21539 2467 21545
rect 2409 21505 2421 21539
rect 2455 21536 2467 21539
rect 2498 21536 2504 21548
rect 2455 21508 2504 21536
rect 2455 21505 2467 21508
rect 2409 21499 2467 21505
rect 1412 21332 1440 21499
rect 2498 21496 2504 21508
rect 2556 21496 2562 21548
rect 4890 21536 4896 21548
rect 4851 21508 4896 21536
rect 4890 21496 4896 21508
rect 4948 21496 4954 21548
rect 5813 21539 5871 21545
rect 5813 21505 5825 21539
rect 5859 21536 5871 21539
rect 6454 21536 6460 21548
rect 5859 21508 6460 21536
rect 5859 21505 5871 21508
rect 5813 21499 5871 21505
rect 2774 21428 2780 21480
rect 2832 21468 2838 21480
rect 2869 21471 2927 21477
rect 2869 21468 2881 21471
rect 2832 21440 2881 21468
rect 2832 21428 2838 21440
rect 2869 21437 2881 21440
rect 2915 21437 2927 21471
rect 4430 21468 4436 21480
rect 2869 21431 2927 21437
rect 4264 21440 4436 21468
rect 4264 21409 4292 21440
rect 4430 21428 4436 21440
rect 4488 21468 4494 21480
rect 5169 21471 5227 21477
rect 5169 21468 5181 21471
rect 4488 21440 5181 21468
rect 4488 21428 4494 21440
rect 5169 21437 5181 21440
rect 5215 21468 5227 21471
rect 5258 21468 5264 21480
rect 5215 21440 5264 21468
rect 5215 21437 5227 21440
rect 5169 21431 5227 21437
rect 5258 21428 5264 21440
rect 5316 21428 5322 21480
rect 4249 21403 4307 21409
rect 4249 21369 4261 21403
rect 4295 21369 4307 21403
rect 5828 21400 5856 21499
rect 6454 21496 6460 21508
rect 6512 21536 6518 21548
rect 6549 21539 6607 21545
rect 6549 21536 6561 21539
rect 6512 21508 6561 21536
rect 6512 21496 6518 21508
rect 6549 21505 6561 21508
rect 6595 21505 6607 21539
rect 7834 21536 7840 21548
rect 7795 21508 7840 21536
rect 6549 21499 6607 21505
rect 7834 21496 7840 21508
rect 7892 21496 7898 21548
rect 8113 21539 8171 21545
rect 8113 21505 8125 21539
rect 8159 21536 8171 21539
rect 8386 21536 8392 21548
rect 8159 21508 8392 21536
rect 8159 21505 8171 21508
rect 8113 21499 8171 21505
rect 8386 21496 8392 21508
rect 8444 21496 8450 21548
rect 9214 21536 9220 21548
rect 9175 21508 9220 21536
rect 9214 21496 9220 21508
rect 9272 21496 9278 21548
rect 6914 21428 6920 21480
rect 6972 21468 6978 21480
rect 7929 21471 7987 21477
rect 7929 21468 7941 21471
rect 6972 21440 7941 21468
rect 6972 21428 6978 21440
rect 7929 21437 7941 21440
rect 7975 21437 7987 21471
rect 7929 21431 7987 21437
rect 8018 21428 8024 21480
rect 8076 21468 8082 21480
rect 9324 21468 9352 21576
rect 9401 21573 9413 21607
rect 9447 21604 9459 21607
rect 12805 21607 12863 21613
rect 12805 21604 12817 21607
rect 9447 21576 12817 21604
rect 9447 21573 9459 21576
rect 9401 21567 9459 21573
rect 12805 21573 12817 21576
rect 12851 21573 12863 21607
rect 13372 21604 13400 21644
rect 13814 21632 13820 21684
rect 13872 21672 13878 21684
rect 13872 21644 15976 21672
rect 13872 21632 13878 21644
rect 14642 21604 14648 21616
rect 13372 21576 14648 21604
rect 12805 21567 12863 21573
rect 14642 21564 14648 21576
rect 14700 21604 14706 21616
rect 15838 21604 15844 21616
rect 14700 21576 15844 21604
rect 14700 21564 14706 21576
rect 15838 21564 15844 21576
rect 15896 21564 15902 21616
rect 15948 21604 15976 21644
rect 16298 21632 16304 21684
rect 16356 21672 16362 21684
rect 20717 21675 20775 21681
rect 16356 21644 20668 21672
rect 16356 21632 16362 21644
rect 16666 21604 16672 21616
rect 15948 21576 16672 21604
rect 16666 21564 16672 21576
rect 16724 21564 16730 21616
rect 16758 21564 16764 21616
rect 16816 21604 16822 21616
rect 16914 21607 16972 21613
rect 16914 21604 16926 21607
rect 16816 21576 16926 21604
rect 16816 21564 16822 21576
rect 16914 21573 16926 21576
rect 16960 21573 16972 21607
rect 19150 21604 19156 21616
rect 16914 21567 16972 21573
rect 17026 21576 19156 21604
rect 9950 21496 9956 21548
rect 10008 21536 10014 21548
rect 10045 21539 10103 21545
rect 10045 21536 10057 21539
rect 10008 21508 10057 21536
rect 10008 21496 10014 21508
rect 10045 21505 10057 21508
rect 10091 21505 10103 21539
rect 10318 21536 10324 21548
rect 10279 21508 10324 21536
rect 10045 21499 10103 21505
rect 10318 21496 10324 21508
rect 10376 21496 10382 21548
rect 10505 21539 10563 21545
rect 10505 21505 10517 21539
rect 10551 21536 10563 21539
rect 10597 21539 10655 21545
rect 10597 21536 10609 21539
rect 10551 21508 10609 21536
rect 10551 21505 10563 21508
rect 10505 21499 10563 21505
rect 10597 21505 10609 21508
rect 10643 21536 10655 21539
rect 10778 21536 10784 21548
rect 10643 21508 10784 21536
rect 10643 21505 10655 21508
rect 10597 21499 10655 21505
rect 10778 21496 10784 21508
rect 10836 21496 10842 21548
rect 11238 21496 11244 21548
rect 11296 21536 11302 21548
rect 11698 21536 11704 21548
rect 11296 21508 11704 21536
rect 11296 21496 11302 21508
rect 11698 21496 11704 21508
rect 11756 21536 11762 21548
rect 12069 21539 12127 21545
rect 12069 21536 12081 21539
rect 11756 21508 12081 21536
rect 11756 21496 11762 21508
rect 12069 21505 12081 21508
rect 12115 21505 12127 21539
rect 12069 21499 12127 21505
rect 12158 21496 12164 21548
rect 12216 21536 12222 21548
rect 12253 21539 12311 21545
rect 12253 21536 12265 21539
rect 12216 21508 12265 21536
rect 12216 21496 12222 21508
rect 12253 21505 12265 21508
rect 12299 21505 12311 21539
rect 12253 21499 12311 21505
rect 12342 21496 12348 21548
rect 12400 21536 12406 21548
rect 12989 21539 13047 21545
rect 12989 21536 13001 21539
rect 12400 21508 13001 21536
rect 12400 21496 12406 21508
rect 12989 21505 13001 21508
rect 13035 21505 13047 21539
rect 12989 21499 13047 21505
rect 13173 21539 13231 21545
rect 13173 21505 13185 21539
rect 13219 21536 13231 21539
rect 13446 21536 13452 21548
rect 13219 21508 13452 21536
rect 13219 21505 13231 21508
rect 13173 21499 13231 21505
rect 13446 21496 13452 21508
rect 13504 21496 13510 21548
rect 14366 21536 14372 21548
rect 14327 21508 14372 21536
rect 14366 21496 14372 21508
rect 14424 21496 14430 21548
rect 14826 21496 14832 21548
rect 14884 21536 14890 21548
rect 15289 21539 15347 21545
rect 15289 21536 15301 21539
rect 14884 21508 15301 21536
rect 14884 21496 14890 21508
rect 15289 21505 15301 21508
rect 15335 21505 15347 21539
rect 15289 21499 15347 21505
rect 15565 21539 15623 21545
rect 15565 21505 15577 21539
rect 15611 21536 15623 21539
rect 15746 21536 15752 21548
rect 15611 21508 15752 21536
rect 15611 21505 15623 21508
rect 15565 21499 15623 21505
rect 15746 21496 15752 21508
rect 15804 21496 15810 21548
rect 17026 21536 17054 21576
rect 19150 21564 19156 21576
rect 19208 21564 19214 21616
rect 19334 21564 19340 21616
rect 19392 21564 19398 21616
rect 19604 21607 19662 21613
rect 19604 21573 19616 21607
rect 19650 21604 19662 21607
rect 20438 21604 20444 21616
rect 19650 21576 20444 21604
rect 19650 21573 19662 21576
rect 19604 21567 19662 21573
rect 20438 21564 20444 21576
rect 20496 21564 20502 21616
rect 20640 21604 20668 21644
rect 20717 21641 20729 21675
rect 20763 21672 20775 21675
rect 20990 21672 20996 21684
rect 20763 21644 20996 21672
rect 20763 21641 20775 21644
rect 20717 21635 20775 21641
rect 20990 21632 20996 21644
rect 21048 21632 21054 21684
rect 21913 21675 21971 21681
rect 21913 21641 21925 21675
rect 21959 21672 21971 21675
rect 22002 21672 22008 21684
rect 21959 21644 22008 21672
rect 21959 21641 21971 21644
rect 21913 21635 21971 21641
rect 22002 21632 22008 21644
rect 22060 21632 22066 21684
rect 22186 21632 22192 21684
rect 22244 21672 22250 21684
rect 22465 21675 22523 21681
rect 22465 21672 22477 21675
rect 22244 21644 22477 21672
rect 22244 21632 22250 21644
rect 22465 21641 22477 21644
rect 22511 21641 22523 21675
rect 22465 21635 22523 21641
rect 22741 21675 22799 21681
rect 22741 21641 22753 21675
rect 22787 21672 22799 21675
rect 22833 21675 22891 21681
rect 22833 21672 22845 21675
rect 22787 21644 22845 21672
rect 22787 21641 22799 21644
rect 22741 21635 22799 21641
rect 22833 21641 22845 21644
rect 22879 21641 22891 21675
rect 23198 21672 23204 21684
rect 23159 21644 23204 21672
rect 22833 21635 22891 21641
rect 23198 21632 23204 21644
rect 23256 21632 23262 21684
rect 24486 21632 24492 21684
rect 24544 21672 24550 21684
rect 24581 21675 24639 21681
rect 24581 21672 24593 21675
rect 24544 21644 24593 21672
rect 24544 21632 24550 21644
rect 24581 21641 24593 21644
rect 24627 21641 24639 21675
rect 25958 21672 25964 21684
rect 25919 21644 25964 21672
rect 24581 21635 24639 21641
rect 25958 21632 25964 21644
rect 26016 21632 26022 21684
rect 26418 21632 26424 21684
rect 26476 21672 26482 21684
rect 27338 21672 27344 21684
rect 26476 21644 27344 21672
rect 26476 21632 26482 21644
rect 27338 21632 27344 21644
rect 27396 21672 27402 21684
rect 31110 21672 31116 21684
rect 27396 21644 28948 21672
rect 27396 21632 27402 21644
rect 21818 21604 21824 21616
rect 20640 21576 21824 21604
rect 21818 21564 21824 21576
rect 21876 21564 21882 21616
rect 23293 21607 23351 21613
rect 23293 21604 23305 21607
rect 21928 21576 23305 21604
rect 15856 21508 17054 21536
rect 18141 21539 18199 21545
rect 11977 21471 12035 21477
rect 11977 21468 11989 21471
rect 8076 21440 8169 21468
rect 9324 21440 11989 21468
rect 8076 21428 8082 21440
rect 11977 21437 11989 21440
rect 12023 21437 12035 21471
rect 11977 21431 12035 21437
rect 12529 21471 12587 21477
rect 12529 21437 12541 21471
rect 12575 21468 12587 21471
rect 14274 21468 14280 21480
rect 12575 21440 14280 21468
rect 12575 21437 12587 21440
rect 12529 21431 12587 21437
rect 14274 21428 14280 21440
rect 14332 21428 14338 21480
rect 14645 21471 14703 21477
rect 14645 21437 14657 21471
rect 14691 21468 14703 21471
rect 14918 21468 14924 21480
rect 14691 21440 14924 21468
rect 14691 21437 14703 21440
rect 14645 21431 14703 21437
rect 14918 21428 14924 21440
rect 14976 21428 14982 21480
rect 15102 21428 15108 21480
rect 15160 21468 15166 21480
rect 15473 21471 15531 21477
rect 15160 21440 15205 21468
rect 15160 21428 15166 21440
rect 15473 21437 15485 21471
rect 15519 21468 15531 21471
rect 15654 21468 15660 21480
rect 15519 21440 15660 21468
rect 15519 21437 15531 21440
rect 15473 21431 15531 21437
rect 6730 21400 6736 21412
rect 4249 21363 4307 21369
rect 4356 21372 5856 21400
rect 6691 21372 6736 21400
rect 768 21304 1440 21332
rect 1581 21335 1639 21341
rect 768 21060 796 21304
rect 1581 21301 1593 21335
rect 1627 21332 1639 21335
rect 1670 21332 1676 21344
rect 1627 21304 1676 21332
rect 1627 21301 1639 21304
rect 1581 21295 1639 21301
rect 1670 21292 1676 21304
rect 1728 21292 1734 21344
rect 2225 21335 2283 21341
rect 2225 21301 2237 21335
rect 2271 21332 2283 21335
rect 2314 21332 2320 21344
rect 2271 21304 2320 21332
rect 2271 21301 2283 21304
rect 2225 21295 2283 21301
rect 2314 21292 2320 21304
rect 2372 21292 2378 21344
rect 3050 21292 3056 21344
rect 3108 21332 3114 21344
rect 4356 21332 4384 21372
rect 6730 21360 6736 21372
rect 6788 21360 6794 21412
rect 8036 21400 8064 21428
rect 9582 21400 9588 21412
rect 8036 21372 9588 21400
rect 9582 21360 9588 21372
rect 9640 21400 9646 21412
rect 10597 21403 10655 21409
rect 10597 21400 10609 21403
rect 9640 21372 10609 21400
rect 9640 21360 9646 21372
rect 10597 21369 10609 21372
rect 10643 21369 10655 21403
rect 10597 21363 10655 21369
rect 10870 21360 10876 21412
rect 10928 21400 10934 21412
rect 12342 21400 12348 21412
rect 10928 21372 12348 21400
rect 10928 21360 10934 21372
rect 12342 21360 12348 21372
rect 12400 21360 12406 21412
rect 12805 21403 12863 21409
rect 12805 21369 12817 21403
rect 12851 21400 12863 21403
rect 14090 21400 14096 21412
rect 12851 21372 14096 21400
rect 12851 21369 12863 21372
rect 12805 21363 12863 21369
rect 14090 21360 14096 21372
rect 14148 21360 14154 21412
rect 14553 21403 14611 21409
rect 14553 21369 14565 21403
rect 14599 21400 14611 21403
rect 15488 21400 15516 21431
rect 15654 21428 15660 21440
rect 15712 21428 15718 21480
rect 14599 21372 15516 21400
rect 14599 21369 14611 21372
rect 14553 21363 14611 21369
rect 4706 21332 4712 21344
rect 3108 21304 4384 21332
rect 4667 21304 4712 21332
rect 3108 21292 3114 21304
rect 4706 21292 4712 21304
rect 4764 21292 4770 21344
rect 4982 21292 4988 21344
rect 5040 21332 5046 21344
rect 5077 21335 5135 21341
rect 5077 21332 5089 21335
rect 5040 21304 5089 21332
rect 5040 21292 5046 21304
rect 5077 21301 5089 21304
rect 5123 21301 5135 21335
rect 6748 21332 6776 21360
rect 11606 21332 11612 21344
rect 6748 21304 11612 21332
rect 5077 21295 5135 21301
rect 11606 21292 11612 21304
rect 11664 21292 11670 21344
rect 12437 21335 12495 21341
rect 12437 21301 12449 21335
rect 12483 21332 12495 21335
rect 12526 21332 12532 21344
rect 12483 21304 12532 21332
rect 12483 21301 12495 21304
rect 12437 21295 12495 21301
rect 12526 21292 12532 21304
rect 12584 21292 12590 21344
rect 12710 21292 12716 21344
rect 12768 21332 12774 21344
rect 13357 21335 13415 21341
rect 13357 21332 13369 21335
rect 12768 21304 13369 21332
rect 12768 21292 12774 21304
rect 13357 21301 13369 21304
rect 13403 21301 13415 21335
rect 14182 21332 14188 21344
rect 14143 21304 14188 21332
rect 13357 21295 13415 21301
rect 14182 21292 14188 21304
rect 14240 21292 14246 21344
rect 15654 21292 15660 21344
rect 15712 21332 15718 21344
rect 15856 21332 15884 21508
rect 18141 21505 18153 21539
rect 18187 21536 18199 21539
rect 18509 21539 18567 21545
rect 18509 21536 18521 21539
rect 18187 21508 18521 21536
rect 18187 21505 18199 21508
rect 18141 21499 18199 21505
rect 18509 21505 18521 21508
rect 18555 21505 18567 21539
rect 18690 21536 18696 21548
rect 18651 21508 18696 21536
rect 18509 21499 18567 21505
rect 18690 21496 18696 21508
rect 18748 21496 18754 21548
rect 18785 21539 18843 21545
rect 18785 21505 18797 21539
rect 18831 21536 18843 21539
rect 18874 21536 18880 21548
rect 18831 21508 18880 21536
rect 18831 21505 18843 21508
rect 18785 21499 18843 21505
rect 18874 21496 18880 21508
rect 18932 21496 18938 21548
rect 19352 21536 19380 21564
rect 19886 21536 19892 21548
rect 19352 21508 19892 21536
rect 19886 21496 19892 21508
rect 19944 21536 19950 21548
rect 21928 21536 21956 21576
rect 23293 21573 23305 21576
rect 23339 21573 23351 21607
rect 24854 21604 24860 21616
rect 23293 21567 23351 21573
rect 23860 21576 24860 21604
rect 19944 21508 21956 21536
rect 22097 21539 22155 21545
rect 19944 21496 19950 21508
rect 22097 21505 22109 21539
rect 22143 21536 22155 21539
rect 22554 21536 22560 21548
rect 22143 21508 22560 21536
rect 22143 21505 22155 21508
rect 22097 21499 22155 21505
rect 22554 21496 22560 21508
rect 22612 21496 22618 21548
rect 22741 21539 22799 21545
rect 22741 21505 22753 21539
rect 22787 21536 22799 21539
rect 23860 21536 23888 21576
rect 24854 21564 24860 21576
rect 24912 21564 24918 21616
rect 26694 21604 26700 21616
rect 24964 21576 26700 21604
rect 24762 21536 24768 21548
rect 22787 21508 23888 21536
rect 24723 21508 24768 21536
rect 22787 21505 22799 21508
rect 22741 21499 22799 21505
rect 24762 21496 24768 21508
rect 24820 21496 24826 21548
rect 24964 21545 24992 21576
rect 24949 21539 25007 21545
rect 24949 21505 24961 21539
rect 24995 21505 25007 21539
rect 26142 21536 26148 21548
rect 26103 21508 26148 21536
rect 24949 21499 25007 21505
rect 26142 21496 26148 21508
rect 26200 21496 26206 21548
rect 26344 21545 26372 21576
rect 26694 21564 26700 21576
rect 26752 21604 26758 21616
rect 27706 21604 27712 21616
rect 26752 21576 27712 21604
rect 26752 21564 26758 21576
rect 27706 21564 27712 21576
rect 27764 21564 27770 21616
rect 26329 21539 26387 21545
rect 26329 21505 26341 21539
rect 26375 21505 26387 21539
rect 27154 21536 27160 21548
rect 27115 21508 27160 21536
rect 26329 21499 26387 21505
rect 27154 21496 27160 21508
rect 27212 21496 27218 21548
rect 27430 21536 27436 21548
rect 27391 21508 27436 21536
rect 27430 21496 27436 21508
rect 27488 21496 27494 21548
rect 27617 21539 27675 21545
rect 27617 21505 27629 21539
rect 27663 21536 27675 21539
rect 27798 21536 27804 21548
rect 27663 21508 27804 21536
rect 27663 21505 27675 21508
rect 27617 21499 27675 21505
rect 27798 21496 27804 21508
rect 27856 21496 27862 21548
rect 28258 21536 28264 21548
rect 28219 21508 28264 21536
rect 28258 21496 28264 21508
rect 28316 21496 28322 21548
rect 16669 21471 16727 21477
rect 16669 21437 16681 21471
rect 16715 21437 16727 21471
rect 19242 21468 19248 21480
rect 16669 21431 16727 21437
rect 17687 21440 19248 21468
rect 15712 21304 15884 21332
rect 15712 21292 15718 21304
rect 16114 21292 16120 21344
rect 16172 21332 16178 21344
rect 16390 21332 16396 21344
rect 16172 21304 16396 21332
rect 16172 21292 16178 21304
rect 16390 21292 16396 21304
rect 16448 21292 16454 21344
rect 16684 21332 16712 21431
rect 17687 21332 17715 21440
rect 19242 21428 19248 21440
rect 19300 21468 19306 21480
rect 19337 21471 19395 21477
rect 19337 21468 19349 21471
rect 19300 21440 19349 21468
rect 19300 21428 19306 21440
rect 19337 21437 19349 21440
rect 19383 21437 19395 21471
rect 19337 21431 19395 21437
rect 22373 21471 22431 21477
rect 22373 21437 22385 21471
rect 22419 21468 22431 21471
rect 23382 21468 23388 21480
rect 22419 21440 23388 21468
rect 22419 21437 22431 21440
rect 22373 21431 22431 21437
rect 23382 21428 23388 21440
rect 23440 21428 23446 21480
rect 25041 21471 25099 21477
rect 25041 21437 25053 21471
rect 25087 21468 25099 21471
rect 25314 21468 25320 21480
rect 25087 21440 25320 21468
rect 25087 21437 25099 21440
rect 25041 21431 25099 21437
rect 25314 21428 25320 21440
rect 25372 21428 25378 21480
rect 25590 21428 25596 21480
rect 25648 21468 25654 21480
rect 26421 21471 26479 21477
rect 26421 21468 26433 21471
rect 25648 21440 26433 21468
rect 25648 21428 25654 21440
rect 26421 21437 26433 21440
rect 26467 21468 26479 21471
rect 27706 21468 27712 21480
rect 26467 21440 27712 21468
rect 26467 21437 26479 21440
rect 26421 21431 26479 21437
rect 27706 21428 27712 21440
rect 27764 21428 27770 21480
rect 28534 21468 28540 21480
rect 28495 21440 28540 21468
rect 28534 21428 28540 21440
rect 28592 21428 28598 21480
rect 28920 21468 28948 21644
rect 29012 21644 31116 21672
rect 29012 21545 29040 21644
rect 31110 21632 31116 21644
rect 31168 21632 31174 21684
rect 29178 21604 29184 21616
rect 29139 21576 29184 21604
rect 29178 21564 29184 21576
rect 29236 21564 29242 21616
rect 29273 21607 29331 21613
rect 29273 21573 29285 21607
rect 29319 21604 29331 21607
rect 29454 21604 29460 21616
rect 29319 21576 29460 21604
rect 29319 21573 29331 21576
rect 29273 21567 29331 21573
rect 29454 21564 29460 21576
rect 29512 21564 29518 21616
rect 28997 21539 29055 21545
rect 28997 21505 29009 21539
rect 29043 21505 29055 21539
rect 28997 21499 29055 21505
rect 29365 21539 29423 21545
rect 29365 21505 29377 21539
rect 29411 21505 29423 21539
rect 29365 21499 29423 21505
rect 29380 21468 29408 21499
rect 30006 21496 30012 21548
rect 30064 21536 30070 21548
rect 30193 21539 30251 21545
rect 30193 21536 30205 21539
rect 30064 21508 30205 21536
rect 30064 21496 30070 21508
rect 30193 21505 30205 21508
rect 30239 21505 30251 21539
rect 30193 21499 30251 21505
rect 30374 21496 30380 21548
rect 30432 21536 30438 21548
rect 30469 21539 30527 21545
rect 30469 21536 30481 21539
rect 30432 21508 30481 21536
rect 30432 21496 30438 21508
rect 30469 21505 30481 21508
rect 30515 21505 30527 21539
rect 30469 21499 30527 21505
rect 30558 21496 30564 21548
rect 30616 21536 30622 21548
rect 30653 21539 30711 21545
rect 30653 21536 30665 21539
rect 30616 21508 30665 21536
rect 30616 21496 30622 21508
rect 30653 21505 30665 21508
rect 30699 21505 30711 21539
rect 30653 21499 30711 21505
rect 30834 21496 30840 21548
rect 30892 21536 30898 21548
rect 31113 21539 31171 21545
rect 31113 21536 31125 21539
rect 30892 21508 31125 21536
rect 30892 21496 30898 21508
rect 31113 21505 31125 21508
rect 31159 21505 31171 21539
rect 31113 21499 31171 21505
rect 30098 21468 30104 21480
rect 28920 21440 30104 21468
rect 30098 21428 30104 21440
rect 30156 21428 30162 21480
rect 17770 21360 17776 21412
rect 17828 21400 17834 21412
rect 18049 21403 18107 21409
rect 18049 21400 18061 21403
rect 17828 21372 18061 21400
rect 17828 21360 17834 21372
rect 18049 21369 18061 21372
rect 18095 21400 18107 21403
rect 18141 21403 18199 21409
rect 18141 21400 18153 21403
rect 18095 21372 18153 21400
rect 18095 21369 18107 21372
rect 18049 21363 18107 21369
rect 18141 21369 18153 21372
rect 18187 21369 18199 21403
rect 18141 21363 18199 21369
rect 20898 21360 20904 21412
rect 20956 21400 20962 21412
rect 24762 21400 24768 21412
rect 20956 21372 24768 21400
rect 20956 21360 20962 21372
rect 24762 21360 24768 21372
rect 24820 21360 24826 21412
rect 27522 21360 27528 21412
rect 27580 21400 27586 21412
rect 28626 21400 28632 21412
rect 27580 21372 28632 21400
rect 27580 21360 27586 21372
rect 28626 21360 28632 21372
rect 28684 21400 28690 21412
rect 31205 21403 31263 21409
rect 31205 21400 31217 21403
rect 28684 21372 31217 21400
rect 28684 21360 28690 21372
rect 31205 21369 31217 21372
rect 31251 21369 31263 21403
rect 31205 21363 31263 21369
rect 16684 21304 17715 21332
rect 18322 21292 18328 21344
rect 18380 21332 18386 21344
rect 18509 21335 18567 21341
rect 18509 21332 18521 21335
rect 18380 21304 18521 21332
rect 18380 21292 18386 21304
rect 18509 21301 18521 21304
rect 18555 21301 18567 21335
rect 18509 21295 18567 21301
rect 18782 21292 18788 21344
rect 18840 21332 18846 21344
rect 22186 21332 22192 21344
rect 18840 21304 22192 21332
rect 18840 21292 18846 21304
rect 22186 21292 22192 21304
rect 22244 21292 22250 21344
rect 22281 21335 22339 21341
rect 22281 21301 22293 21335
rect 22327 21332 22339 21335
rect 22465 21335 22523 21341
rect 22465 21332 22477 21335
rect 22327 21304 22477 21332
rect 22327 21301 22339 21304
rect 22281 21295 22339 21301
rect 22465 21301 22477 21304
rect 22511 21332 22523 21335
rect 22922 21332 22928 21344
rect 22511 21304 22928 21332
rect 22511 21301 22523 21304
rect 22465 21295 22523 21301
rect 22922 21292 22928 21304
rect 22980 21292 22986 21344
rect 24780 21332 24808 21360
rect 25038 21332 25044 21344
rect 24780 21304 25044 21332
rect 25038 21292 25044 21304
rect 25096 21292 25102 21344
rect 26510 21292 26516 21344
rect 26568 21332 26574 21344
rect 26973 21335 27031 21341
rect 26973 21332 26985 21335
rect 26568 21304 26985 21332
rect 26568 21292 26574 21304
rect 26973 21301 26985 21304
rect 27019 21301 27031 21335
rect 26973 21295 27031 21301
rect 27982 21292 27988 21344
rect 28040 21332 28046 21344
rect 28077 21335 28135 21341
rect 28077 21332 28089 21335
rect 28040 21304 28089 21332
rect 28040 21292 28046 21304
rect 28077 21301 28089 21304
rect 28123 21301 28135 21335
rect 28077 21295 28135 21301
rect 28166 21292 28172 21344
rect 28224 21332 28230 21344
rect 28445 21335 28503 21341
rect 28445 21332 28457 21335
rect 28224 21304 28457 21332
rect 28224 21292 28230 21304
rect 28445 21301 28457 21304
rect 28491 21301 28503 21335
rect 28445 21295 28503 21301
rect 28902 21292 28908 21344
rect 28960 21332 28966 21344
rect 29549 21335 29607 21341
rect 29549 21332 29561 21335
rect 28960 21304 29561 21332
rect 28960 21292 28966 21304
rect 29549 21301 29561 21304
rect 29595 21301 29607 21335
rect 29549 21295 29607 21301
rect 30009 21335 30067 21341
rect 30009 21301 30021 21335
rect 30055 21332 30067 21335
rect 30926 21332 30932 21344
rect 30055 21304 30932 21332
rect 30055 21301 30067 21304
rect 30009 21295 30067 21301
rect 30926 21292 30932 21304
rect 30984 21292 30990 21344
rect 1104 21242 32016 21264
rect 1104 21190 2136 21242
rect 2188 21190 12440 21242
rect 12492 21190 22744 21242
rect 22796 21190 32016 21242
rect 1104 21168 32016 21190
rect 2590 21088 2596 21140
rect 2648 21128 2654 21140
rect 2777 21131 2835 21137
rect 2777 21128 2789 21131
rect 2648 21100 2789 21128
rect 2648 21088 2654 21100
rect 2777 21097 2789 21100
rect 2823 21128 2835 21131
rect 2866 21128 2872 21140
rect 2823 21100 2872 21128
rect 2823 21097 2835 21100
rect 2777 21091 2835 21097
rect 2866 21088 2872 21100
rect 2924 21088 2930 21140
rect 3510 21088 3516 21140
rect 3568 21128 3574 21140
rect 6273 21131 6331 21137
rect 3568 21100 6224 21128
rect 3568 21088 3574 21100
rect 768 21032 888 21060
rect 0 20856 800 20870
rect 860 20856 888 21032
rect 5626 21020 5632 21072
rect 5684 21060 5690 21072
rect 5902 21060 5908 21072
rect 5684 21032 5908 21060
rect 5684 21020 5690 21032
rect 5902 21020 5908 21032
rect 5960 21020 5966 21072
rect 6196 21060 6224 21100
rect 6273 21097 6285 21131
rect 6319 21128 6331 21131
rect 8113 21131 8171 21137
rect 6319 21100 8064 21128
rect 6319 21097 6331 21100
rect 6273 21091 6331 21097
rect 7653 21063 7711 21069
rect 7653 21060 7665 21063
rect 6196 21032 7665 21060
rect 7653 21029 7665 21032
rect 7699 21029 7711 21063
rect 8036 21060 8064 21100
rect 8113 21097 8125 21131
rect 8159 21128 8171 21131
rect 8662 21128 8668 21140
rect 8159 21100 8668 21128
rect 8159 21097 8171 21100
rect 8113 21091 8171 21097
rect 8662 21088 8668 21100
rect 8720 21088 8726 21140
rect 9214 21088 9220 21140
rect 9272 21128 9278 21140
rect 10778 21128 10784 21140
rect 9272 21100 10784 21128
rect 9272 21088 9278 21100
rect 10778 21088 10784 21100
rect 10836 21088 10842 21140
rect 11054 21088 11060 21140
rect 11112 21128 11118 21140
rect 11425 21131 11483 21137
rect 11425 21128 11437 21131
rect 11112 21100 11437 21128
rect 11112 21088 11118 21100
rect 11425 21097 11437 21100
rect 11471 21097 11483 21131
rect 17773 21131 17831 21137
rect 11425 21091 11483 21097
rect 12268 21100 16344 21128
rect 9398 21060 9404 21072
rect 8036 21032 9404 21060
rect 7653 21023 7711 21029
rect 9398 21020 9404 21032
rect 9456 21020 9462 21072
rect 9674 21020 9680 21072
rect 9732 21060 9738 21072
rect 10045 21063 10103 21069
rect 10045 21060 10057 21063
rect 9732 21032 10057 21060
rect 9732 21020 9738 21032
rect 10045 21029 10057 21032
rect 10091 21029 10103 21063
rect 12268 21060 12296 21100
rect 10045 21023 10103 21029
rect 10888 21032 12296 21060
rect 7190 20952 7196 21004
rect 7248 20992 7254 21004
rect 10888 20992 10916 21032
rect 12342 21020 12348 21072
rect 12400 21060 12406 21072
rect 12894 21060 12900 21072
rect 12400 21032 12900 21060
rect 12400 21020 12406 21032
rect 12894 21020 12900 21032
rect 12952 21020 12958 21072
rect 12158 20992 12164 21004
rect 7248 20964 10916 20992
rect 11164 20964 12164 20992
rect 7248 20952 7254 20964
rect 1397 20927 1455 20933
rect 1397 20893 1409 20927
rect 1443 20924 1455 20927
rect 2774 20924 2780 20936
rect 1443 20896 2780 20924
rect 1443 20893 1455 20896
rect 1397 20887 1455 20893
rect 2774 20884 2780 20896
rect 2832 20884 2838 20936
rect 4157 20927 4215 20933
rect 4157 20893 4169 20927
rect 4203 20924 4215 20927
rect 5626 20924 5632 20936
rect 4203 20896 5632 20924
rect 4203 20893 4215 20896
rect 4157 20887 4215 20893
rect 5626 20884 5632 20896
rect 5684 20884 5690 20936
rect 6457 20927 6515 20933
rect 6457 20893 6469 20927
rect 6503 20893 6515 20927
rect 6457 20887 6515 20893
rect 6549 20927 6607 20933
rect 6549 20893 6561 20927
rect 6595 20893 6607 20927
rect 6730 20924 6736 20936
rect 6691 20896 6736 20924
rect 6549 20887 6607 20893
rect 0 20828 888 20856
rect 1664 20859 1722 20865
rect 0 20814 800 20828
rect 1664 20825 1676 20859
rect 1710 20856 1722 20859
rect 1854 20856 1860 20868
rect 1710 20828 1860 20856
rect 1710 20825 1722 20828
rect 1664 20819 1722 20825
rect 1854 20816 1860 20828
rect 1912 20816 1918 20868
rect 4424 20859 4482 20865
rect 4424 20825 4436 20859
rect 4470 20856 4482 20859
rect 4706 20856 4712 20868
rect 4470 20828 4712 20856
rect 4470 20825 4482 20828
rect 4424 20819 4482 20825
rect 4706 20816 4712 20828
rect 4764 20816 4770 20868
rect 5074 20816 5080 20868
rect 5132 20856 5138 20868
rect 6472 20856 6500 20887
rect 5132 20828 6500 20856
rect 6564 20856 6592 20887
rect 6730 20884 6736 20896
rect 6788 20884 6794 20936
rect 6822 20884 6828 20936
rect 6880 20924 6886 20936
rect 6880 20896 6925 20924
rect 6880 20884 6886 20896
rect 7466 20884 7472 20936
rect 7524 20924 7530 20936
rect 7745 20927 7803 20933
rect 7745 20924 7757 20927
rect 7524 20896 7757 20924
rect 7524 20884 7530 20896
rect 7745 20893 7757 20896
rect 7791 20893 7803 20927
rect 7745 20887 7803 20893
rect 7834 20884 7840 20936
rect 7892 20924 7898 20936
rect 7929 20927 7987 20933
rect 7929 20924 7941 20927
rect 7892 20896 7941 20924
rect 7892 20884 7898 20896
rect 7929 20893 7941 20896
rect 7975 20893 7987 20927
rect 7929 20887 7987 20893
rect 8570 20884 8576 20936
rect 8628 20924 8634 20936
rect 9214 20924 9220 20936
rect 8628 20896 9220 20924
rect 8628 20884 8634 20896
rect 9214 20884 9220 20896
rect 9272 20924 9278 20936
rect 9309 20927 9367 20933
rect 9309 20924 9321 20927
rect 9272 20896 9321 20924
rect 9272 20884 9278 20896
rect 9309 20893 9321 20896
rect 9355 20893 9367 20927
rect 10686 20924 10692 20936
rect 9683 20914 10272 20924
rect 9309 20887 9367 20893
rect 9646 20896 10272 20914
rect 10647 20896 10692 20924
rect 9646 20886 9711 20896
rect 7006 20856 7012 20868
rect 6564 20828 7012 20856
rect 5132 20816 5138 20828
rect 7006 20816 7012 20828
rect 7064 20816 7070 20868
rect 7558 20816 7564 20868
rect 7616 20816 7622 20868
rect 7653 20859 7711 20865
rect 7653 20825 7665 20859
rect 7699 20856 7711 20859
rect 9646 20856 9674 20886
rect 9766 20856 9772 20868
rect 7699 20828 9674 20856
rect 9727 20828 9772 20856
rect 7699 20825 7711 20828
rect 7653 20819 7711 20825
rect 9766 20816 9772 20828
rect 9824 20816 9830 20868
rect 9950 20816 9956 20868
rect 10008 20856 10014 20868
rect 10244 20856 10272 20896
rect 10686 20884 10692 20896
rect 10744 20884 10750 20936
rect 10873 20927 10931 20933
rect 10873 20893 10885 20927
rect 10919 20924 10931 20927
rect 11164 20924 11192 20964
rect 12158 20952 12164 20964
rect 12216 20992 12222 21004
rect 12529 20995 12587 21001
rect 12529 20992 12541 20995
rect 12216 20964 12541 20992
rect 12216 20952 12222 20964
rect 12529 20961 12541 20964
rect 12575 20961 12587 20995
rect 12529 20955 12587 20961
rect 12802 20952 12808 21004
rect 12860 20992 12866 21004
rect 14737 20995 14795 21001
rect 14737 20992 14749 20995
rect 12860 20964 14749 20992
rect 12860 20952 12866 20964
rect 14737 20961 14749 20964
rect 14783 20961 14795 20995
rect 16316 20992 16344 21100
rect 17773 21097 17785 21131
rect 17819 21128 17831 21131
rect 18414 21128 18420 21140
rect 17819 21100 18420 21128
rect 17819 21097 17831 21100
rect 17773 21091 17831 21097
rect 18414 21088 18420 21100
rect 18472 21088 18478 21140
rect 19245 21131 19303 21137
rect 19245 21097 19257 21131
rect 19291 21128 19303 21131
rect 20622 21128 20628 21140
rect 19291 21100 20628 21128
rect 19291 21097 19303 21100
rect 19245 21091 19303 21097
rect 20622 21088 20628 21100
rect 20680 21088 20686 21140
rect 20714 21088 20720 21140
rect 20772 21128 20778 21140
rect 21266 21128 21272 21140
rect 20772 21100 21272 21128
rect 20772 21088 20778 21100
rect 21266 21088 21272 21100
rect 21324 21128 21330 21140
rect 24026 21128 24032 21140
rect 21324 21100 24032 21128
rect 21324 21088 21330 21100
rect 24026 21088 24032 21100
rect 24084 21128 24090 21140
rect 25777 21131 25835 21137
rect 25777 21128 25789 21131
rect 24084 21100 25789 21128
rect 24084 21088 24090 21100
rect 25777 21097 25789 21100
rect 25823 21097 25835 21131
rect 26694 21128 26700 21140
rect 26655 21100 26700 21128
rect 25777 21091 25835 21097
rect 26694 21088 26700 21100
rect 26752 21088 26758 21140
rect 26804 21100 28033 21128
rect 26804 21060 26832 21100
rect 17236 21032 26832 21060
rect 17236 20992 17264 21032
rect 27338 21020 27344 21072
rect 27396 21060 27402 21072
rect 28005 21060 28033 21100
rect 28534 21088 28540 21140
rect 28592 21128 28598 21140
rect 28997 21131 29055 21137
rect 28997 21128 29009 21131
rect 28592 21100 29009 21128
rect 28592 21088 28598 21100
rect 28997 21097 29009 21100
rect 29043 21097 29055 21131
rect 30742 21128 30748 21140
rect 30703 21100 30748 21128
rect 28997 21091 29055 21097
rect 30742 21088 30748 21100
rect 30800 21088 30806 21140
rect 28074 21060 28080 21072
rect 27396 21032 27933 21060
rect 28005 21032 28080 21060
rect 27396 21020 27402 21032
rect 21910 20992 21916 21004
rect 16316 20964 17264 20992
rect 17328 20964 18276 20992
rect 14737 20955 14795 20961
rect 10919 20896 11192 20924
rect 10919 20893 10931 20896
rect 10873 20887 10931 20893
rect 11238 20884 11244 20936
rect 11296 20924 11302 20936
rect 11333 20927 11391 20933
rect 11333 20924 11345 20927
rect 11296 20896 11345 20924
rect 11296 20884 11302 20896
rect 11333 20893 11345 20896
rect 11379 20893 11391 20927
rect 11333 20887 11391 20893
rect 11790 20884 11796 20936
rect 11848 20924 11854 20936
rect 12066 20924 12072 20936
rect 11848 20896 12072 20924
rect 11848 20884 11854 20896
rect 12066 20884 12072 20896
rect 12124 20884 12130 20936
rect 12250 20924 12256 20936
rect 12211 20896 12256 20924
rect 12250 20884 12256 20896
rect 12308 20884 12314 20936
rect 12342 20884 12348 20936
rect 12400 20924 12406 20936
rect 12710 20924 12716 20936
rect 12400 20896 12716 20924
rect 12400 20884 12406 20896
rect 12710 20884 12716 20896
rect 12768 20884 12774 20936
rect 14090 20924 14096 20936
rect 14051 20896 14096 20924
rect 14090 20884 14096 20896
rect 14148 20884 14154 20936
rect 14277 20927 14335 20933
rect 14277 20893 14289 20927
rect 14323 20924 14335 20927
rect 14366 20924 14372 20936
rect 14323 20896 14372 20924
rect 14323 20893 14335 20896
rect 14277 20887 14335 20893
rect 14366 20884 14372 20896
rect 14424 20884 14430 20936
rect 15010 20933 15016 20936
rect 15004 20924 15016 20933
rect 14971 20896 15016 20924
rect 15004 20887 15016 20896
rect 15010 20884 15016 20887
rect 15068 20884 15074 20936
rect 15930 20924 15936 20936
rect 15120 20896 15936 20924
rect 10781 20859 10839 20865
rect 10008 20828 10180 20856
rect 10244 20828 10732 20856
rect 10008 20816 10014 20828
rect 5537 20791 5595 20797
rect 5537 20757 5549 20791
rect 5583 20788 5595 20791
rect 5718 20788 5724 20800
rect 5583 20760 5724 20788
rect 5583 20757 5595 20760
rect 5537 20751 5595 20757
rect 5718 20748 5724 20760
rect 5776 20748 5782 20800
rect 7576 20788 7604 20816
rect 8570 20788 8576 20800
rect 7576 20760 8576 20788
rect 8570 20748 8576 20760
rect 8628 20748 8634 20800
rect 9125 20791 9183 20797
rect 9125 20757 9137 20791
rect 9171 20788 9183 20791
rect 10042 20788 10048 20800
rect 9171 20760 10048 20788
rect 9171 20757 9183 20760
rect 9125 20751 9183 20757
rect 10042 20748 10048 20760
rect 10100 20748 10106 20800
rect 10152 20788 10180 20828
rect 10229 20791 10287 20797
rect 10229 20788 10241 20791
rect 10152 20760 10241 20788
rect 10229 20757 10241 20760
rect 10275 20757 10287 20791
rect 10704 20788 10732 20828
rect 10781 20825 10793 20859
rect 10827 20856 10839 20859
rect 10827 20828 11376 20856
rect 10827 20825 10839 20828
rect 10781 20819 10839 20825
rect 11054 20788 11060 20800
rect 10704 20760 11060 20788
rect 10229 20751 10287 20757
rect 11054 20748 11060 20760
rect 11112 20748 11118 20800
rect 11348 20788 11376 20828
rect 11974 20816 11980 20868
rect 12032 20856 12038 20868
rect 15120 20856 15148 20896
rect 15930 20884 15936 20896
rect 15988 20884 15994 20936
rect 17126 20924 17132 20936
rect 17087 20896 17132 20924
rect 17126 20884 17132 20896
rect 17184 20918 17190 20936
rect 17328 20924 17356 20964
rect 17297 20918 17356 20924
rect 17184 20896 17356 20918
rect 17398 20927 17456 20933
rect 17184 20890 17325 20896
rect 17398 20893 17410 20927
rect 17444 20924 17456 20927
rect 17589 20927 17647 20933
rect 17444 20896 17540 20924
rect 17444 20893 17456 20896
rect 17184 20884 17190 20890
rect 17398 20887 17456 20893
rect 12032 20828 15148 20856
rect 12032 20816 12038 20828
rect 15378 20816 15384 20868
rect 15436 20856 15442 20868
rect 15746 20856 15752 20868
rect 15436 20828 15752 20856
rect 15436 20816 15442 20828
rect 15746 20816 15752 20828
rect 15804 20856 15810 20868
rect 16298 20856 16304 20868
rect 15804 20828 16304 20856
rect 15804 20816 15810 20828
rect 16298 20816 16304 20828
rect 16356 20816 16362 20868
rect 17512 20856 17540 20896
rect 17589 20893 17601 20927
rect 17635 20924 17647 20927
rect 17678 20924 17684 20936
rect 17635 20896 17684 20924
rect 17635 20893 17647 20896
rect 17589 20887 17647 20893
rect 17678 20884 17684 20896
rect 17736 20924 17742 20936
rect 17770 20924 17776 20936
rect 17736 20896 17776 20924
rect 17736 20884 17742 20896
rect 17770 20884 17776 20896
rect 17828 20884 17834 20936
rect 18046 20924 18052 20936
rect 18007 20896 18052 20924
rect 18046 20884 18052 20896
rect 18104 20884 18110 20936
rect 18248 20933 18276 20964
rect 19720 20964 21916 20992
rect 18233 20927 18291 20933
rect 18233 20893 18245 20927
rect 18279 20924 18291 20927
rect 18414 20924 18420 20936
rect 18279 20896 18420 20924
rect 18279 20893 18291 20896
rect 18233 20887 18291 20893
rect 18414 20884 18420 20896
rect 18472 20884 18478 20936
rect 18509 20927 18567 20933
rect 18509 20893 18521 20927
rect 18555 20893 18567 20927
rect 18690 20924 18696 20936
rect 18651 20896 18696 20924
rect 18509 20887 18567 20893
rect 18138 20856 18144 20868
rect 17512 20828 18144 20856
rect 18138 20816 18144 20828
rect 18196 20856 18202 20868
rect 18524 20856 18552 20887
rect 18690 20884 18696 20896
rect 18748 20884 18754 20936
rect 19426 20924 19432 20936
rect 19387 20896 19432 20924
rect 19426 20884 19432 20896
rect 19484 20884 19490 20936
rect 19720 20933 19748 20964
rect 21910 20952 21916 20964
rect 21968 20952 21974 21004
rect 22370 20952 22376 21004
rect 22428 20992 22434 21004
rect 22557 20995 22615 21001
rect 22557 20992 22569 20995
rect 22428 20964 22569 20992
rect 22428 20952 22434 20964
rect 22557 20961 22569 20964
rect 22603 20961 22615 20995
rect 23106 20992 23112 21004
rect 23067 20964 23112 20992
rect 22557 20955 22615 20961
rect 23106 20952 23112 20964
rect 23164 20952 23170 21004
rect 23201 20995 23259 21001
rect 23201 20961 23213 20995
rect 23247 20961 23259 20995
rect 23201 20955 23259 20961
rect 25041 20995 25099 21001
rect 25041 20961 25053 20995
rect 25087 20992 25099 20995
rect 26418 20992 26424 21004
rect 25087 20964 26424 20992
rect 25087 20961 25099 20964
rect 25041 20955 25099 20961
rect 19705 20927 19763 20933
rect 19705 20893 19717 20927
rect 19751 20893 19763 20927
rect 19705 20887 19763 20893
rect 19889 20927 19947 20933
rect 19889 20893 19901 20927
rect 19935 20924 19947 20927
rect 20990 20924 20996 20936
rect 19935 20896 20996 20924
rect 19935 20893 19947 20896
rect 19889 20887 19947 20893
rect 20990 20884 20996 20896
rect 21048 20884 21054 20936
rect 21542 20884 21548 20936
rect 21600 20924 21606 20936
rect 22462 20924 22468 20936
rect 21600 20896 22468 20924
rect 21600 20884 21606 20896
rect 22462 20884 22468 20896
rect 22520 20924 22526 20936
rect 23216 20924 23244 20955
rect 26418 20952 26424 20964
rect 26476 20952 26482 21004
rect 26789 20995 26847 21001
rect 26789 20961 26801 20995
rect 26835 20992 26847 20995
rect 27246 20992 27252 21004
rect 26835 20964 27252 20992
rect 26835 20961 26847 20964
rect 26789 20955 26847 20961
rect 27246 20952 27252 20964
rect 27304 20992 27310 21004
rect 27905 20992 27933 21032
rect 28074 21020 28080 21032
rect 28132 21020 28138 21072
rect 28166 21020 28172 21072
rect 28224 21060 28230 21072
rect 30285 21063 30343 21069
rect 30285 21060 30297 21063
rect 28224 21032 28269 21060
rect 28644 21032 30297 21060
rect 28224 21020 28230 21032
rect 27304 20964 27660 20992
rect 27905 20964 28033 20992
rect 27304 20952 27310 20964
rect 24762 20924 24768 20936
rect 22520 20896 23244 20924
rect 24723 20896 24768 20924
rect 22520 20884 22526 20896
rect 24762 20884 24768 20896
rect 24820 20884 24826 20936
rect 24946 20924 24952 20936
rect 24907 20896 24952 20924
rect 24946 20884 24952 20896
rect 25004 20884 25010 20936
rect 25593 20927 25651 20933
rect 25593 20924 25605 20927
rect 25148 20896 25605 20924
rect 25148 20868 25176 20896
rect 25593 20893 25605 20896
rect 25639 20893 25651 20927
rect 26510 20924 26516 20936
rect 26471 20896 26516 20924
rect 25593 20887 25651 20893
rect 26510 20884 26516 20896
rect 26568 20884 26574 20936
rect 27522 20924 27528 20936
rect 27483 20896 27528 20924
rect 27522 20884 27528 20896
rect 27580 20884 27586 20936
rect 27632 20933 27660 20964
rect 27618 20927 27676 20933
rect 27618 20893 27630 20927
rect 27664 20893 27676 20927
rect 27618 20887 27676 20893
rect 27706 20884 27712 20936
rect 27764 20924 27770 20936
rect 28005 20933 28033 20964
rect 28534 20952 28540 21004
rect 28592 20992 28598 21004
rect 28644 20992 28672 21032
rect 30285 21029 30297 21032
rect 30331 21029 30343 21063
rect 30285 21023 30343 21029
rect 31205 20995 31263 21001
rect 31205 20992 31217 20995
rect 28592 20964 28672 20992
rect 28736 20964 28994 20992
rect 28592 20952 28598 20964
rect 27990 20927 28048 20933
rect 27764 20896 27927 20924
rect 27764 20884 27770 20896
rect 18966 20856 18972 20868
rect 18196 20828 18972 20856
rect 18196 20816 18202 20828
rect 18966 20816 18972 20828
rect 19024 20816 19030 20868
rect 19150 20816 19156 20868
rect 19208 20856 19214 20868
rect 19610 20856 19616 20868
rect 19208 20828 19616 20856
rect 19208 20816 19214 20828
rect 19610 20816 19616 20828
rect 19668 20816 19674 20868
rect 20438 20856 20444 20868
rect 20399 20828 20444 20856
rect 20438 20816 20444 20828
rect 20496 20816 20502 20868
rect 22370 20856 22376 20868
rect 20548 20828 22376 20856
rect 12526 20788 12532 20800
rect 11348 20760 12532 20788
rect 12526 20748 12532 20760
rect 12584 20748 12590 20800
rect 13722 20748 13728 20800
rect 13780 20788 13786 20800
rect 14185 20791 14243 20797
rect 14185 20788 14197 20791
rect 13780 20760 14197 20788
rect 13780 20748 13786 20760
rect 14185 20757 14197 20760
rect 14231 20757 14243 20791
rect 14185 20751 14243 20757
rect 14918 20748 14924 20800
rect 14976 20788 14982 20800
rect 16117 20791 16175 20797
rect 16117 20788 16129 20791
rect 14976 20760 16129 20788
rect 14976 20748 14982 20760
rect 16117 20757 16129 20760
rect 16163 20757 16175 20791
rect 16942 20788 16948 20800
rect 16903 20760 16948 20788
rect 16117 20751 16175 20757
rect 16942 20748 16948 20760
rect 17000 20748 17006 20800
rect 17034 20748 17040 20800
rect 17092 20788 17098 20800
rect 17218 20788 17224 20800
rect 17092 20760 17224 20788
rect 17092 20748 17098 20760
rect 17218 20748 17224 20760
rect 17276 20748 17282 20800
rect 17770 20788 17776 20800
rect 17731 20760 17776 20788
rect 17770 20748 17776 20760
rect 17828 20748 17834 20800
rect 17862 20748 17868 20800
rect 17920 20788 17926 20800
rect 19334 20788 19340 20800
rect 17920 20760 19340 20788
rect 17920 20748 17926 20760
rect 19334 20748 19340 20760
rect 19392 20748 19398 20800
rect 20254 20748 20260 20800
rect 20312 20788 20318 20800
rect 20548 20788 20576 20828
rect 22370 20816 22376 20828
rect 22428 20816 22434 20868
rect 23017 20859 23075 20865
rect 23017 20856 23029 20859
rect 22480 20828 23029 20856
rect 20312 20760 20576 20788
rect 20312 20748 20318 20760
rect 20806 20748 20812 20800
rect 20864 20788 20870 20800
rect 21729 20791 21787 20797
rect 21729 20788 21741 20791
rect 20864 20760 21741 20788
rect 20864 20748 20870 20760
rect 21729 20757 21741 20760
rect 21775 20757 21787 20791
rect 21729 20751 21787 20757
rect 21818 20748 21824 20800
rect 21876 20788 21882 20800
rect 22480 20788 22508 20828
rect 23017 20825 23029 20828
rect 23063 20825 23075 20859
rect 23017 20819 23075 20825
rect 25130 20816 25136 20868
rect 25188 20856 25194 20868
rect 25188 20828 25233 20856
rect 25188 20816 25194 20828
rect 27430 20816 27436 20868
rect 27488 20856 27494 20868
rect 27899 20865 27927 20896
rect 27990 20893 28002 20927
rect 28036 20893 28048 20927
rect 27990 20887 28048 20893
rect 28442 20884 28448 20936
rect 28500 20924 28506 20936
rect 28629 20927 28687 20933
rect 28629 20924 28641 20927
rect 28500 20896 28641 20924
rect 28500 20884 28506 20896
rect 28629 20893 28641 20896
rect 28675 20893 28687 20927
rect 28629 20887 28687 20893
rect 27801 20859 27859 20865
rect 27801 20856 27813 20859
rect 27488 20828 27813 20856
rect 27488 20816 27494 20828
rect 27801 20825 27813 20828
rect 27847 20825 27859 20859
rect 27801 20819 27859 20825
rect 27893 20859 27951 20865
rect 27893 20825 27905 20859
rect 27939 20825 27951 20859
rect 27893 20819 27951 20825
rect 28166 20816 28172 20868
rect 28224 20856 28230 20868
rect 28736 20856 28764 20964
rect 28813 20927 28871 20933
rect 28813 20893 28825 20927
rect 28859 20893 28871 20927
rect 28813 20887 28871 20893
rect 28224 20828 28764 20856
rect 28224 20816 28230 20828
rect 21876 20760 22508 20788
rect 22557 20791 22615 20797
rect 21876 20748 21882 20760
rect 22557 20757 22569 20791
rect 22603 20788 22615 20791
rect 22649 20791 22707 20797
rect 22649 20788 22661 20791
rect 22603 20760 22661 20788
rect 22603 20757 22615 20760
rect 22557 20751 22615 20757
rect 22649 20757 22661 20760
rect 22695 20757 22707 20791
rect 22649 20751 22707 20757
rect 26142 20748 26148 20800
rect 26200 20788 26206 20800
rect 26329 20791 26387 20797
rect 26329 20788 26341 20791
rect 26200 20760 26341 20788
rect 26200 20748 26206 20760
rect 26329 20757 26341 20760
rect 26375 20757 26387 20791
rect 26329 20751 26387 20757
rect 27246 20748 27252 20800
rect 27304 20788 27310 20800
rect 28828 20788 28856 20887
rect 27304 20760 28856 20788
rect 28966 20788 28994 20964
rect 30024 20964 31217 20992
rect 29638 20924 29644 20936
rect 29599 20896 29644 20924
rect 29638 20884 29644 20896
rect 29696 20884 29702 20936
rect 29789 20927 29847 20933
rect 29789 20893 29801 20927
rect 29835 20924 29847 20927
rect 30024 20924 30052 20964
rect 31205 20961 31217 20964
rect 31251 20992 31263 20995
rect 31294 20992 31300 21004
rect 31251 20964 31300 20992
rect 31251 20961 31263 20964
rect 31205 20955 31263 20961
rect 31294 20952 31300 20964
rect 31352 20952 31358 21004
rect 29835 20896 30052 20924
rect 29835 20893 29847 20896
rect 29789 20887 29847 20893
rect 30098 20884 30104 20936
rect 30156 20933 30162 20936
rect 30156 20924 30164 20933
rect 30926 20924 30932 20936
rect 30156 20896 30201 20924
rect 30887 20896 30932 20924
rect 30156 20887 30164 20896
rect 30156 20884 30162 20887
rect 30926 20884 30932 20896
rect 30984 20884 30990 20936
rect 31113 20927 31171 20933
rect 31113 20893 31125 20927
rect 31159 20893 31171 20927
rect 31113 20887 31171 20893
rect 29454 20816 29460 20868
rect 29512 20856 29518 20868
rect 29917 20859 29975 20865
rect 29917 20856 29929 20859
rect 29512 20828 29929 20856
rect 29512 20816 29518 20828
rect 29917 20825 29929 20828
rect 29963 20825 29975 20859
rect 29917 20819 29975 20825
rect 30009 20859 30067 20865
rect 30009 20825 30021 20859
rect 30055 20856 30067 20859
rect 30466 20856 30472 20868
rect 30055 20828 30472 20856
rect 30055 20825 30067 20828
rect 30009 20819 30067 20825
rect 30466 20816 30472 20828
rect 30524 20816 30530 20868
rect 31128 20856 31156 20887
rect 31202 20856 31208 20868
rect 31128 20828 31208 20856
rect 31202 20816 31208 20828
rect 31260 20816 31266 20868
rect 32320 20856 33120 20870
rect 31726 20828 33120 20856
rect 31726 20788 31754 20828
rect 32320 20814 33120 20828
rect 28966 20760 31754 20788
rect 27304 20748 27310 20760
rect 1104 20698 32016 20720
rect 1104 20646 7288 20698
rect 7340 20646 17592 20698
rect 17644 20646 27896 20698
rect 27948 20646 32016 20698
rect 1104 20624 32016 20646
rect 1854 20584 1860 20596
rect 1815 20556 1860 20584
rect 1854 20544 1860 20556
rect 1912 20544 1918 20596
rect 2038 20544 2044 20596
rect 2096 20584 2102 20596
rect 5074 20584 5080 20596
rect 2096 20556 3924 20584
rect 5035 20556 5080 20584
rect 2096 20544 2102 20556
rect 1670 20476 1676 20528
rect 1728 20516 1734 20528
rect 1728 20488 3832 20516
rect 1728 20476 1734 20488
rect 2038 20448 2044 20460
rect 1999 20420 2044 20448
rect 2038 20408 2044 20420
rect 2096 20408 2102 20460
rect 2222 20408 2228 20460
rect 2280 20448 2286 20460
rect 2682 20448 2688 20460
rect 2280 20420 2688 20448
rect 2280 20408 2286 20420
rect 2682 20408 2688 20420
rect 2740 20448 2746 20460
rect 3329 20451 3387 20457
rect 3329 20448 3341 20451
rect 2740 20420 3341 20448
rect 2740 20408 2746 20420
rect 3329 20417 3341 20420
rect 3375 20417 3387 20451
rect 3329 20411 3387 20417
rect 2317 20383 2375 20389
rect 2317 20349 2329 20383
rect 2363 20380 2375 20383
rect 2590 20380 2596 20392
rect 2363 20352 2596 20380
rect 2363 20349 2375 20352
rect 2317 20343 2375 20349
rect 2590 20340 2596 20352
rect 2648 20340 2654 20392
rect 3050 20380 3056 20392
rect 3011 20352 3056 20380
rect 3050 20340 3056 20352
rect 3108 20340 3114 20392
rect 2222 20244 2228 20256
rect 2183 20216 2228 20244
rect 2222 20204 2228 20216
rect 2280 20204 2286 20256
rect 3804 20244 3832 20488
rect 3896 20380 3924 20556
rect 5074 20544 5080 20556
rect 5132 20544 5138 20596
rect 5537 20587 5595 20593
rect 5537 20553 5549 20587
rect 5583 20584 5595 20587
rect 6178 20584 6184 20596
rect 5583 20556 6184 20584
rect 5583 20553 5595 20556
rect 5537 20547 5595 20553
rect 6178 20544 6184 20556
rect 6236 20544 6242 20596
rect 6822 20544 6828 20596
rect 6880 20584 6886 20596
rect 6880 20556 8294 20584
rect 6880 20544 6886 20556
rect 4617 20519 4675 20525
rect 4617 20485 4629 20519
rect 4663 20516 4675 20519
rect 4982 20516 4988 20528
rect 4663 20488 4988 20516
rect 4663 20485 4675 20488
rect 4617 20479 4675 20485
rect 4982 20476 4988 20488
rect 5040 20476 5046 20528
rect 6638 20476 6644 20528
rect 6696 20516 6702 20528
rect 6696 20488 7052 20516
rect 6696 20476 6702 20488
rect 4433 20451 4491 20457
rect 4433 20417 4445 20451
rect 4479 20448 4491 20451
rect 4706 20448 4712 20460
rect 4479 20420 4712 20448
rect 4479 20417 4491 20420
rect 4433 20411 4491 20417
rect 4706 20408 4712 20420
rect 4764 20408 4770 20460
rect 5350 20408 5356 20460
rect 5408 20448 5414 20460
rect 5445 20451 5503 20457
rect 5445 20448 5457 20451
rect 5408 20420 5457 20448
rect 5408 20408 5414 20420
rect 5445 20417 5457 20420
rect 5491 20417 5503 20451
rect 6914 20448 6920 20460
rect 5445 20411 5503 20417
rect 5552 20420 5764 20448
rect 6875 20420 6920 20448
rect 4246 20380 4252 20392
rect 3896 20352 4252 20380
rect 4246 20340 4252 20352
rect 4304 20380 4310 20392
rect 5552 20380 5580 20420
rect 4304 20352 5580 20380
rect 5629 20383 5687 20389
rect 4304 20340 4310 20352
rect 5629 20349 5641 20383
rect 5675 20349 5687 20383
rect 5736 20380 5764 20420
rect 6914 20408 6920 20420
rect 6972 20408 6978 20460
rect 7024 20448 7052 20488
rect 7374 20476 7380 20528
rect 7432 20516 7438 20528
rect 8110 20516 8116 20528
rect 7432 20488 8116 20516
rect 7432 20476 7438 20488
rect 8110 20476 8116 20488
rect 8168 20476 8174 20528
rect 8266 20516 8294 20556
rect 8478 20544 8484 20596
rect 8536 20584 8542 20596
rect 8536 20556 9444 20584
rect 8536 20544 8542 20556
rect 9416 20525 9444 20556
rect 9766 20544 9772 20596
rect 9824 20584 9830 20596
rect 9929 20587 9987 20593
rect 9929 20584 9941 20587
rect 9824 20556 9941 20584
rect 9824 20544 9830 20556
rect 9929 20553 9941 20556
rect 9975 20553 9987 20587
rect 9929 20547 9987 20553
rect 10045 20587 10103 20593
rect 10045 20553 10057 20587
rect 10091 20584 10103 20587
rect 10502 20584 10508 20596
rect 10091 20556 10508 20584
rect 10091 20553 10103 20556
rect 10045 20547 10103 20553
rect 10502 20544 10508 20556
rect 10560 20544 10566 20596
rect 10686 20544 10692 20596
rect 10744 20584 10750 20596
rect 10873 20587 10931 20593
rect 10873 20584 10885 20587
rect 10744 20556 10885 20584
rect 10744 20544 10750 20556
rect 10873 20553 10885 20556
rect 10919 20553 10931 20587
rect 11238 20584 11244 20596
rect 10873 20547 10931 20553
rect 10980 20556 11244 20584
rect 9401 20519 9459 20525
rect 8266 20488 8800 20516
rect 7929 20451 7987 20457
rect 7929 20448 7941 20451
rect 7024 20420 7144 20448
rect 7116 20389 7144 20420
rect 7300 20420 7941 20448
rect 7009 20383 7067 20389
rect 7009 20380 7021 20383
rect 5736 20352 7021 20380
rect 5629 20343 5687 20349
rect 7009 20349 7021 20352
rect 7055 20349 7067 20383
rect 7009 20343 7067 20349
rect 7101 20383 7159 20389
rect 7101 20349 7113 20383
rect 7147 20349 7159 20383
rect 7101 20343 7159 20349
rect 5166 20272 5172 20324
rect 5224 20312 5230 20324
rect 5644 20312 5672 20343
rect 5224 20284 5672 20312
rect 6549 20315 6607 20321
rect 5224 20272 5230 20284
rect 6549 20281 6561 20315
rect 6595 20312 6607 20315
rect 7300 20312 7328 20420
rect 7929 20417 7941 20420
rect 7975 20417 7987 20451
rect 7929 20411 7987 20417
rect 8018 20408 8024 20460
rect 8076 20448 8082 20460
rect 8202 20448 8208 20460
rect 8076 20420 8121 20448
rect 8163 20420 8208 20448
rect 8076 20408 8082 20420
rect 8202 20408 8208 20420
rect 8260 20408 8266 20460
rect 8772 20457 8800 20488
rect 9401 20485 9413 20519
rect 9447 20485 9459 20519
rect 9585 20519 9643 20525
rect 9585 20516 9597 20519
rect 9401 20479 9459 20485
rect 9508 20488 9597 20516
rect 8297 20451 8355 20457
rect 8297 20417 8309 20451
rect 8343 20417 8355 20451
rect 8297 20411 8355 20417
rect 8757 20451 8815 20457
rect 8757 20417 8769 20451
rect 8803 20448 8815 20451
rect 9030 20448 9036 20460
rect 8803 20420 9036 20448
rect 8803 20417 8815 20420
rect 8757 20411 8815 20417
rect 8312 20380 8340 20411
rect 9030 20408 9036 20420
rect 9088 20408 9094 20460
rect 9122 20408 9128 20460
rect 9180 20448 9186 20460
rect 9508 20448 9536 20488
rect 9585 20485 9597 20488
rect 9631 20516 9643 20519
rect 10980 20516 11008 20556
rect 11238 20544 11244 20556
rect 11296 20544 11302 20596
rect 11330 20544 11336 20596
rect 11388 20584 11394 20596
rect 12989 20587 13047 20593
rect 11388 20556 11928 20584
rect 11388 20544 11394 20556
rect 11900 20528 11928 20556
rect 12989 20553 13001 20587
rect 13035 20584 13047 20587
rect 17218 20584 17224 20596
rect 13035 20556 17224 20584
rect 13035 20553 13047 20556
rect 12989 20547 13047 20553
rect 17218 20544 17224 20556
rect 17276 20544 17282 20596
rect 18598 20584 18604 20596
rect 17972 20556 18604 20584
rect 9631 20488 11008 20516
rect 9631 20485 9643 20488
rect 9585 20479 9643 20485
rect 11054 20476 11060 20528
rect 11112 20516 11118 20528
rect 11112 20488 11468 20516
rect 11112 20476 11118 20488
rect 9180 20420 9536 20448
rect 9841 20451 9899 20457
rect 9180 20408 9186 20420
rect 9841 20417 9853 20451
rect 9887 20448 9899 20451
rect 9950 20448 9956 20460
rect 9887 20420 9956 20448
rect 9887 20417 9899 20420
rect 9841 20411 9899 20417
rect 9950 20408 9956 20420
rect 10008 20408 10014 20460
rect 10137 20451 10195 20457
rect 10137 20417 10149 20451
rect 10183 20417 10195 20451
rect 10137 20411 10195 20417
rect 8849 20383 8907 20389
rect 8849 20380 8861 20383
rect 8036 20352 8861 20380
rect 6595 20284 7328 20312
rect 6595 20281 6607 20284
rect 6549 20275 6607 20281
rect 7650 20272 7656 20324
rect 7708 20312 7714 20324
rect 8036 20312 8064 20352
rect 8849 20349 8861 20352
rect 8895 20349 8907 20383
rect 10152 20380 10180 20411
rect 10778 20408 10784 20460
rect 10836 20448 10842 20460
rect 11333 20451 11391 20457
rect 11333 20448 11345 20451
rect 10836 20420 11345 20448
rect 10836 20408 10842 20420
rect 11333 20417 11345 20420
rect 11379 20417 11391 20451
rect 11333 20411 11391 20417
rect 11238 20380 11244 20392
rect 10152 20352 11244 20380
rect 8849 20343 8907 20349
rect 11238 20340 11244 20352
rect 11296 20340 11302 20392
rect 11440 20380 11468 20488
rect 11882 20476 11888 20528
rect 11940 20516 11946 20528
rect 12897 20519 12955 20525
rect 12897 20516 12909 20519
rect 11940 20488 12909 20516
rect 11940 20476 11946 20488
rect 12897 20485 12909 20488
rect 12943 20485 12955 20519
rect 12897 20479 12955 20485
rect 13808 20519 13866 20525
rect 13808 20485 13820 20519
rect 13854 20516 13866 20519
rect 14182 20516 14188 20528
rect 13854 20488 14188 20516
rect 13854 20485 13866 20488
rect 13808 20479 13866 20485
rect 14182 20476 14188 20488
rect 14240 20476 14246 20528
rect 14550 20476 14556 20528
rect 14608 20516 14614 20528
rect 15102 20516 15108 20528
rect 14608 20488 15108 20516
rect 14608 20476 14614 20488
rect 15102 20476 15108 20488
rect 15160 20476 15166 20528
rect 15470 20476 15476 20528
rect 15528 20516 15534 20528
rect 16114 20516 16120 20528
rect 15528 20488 16120 20516
rect 15528 20476 15534 20488
rect 16114 20476 16120 20488
rect 16172 20476 16178 20528
rect 16485 20519 16543 20525
rect 16485 20485 16497 20519
rect 16531 20516 16543 20519
rect 16666 20516 16672 20528
rect 16531 20488 16672 20516
rect 16531 20485 16543 20488
rect 16485 20479 16543 20485
rect 16666 20476 16672 20488
rect 16724 20476 16730 20528
rect 16758 20476 16764 20528
rect 16816 20516 16822 20528
rect 17865 20519 17923 20525
rect 17865 20516 17877 20519
rect 16816 20488 17877 20516
rect 16816 20476 16822 20488
rect 17865 20485 17877 20488
rect 17911 20485 17923 20519
rect 17865 20479 17923 20485
rect 11606 20448 11612 20460
rect 11567 20420 11612 20448
rect 11606 20408 11612 20420
rect 11664 20408 11670 20460
rect 11790 20448 11796 20460
rect 11716 20420 11796 20448
rect 11716 20380 11744 20420
rect 11790 20408 11796 20420
rect 11848 20408 11854 20460
rect 12158 20448 12164 20460
rect 12119 20420 12164 20448
rect 12158 20408 12164 20420
rect 12216 20448 12222 20460
rect 12526 20448 12532 20460
rect 12216 20420 12532 20448
rect 12216 20408 12222 20420
rect 12526 20408 12532 20420
rect 12584 20408 12590 20460
rect 14918 20408 14924 20460
rect 14976 20448 14982 20460
rect 15378 20448 15384 20460
rect 14976 20420 15384 20448
rect 14976 20408 14982 20420
rect 15378 20408 15384 20420
rect 15436 20408 15442 20460
rect 15565 20451 15623 20457
rect 15565 20417 15577 20451
rect 15611 20448 15623 20451
rect 15654 20448 15660 20460
rect 15611 20420 15660 20448
rect 15611 20417 15623 20420
rect 15565 20411 15623 20417
rect 15654 20408 15660 20420
rect 15712 20408 15718 20460
rect 16022 20408 16028 20460
rect 16080 20408 16086 20460
rect 16853 20451 16911 20457
rect 16853 20448 16865 20451
rect 16592 20420 16865 20448
rect 11440 20352 11744 20380
rect 11885 20383 11943 20389
rect 11885 20349 11897 20383
rect 11931 20349 11943 20383
rect 11885 20343 11943 20349
rect 11977 20383 12035 20389
rect 11977 20349 11989 20383
rect 12023 20380 12035 20383
rect 12342 20380 12348 20392
rect 12023 20352 12348 20380
rect 12023 20349 12035 20352
rect 11977 20343 12035 20349
rect 7708 20284 8064 20312
rect 7708 20272 7714 20284
rect 8110 20272 8116 20324
rect 8168 20312 8174 20324
rect 11517 20315 11575 20321
rect 8168 20284 11192 20312
rect 8168 20272 8174 20284
rect 5350 20244 5356 20256
rect 3804 20216 5356 20244
rect 5350 20204 5356 20216
rect 5408 20204 5414 20256
rect 6914 20204 6920 20256
rect 6972 20244 6978 20256
rect 7374 20244 7380 20256
rect 6972 20216 7380 20244
rect 6972 20204 6978 20216
rect 7374 20204 7380 20216
rect 7432 20204 7438 20256
rect 7745 20247 7803 20253
rect 7745 20213 7757 20247
rect 7791 20244 7803 20247
rect 8478 20244 8484 20256
rect 7791 20216 8484 20244
rect 7791 20213 7803 20216
rect 7745 20207 7803 20213
rect 8478 20204 8484 20216
rect 8536 20204 8542 20256
rect 9398 20204 9404 20256
rect 9456 20244 9462 20256
rect 11054 20244 11060 20256
rect 9456 20216 11060 20244
rect 9456 20204 9462 20216
rect 11054 20204 11060 20216
rect 11112 20204 11118 20256
rect 11164 20244 11192 20284
rect 11517 20281 11529 20315
rect 11563 20312 11575 20315
rect 11698 20312 11704 20324
rect 11563 20284 11704 20312
rect 11563 20281 11575 20284
rect 11517 20275 11575 20281
rect 11698 20272 11704 20284
rect 11756 20272 11762 20324
rect 11900 20312 11928 20343
rect 12342 20340 12348 20352
rect 12400 20340 12406 20392
rect 12802 20340 12808 20392
rect 12860 20380 12866 20392
rect 13541 20383 13599 20389
rect 13541 20380 13553 20383
rect 12860 20352 13553 20380
rect 12860 20340 12866 20352
rect 13541 20349 13553 20352
rect 13587 20349 13599 20383
rect 13541 20343 13599 20349
rect 14642 20340 14648 20392
rect 14700 20380 14706 20392
rect 16040 20380 16068 20408
rect 16592 20380 16620 20420
rect 16853 20417 16865 20420
rect 16899 20417 16911 20451
rect 16853 20411 16911 20417
rect 16942 20408 16948 20460
rect 17000 20448 17006 20460
rect 17972 20457 18000 20556
rect 18598 20544 18604 20556
rect 18656 20544 18662 20596
rect 18874 20544 18880 20596
rect 18932 20584 18938 20596
rect 23474 20584 23480 20596
rect 18932 20556 23143 20584
rect 23435 20556 23480 20584
rect 18932 20544 18938 20556
rect 18230 20525 18236 20528
rect 18213 20519 18236 20525
rect 18213 20485 18225 20519
rect 18213 20479 18236 20485
rect 18230 20476 18236 20479
rect 18288 20476 18294 20528
rect 19429 20519 19487 20525
rect 19429 20516 19441 20519
rect 18708 20488 19441 20516
rect 18708 20460 18736 20488
rect 19429 20485 19441 20488
rect 19475 20485 19487 20519
rect 19429 20479 19487 20485
rect 19610 20476 19616 20528
rect 19668 20516 19674 20528
rect 20070 20516 20076 20528
rect 19668 20488 20076 20516
rect 19668 20476 19674 20488
rect 20070 20476 20076 20488
rect 20128 20516 20134 20528
rect 20128 20488 21312 20516
rect 20128 20476 20134 20488
rect 17221 20451 17279 20457
rect 17000 20420 17045 20448
rect 17000 20408 17006 20420
rect 17221 20417 17233 20451
rect 17267 20417 17279 20451
rect 17221 20411 17279 20417
rect 17957 20451 18015 20457
rect 17957 20417 17969 20451
rect 18003 20417 18015 20451
rect 18690 20448 18696 20460
rect 17957 20411 18015 20417
rect 18064 20420 18696 20448
rect 14700 20352 16620 20380
rect 14700 20340 14706 20352
rect 16666 20340 16672 20392
rect 16724 20380 16730 20392
rect 17236 20380 17264 20411
rect 18064 20380 18092 20420
rect 18690 20408 18696 20420
rect 18748 20408 18754 20460
rect 18966 20408 18972 20460
rect 19024 20448 19030 20460
rect 19024 20420 20116 20448
rect 19024 20408 19030 20420
rect 16724 20352 18092 20380
rect 19797 20383 19855 20389
rect 16724 20340 16730 20352
rect 19797 20349 19809 20383
rect 19843 20380 19855 20383
rect 19978 20380 19984 20392
rect 19843 20352 19984 20380
rect 19843 20349 19855 20352
rect 19797 20343 19855 20349
rect 19978 20340 19984 20352
rect 20036 20340 20042 20392
rect 20088 20389 20116 20420
rect 20714 20408 20720 20460
rect 20772 20448 20778 20460
rect 21284 20457 21312 20488
rect 21450 20476 21456 20528
rect 21508 20516 21514 20528
rect 23115 20516 23143 20556
rect 23474 20544 23480 20556
rect 23532 20544 23538 20596
rect 23661 20587 23719 20593
rect 23661 20553 23673 20587
rect 23707 20584 23719 20587
rect 24578 20584 24584 20596
rect 23707 20556 24584 20584
rect 23707 20553 23719 20556
rect 23661 20547 23719 20553
rect 24578 20544 24584 20556
rect 24636 20544 24642 20596
rect 27246 20584 27252 20596
rect 27207 20556 27252 20584
rect 27246 20544 27252 20556
rect 27304 20544 27310 20596
rect 27614 20584 27620 20596
rect 27575 20556 27620 20584
rect 27614 20544 27620 20556
rect 27672 20544 27678 20596
rect 27709 20587 27767 20593
rect 27709 20553 27721 20587
rect 27755 20584 27767 20587
rect 27798 20584 27804 20596
rect 27755 20556 27804 20584
rect 27755 20553 27767 20556
rect 27709 20547 27767 20553
rect 27798 20544 27804 20556
rect 27856 20544 27862 20596
rect 29086 20584 29092 20596
rect 28966 20556 29092 20584
rect 28966 20516 28994 20556
rect 29086 20544 29092 20556
rect 29144 20544 29150 20596
rect 29178 20544 29184 20596
rect 29236 20544 29242 20596
rect 29638 20544 29644 20596
rect 29696 20584 29702 20596
rect 29825 20587 29883 20593
rect 29825 20584 29837 20587
rect 29696 20556 29837 20584
rect 29696 20544 29702 20556
rect 29825 20553 29837 20556
rect 29871 20553 29883 20587
rect 29825 20547 29883 20553
rect 30193 20587 30251 20593
rect 30193 20553 30205 20587
rect 30239 20584 30251 20587
rect 31110 20584 31116 20596
rect 30239 20556 31116 20584
rect 30239 20553 30251 20556
rect 30193 20547 30251 20553
rect 31110 20544 31116 20556
rect 31168 20544 31174 20596
rect 21508 20488 23060 20516
rect 23115 20488 28994 20516
rect 29196 20516 29224 20544
rect 29196 20488 30328 20516
rect 21508 20476 21514 20488
rect 21085 20451 21143 20457
rect 21085 20448 21097 20451
rect 20772 20420 21097 20448
rect 20772 20408 20778 20420
rect 21085 20417 21097 20420
rect 21131 20417 21143 20451
rect 21085 20411 21143 20417
rect 21269 20451 21327 20457
rect 21269 20417 21281 20451
rect 21315 20417 21327 20451
rect 21269 20411 21327 20417
rect 21818 20408 21824 20460
rect 21876 20448 21882 20460
rect 22005 20451 22063 20457
rect 22005 20448 22017 20451
rect 21876 20420 22017 20448
rect 21876 20408 21882 20420
rect 22005 20417 22017 20420
rect 22051 20417 22063 20451
rect 22005 20411 22063 20417
rect 22189 20451 22247 20457
rect 22189 20417 22201 20451
rect 22235 20448 22247 20451
rect 22922 20448 22928 20460
rect 22235 20420 22928 20448
rect 22235 20417 22247 20420
rect 22189 20411 22247 20417
rect 22922 20408 22928 20420
rect 22980 20408 22986 20460
rect 20073 20383 20131 20389
rect 20073 20349 20085 20383
rect 20119 20349 20131 20383
rect 20990 20380 20996 20392
rect 20073 20343 20131 20349
rect 20180 20352 20996 20380
rect 12158 20312 12164 20324
rect 11900 20284 12164 20312
rect 12158 20272 12164 20284
rect 12216 20272 12222 20324
rect 14921 20315 14979 20321
rect 14921 20281 14933 20315
rect 14967 20312 14979 20315
rect 15562 20312 15568 20324
rect 14967 20284 15568 20312
rect 14967 20281 14979 20284
rect 14921 20275 14979 20281
rect 15562 20272 15568 20284
rect 15620 20312 15626 20324
rect 16022 20312 16028 20324
rect 15620 20284 16028 20312
rect 15620 20272 15626 20284
rect 16022 20272 16028 20284
rect 16080 20272 16086 20324
rect 16298 20272 16304 20324
rect 16356 20312 16362 20324
rect 16485 20315 16543 20321
rect 16485 20312 16497 20315
rect 16356 20284 16497 20312
rect 16356 20272 16362 20284
rect 16485 20281 16497 20284
rect 16531 20312 16543 20315
rect 17129 20315 17187 20321
rect 17129 20312 17141 20315
rect 16531 20284 17141 20312
rect 16531 20281 16543 20284
rect 16485 20275 16543 20281
rect 17129 20281 17141 20284
rect 17175 20281 17187 20315
rect 20180 20312 20208 20352
rect 20990 20340 20996 20352
rect 21048 20340 21054 20392
rect 21726 20340 21732 20392
rect 21784 20380 21790 20392
rect 22281 20383 22339 20389
rect 22281 20380 22293 20383
rect 21784 20352 22293 20380
rect 21784 20340 21790 20352
rect 22281 20349 22293 20352
rect 22327 20349 22339 20383
rect 23032 20380 23060 20488
rect 23109 20451 23167 20457
rect 23109 20417 23121 20451
rect 23155 20448 23167 20451
rect 23750 20448 23756 20460
rect 23155 20420 23756 20448
rect 23155 20417 23167 20420
rect 23109 20411 23167 20417
rect 23750 20408 23756 20420
rect 23808 20408 23814 20460
rect 24121 20451 24179 20457
rect 24121 20417 24133 20451
rect 24167 20448 24179 20451
rect 24762 20448 24768 20460
rect 24167 20420 24768 20448
rect 24167 20417 24179 20420
rect 24121 20411 24179 20417
rect 24762 20408 24768 20420
rect 24820 20408 24826 20460
rect 24854 20408 24860 20460
rect 24912 20448 24918 20460
rect 25317 20451 25375 20457
rect 25317 20448 25329 20451
rect 24912 20420 25329 20448
rect 24912 20408 24918 20420
rect 25317 20417 25329 20420
rect 25363 20417 25375 20451
rect 25317 20411 25375 20417
rect 26145 20451 26203 20457
rect 26145 20417 26157 20451
rect 26191 20448 26203 20451
rect 26970 20448 26976 20460
rect 26191 20420 26976 20448
rect 26191 20417 26203 20420
rect 26145 20411 26203 20417
rect 26970 20408 26976 20420
rect 27028 20408 27034 20460
rect 29089 20451 29147 20457
rect 29089 20448 29101 20451
rect 27816 20420 29101 20448
rect 24210 20380 24216 20392
rect 23032 20352 24216 20380
rect 22281 20343 22339 20349
rect 24210 20340 24216 20352
rect 24268 20380 24274 20392
rect 24305 20383 24363 20389
rect 24305 20380 24317 20383
rect 24268 20352 24317 20380
rect 24268 20340 24274 20352
rect 24305 20349 24317 20352
rect 24351 20349 24363 20383
rect 24305 20343 24363 20349
rect 25133 20383 25191 20389
rect 25133 20349 25145 20383
rect 25179 20380 25191 20383
rect 25406 20380 25412 20392
rect 25179 20352 25412 20380
rect 25179 20349 25191 20352
rect 25133 20343 25191 20349
rect 25406 20340 25412 20352
rect 25464 20340 25470 20392
rect 25590 20340 25596 20392
rect 25648 20380 25654 20392
rect 26421 20383 26479 20389
rect 26421 20380 26433 20383
rect 25648 20352 26433 20380
rect 25648 20340 25654 20352
rect 26421 20349 26433 20352
rect 26467 20349 26479 20383
rect 26421 20343 26479 20349
rect 27706 20340 27712 20392
rect 27764 20380 27770 20392
rect 27816 20389 27844 20420
rect 29089 20417 29101 20420
rect 29135 20417 29147 20451
rect 29089 20411 29147 20417
rect 29181 20454 29239 20457
rect 29181 20451 29316 20454
rect 29181 20417 29193 20451
rect 29227 20448 29316 20451
rect 29730 20448 29736 20460
rect 29227 20426 29736 20448
rect 29227 20417 29239 20426
rect 29288 20420 29736 20426
rect 29181 20411 29239 20417
rect 29730 20408 29736 20420
rect 29788 20408 29794 20460
rect 30300 20457 30328 20488
rect 30558 20476 30564 20528
rect 30616 20516 30622 20528
rect 30616 20488 31064 20516
rect 30616 20476 30622 20488
rect 30009 20451 30067 20457
rect 30009 20417 30021 20451
rect 30055 20417 30067 20451
rect 30009 20411 30067 20417
rect 30285 20451 30343 20457
rect 30285 20417 30297 20451
rect 30331 20417 30343 20451
rect 30285 20411 30343 20417
rect 30929 20451 30987 20457
rect 30929 20417 30941 20451
rect 30975 20417 30987 20451
rect 30929 20411 30987 20417
rect 27801 20383 27859 20389
rect 27801 20380 27813 20383
rect 27764 20352 27813 20380
rect 27764 20340 27770 20352
rect 27801 20349 27813 20352
rect 27847 20349 27859 20383
rect 27801 20343 27859 20349
rect 28997 20383 29055 20389
rect 28997 20349 29009 20383
rect 29043 20349 29055 20383
rect 28997 20343 29055 20349
rect 29273 20383 29331 20389
rect 29273 20349 29285 20383
rect 29319 20349 29331 20383
rect 29273 20343 29331 20349
rect 17129 20275 17187 20281
rect 18892 20284 20208 20312
rect 12253 20247 12311 20253
rect 12253 20244 12265 20247
rect 11164 20216 12265 20244
rect 12253 20213 12265 20216
rect 12299 20213 12311 20247
rect 12253 20207 12311 20213
rect 12342 20204 12348 20256
rect 12400 20244 12406 20256
rect 14734 20244 14740 20256
rect 12400 20216 14740 20244
rect 12400 20204 12406 20216
rect 14734 20204 14740 20216
rect 14792 20204 14798 20256
rect 15470 20204 15476 20256
rect 15528 20244 15534 20256
rect 15749 20247 15807 20253
rect 15749 20244 15761 20247
rect 15528 20216 15761 20244
rect 15528 20204 15534 20216
rect 15749 20213 15761 20216
rect 15795 20213 15807 20247
rect 15749 20207 15807 20213
rect 16669 20247 16727 20253
rect 16669 20213 16681 20247
rect 16715 20244 16727 20247
rect 16850 20244 16856 20256
rect 16715 20216 16856 20244
rect 16715 20213 16727 20216
rect 16669 20207 16727 20213
rect 16850 20204 16856 20216
rect 16908 20204 16914 20256
rect 17865 20247 17923 20253
rect 17865 20213 17877 20247
rect 17911 20244 17923 20247
rect 18892 20244 18920 20284
rect 20254 20272 20260 20324
rect 20312 20312 20318 20324
rect 21177 20315 21235 20321
rect 21177 20312 21189 20315
rect 20312 20284 21189 20312
rect 20312 20272 20318 20284
rect 21177 20281 21189 20284
rect 21223 20281 21235 20315
rect 21177 20275 21235 20281
rect 21910 20272 21916 20324
rect 21968 20312 21974 20324
rect 22554 20312 22560 20324
rect 21968 20284 22560 20312
rect 21968 20272 21974 20284
rect 22554 20272 22560 20284
rect 22612 20272 22618 20324
rect 23014 20272 23020 20324
rect 23072 20312 23078 20324
rect 24854 20312 24860 20324
rect 23072 20284 24860 20312
rect 23072 20272 23078 20284
rect 24854 20272 24860 20284
rect 24912 20272 24918 20324
rect 27614 20272 27620 20324
rect 27672 20312 27678 20324
rect 28442 20312 28448 20324
rect 27672 20284 28448 20312
rect 27672 20272 27678 20284
rect 28442 20272 28448 20284
rect 28500 20312 28506 20324
rect 29012 20312 29040 20343
rect 28500 20284 29040 20312
rect 28500 20272 28506 20284
rect 29086 20272 29092 20324
rect 29144 20312 29150 20324
rect 29288 20312 29316 20343
rect 29362 20340 29368 20392
rect 29420 20380 29426 20392
rect 30024 20380 30052 20411
rect 30834 20380 30840 20392
rect 29420 20352 30052 20380
rect 30116 20352 30840 20380
rect 29420 20340 29426 20352
rect 30116 20312 30144 20352
rect 30834 20340 30840 20352
rect 30892 20340 30898 20392
rect 29144 20284 30144 20312
rect 29144 20272 29150 20284
rect 30190 20272 30196 20324
rect 30248 20312 30254 20324
rect 30944 20312 30972 20411
rect 30248 20284 30972 20312
rect 31036 20380 31064 20488
rect 31205 20383 31263 20389
rect 31205 20380 31217 20383
rect 31036 20352 31217 20380
rect 30248 20272 30254 20284
rect 17911 20216 18920 20244
rect 19337 20247 19395 20253
rect 17911 20213 17923 20216
rect 17865 20207 17923 20213
rect 19337 20213 19349 20247
rect 19383 20244 19395 20247
rect 19429 20247 19487 20253
rect 19429 20244 19441 20247
rect 19383 20216 19441 20244
rect 19383 20213 19395 20216
rect 19337 20207 19395 20213
rect 19429 20213 19441 20216
rect 19475 20213 19487 20247
rect 19429 20207 19487 20213
rect 20070 20204 20076 20256
rect 20128 20244 20134 20256
rect 20622 20244 20628 20256
rect 20128 20216 20628 20244
rect 20128 20204 20134 20216
rect 20622 20204 20628 20216
rect 20680 20204 20686 20256
rect 21821 20247 21879 20253
rect 21821 20213 21833 20247
rect 21867 20244 21879 20247
rect 22002 20244 22008 20256
rect 21867 20216 22008 20244
rect 21867 20213 21879 20216
rect 21821 20207 21879 20213
rect 22002 20204 22008 20216
rect 22060 20204 22066 20256
rect 22278 20204 22284 20256
rect 22336 20244 22342 20256
rect 22462 20244 22468 20256
rect 22336 20216 22468 20244
rect 22336 20204 22342 20216
rect 22462 20204 22468 20216
rect 22520 20204 22526 20256
rect 23382 20204 23388 20256
rect 23440 20244 23446 20256
rect 23477 20247 23535 20253
rect 23477 20244 23489 20247
rect 23440 20216 23489 20244
rect 23440 20204 23446 20216
rect 23477 20213 23489 20216
rect 23523 20213 23535 20247
rect 23477 20207 23535 20213
rect 24302 20204 24308 20256
rect 24360 20244 24366 20256
rect 24670 20244 24676 20256
rect 24360 20216 24676 20244
rect 24360 20204 24366 20216
rect 24670 20204 24676 20216
rect 24728 20204 24734 20256
rect 25130 20204 25136 20256
rect 25188 20244 25194 20256
rect 25501 20247 25559 20253
rect 25501 20244 25513 20247
rect 25188 20216 25513 20244
rect 25188 20204 25194 20216
rect 25501 20213 25513 20216
rect 25547 20213 25559 20247
rect 25501 20207 25559 20213
rect 25961 20247 26019 20253
rect 25961 20213 25973 20247
rect 26007 20244 26019 20247
rect 26050 20244 26056 20256
rect 26007 20216 26056 20244
rect 26007 20213 26019 20216
rect 25961 20207 26019 20213
rect 26050 20204 26056 20216
rect 26108 20204 26114 20256
rect 26326 20244 26332 20256
rect 26287 20216 26332 20244
rect 26326 20204 26332 20216
rect 26384 20204 26390 20256
rect 28810 20244 28816 20256
rect 28771 20216 28816 20244
rect 28810 20204 28816 20216
rect 28868 20204 28874 20256
rect 29454 20204 29460 20256
rect 29512 20244 29518 20256
rect 30282 20244 30288 20256
rect 29512 20216 30288 20244
rect 29512 20204 29518 20216
rect 30282 20204 30288 20216
rect 30340 20204 30346 20256
rect 30742 20244 30748 20256
rect 30703 20216 30748 20244
rect 30742 20204 30748 20216
rect 30800 20204 30806 20256
rect 30834 20204 30840 20256
rect 30892 20244 30898 20256
rect 31036 20244 31064 20352
rect 31205 20349 31217 20352
rect 31251 20349 31263 20383
rect 31205 20343 31263 20349
rect 30892 20216 31064 20244
rect 31113 20247 31171 20253
rect 30892 20204 30898 20216
rect 31113 20213 31125 20247
rect 31159 20244 31171 20247
rect 31202 20244 31208 20256
rect 31159 20216 31208 20244
rect 31159 20213 31171 20216
rect 31113 20207 31171 20213
rect 31202 20204 31208 20216
rect 31260 20204 31266 20256
rect 1104 20154 32016 20176
rect 1104 20102 2136 20154
rect 2188 20102 12440 20154
rect 12492 20102 22744 20154
rect 22796 20102 32016 20154
rect 1104 20080 32016 20102
rect 2038 20000 2044 20052
rect 2096 20040 2102 20052
rect 2133 20043 2191 20049
rect 2133 20040 2145 20043
rect 2096 20012 2145 20040
rect 2096 20000 2102 20012
rect 2133 20009 2145 20012
rect 2179 20009 2191 20043
rect 5166 20040 5172 20052
rect 2133 20003 2191 20009
rect 2746 20012 4752 20040
rect 5127 20012 5172 20040
rect 1581 19975 1639 19981
rect 1581 19941 1593 19975
rect 1627 19972 1639 19975
rect 2746 19972 2774 20012
rect 1627 19944 2774 19972
rect 4724 19972 4752 20012
rect 5166 20000 5172 20012
rect 5224 20000 5230 20052
rect 5994 20040 6000 20052
rect 5276 20012 6000 20040
rect 5276 19972 5304 20012
rect 5994 20000 6000 20012
rect 6052 20000 6058 20052
rect 6362 20000 6368 20052
rect 6420 20040 6426 20052
rect 7006 20040 7012 20052
rect 6420 20012 6914 20040
rect 6967 20012 7012 20040
rect 6420 20000 6426 20012
rect 4724 19944 5304 19972
rect 6886 19972 6914 20012
rect 7006 20000 7012 20012
rect 7064 20000 7070 20052
rect 8754 20040 8760 20052
rect 7576 20012 8760 20040
rect 7576 19972 7604 20012
rect 8754 20000 8760 20012
rect 8812 20000 8818 20052
rect 8846 20000 8852 20052
rect 8904 20040 8910 20052
rect 13633 20043 13691 20049
rect 13633 20040 13645 20043
rect 8904 20012 13645 20040
rect 8904 20000 8910 20012
rect 13633 20009 13645 20012
rect 13679 20009 13691 20043
rect 15654 20040 15660 20052
rect 13633 20003 13691 20009
rect 13740 20012 15660 20040
rect 6886 19944 7604 19972
rect 7653 19975 7711 19981
rect 1627 19941 1639 19944
rect 1581 19935 1639 19941
rect 7653 19941 7665 19975
rect 7699 19972 7711 19975
rect 8662 19972 8668 19984
rect 7699 19944 8668 19972
rect 7699 19941 7711 19944
rect 7653 19935 7711 19941
rect 8662 19932 8668 19944
rect 8720 19932 8726 19984
rect 9306 19932 9312 19984
rect 9364 19972 9370 19984
rect 9401 19975 9459 19981
rect 9401 19972 9413 19975
rect 9364 19944 9413 19972
rect 9364 19932 9370 19944
rect 9401 19941 9413 19944
rect 9447 19941 9459 19975
rect 9401 19935 9459 19941
rect 9646 19944 10180 19972
rect 3510 19904 3516 19916
rect 2608 19876 3516 19904
rect 1302 19796 1308 19848
rect 1360 19836 1366 19848
rect 2608 19845 2636 19876
rect 3510 19864 3516 19876
rect 3568 19864 3574 19916
rect 5626 19904 5632 19916
rect 5587 19876 5632 19904
rect 5626 19864 5632 19876
rect 5684 19864 5690 19916
rect 8297 19907 8355 19913
rect 8297 19873 8309 19907
rect 8343 19904 8355 19907
rect 8386 19904 8392 19916
rect 8343 19876 8392 19904
rect 8343 19873 8355 19876
rect 8297 19867 8355 19873
rect 8386 19864 8392 19876
rect 8444 19864 8450 19916
rect 9646 19904 9674 19944
rect 8588 19876 9674 19904
rect 10152 19904 10180 19944
rect 10686 19932 10692 19984
rect 10744 19972 10750 19984
rect 11974 19972 11980 19984
rect 10744 19944 11980 19972
rect 10744 19932 10750 19944
rect 11974 19932 11980 19944
rect 12032 19932 12038 19984
rect 13740 19972 13768 20012
rect 15654 20000 15660 20012
rect 15712 20000 15718 20052
rect 17405 20043 17463 20049
rect 17405 20009 17417 20043
rect 17451 20040 17463 20043
rect 17773 20043 17831 20049
rect 17451 20012 17724 20040
rect 17451 20009 17463 20012
rect 17405 20003 17463 20009
rect 12084 19944 13768 19972
rect 10410 19904 10416 19916
rect 10152 19876 10416 19904
rect 1397 19839 1455 19845
rect 1397 19836 1409 19839
rect 1360 19808 1409 19836
rect 1360 19796 1366 19808
rect 1397 19805 1409 19808
rect 1443 19805 1455 19839
rect 1397 19799 1455 19805
rect 2317 19839 2375 19845
rect 2317 19805 2329 19839
rect 2363 19805 2375 19839
rect 2317 19799 2375 19805
rect 2593 19839 2651 19845
rect 2593 19805 2605 19839
rect 2639 19805 2651 19839
rect 2593 19799 2651 19805
rect 2777 19839 2835 19845
rect 2777 19805 2789 19839
rect 2823 19836 2835 19839
rect 2866 19836 2872 19848
rect 2823 19808 2872 19836
rect 2823 19805 2835 19808
rect 2777 19799 2835 19805
rect 1118 19728 1124 19780
rect 1176 19768 1182 19780
rect 1670 19768 1676 19780
rect 1176 19740 1676 19768
rect 1176 19728 1182 19740
rect 1670 19728 1676 19740
rect 1728 19728 1734 19780
rect 937 19703 995 19709
rect 937 19669 949 19703
rect 983 19700 995 19703
rect 1578 19700 1584 19712
rect 983 19672 1584 19700
rect 983 19669 995 19672
rect 937 19663 995 19669
rect 1578 19660 1584 19672
rect 1636 19660 1642 19712
rect 2332 19700 2360 19799
rect 2866 19796 2872 19808
rect 2924 19796 2930 19848
rect 3789 19839 3847 19845
rect 3789 19805 3801 19839
rect 3835 19836 3847 19839
rect 3878 19836 3884 19848
rect 3835 19808 3884 19836
rect 3835 19805 3847 19808
rect 3789 19799 3847 19805
rect 3878 19796 3884 19808
rect 3936 19796 3942 19848
rect 3050 19728 3056 19780
rect 3108 19768 3114 19780
rect 4034 19771 4092 19777
rect 4034 19768 4046 19771
rect 3108 19740 4046 19768
rect 3108 19728 3114 19740
rect 4034 19737 4046 19740
rect 4080 19737 4092 19771
rect 4034 19731 4092 19737
rect 5896 19771 5954 19777
rect 5896 19737 5908 19771
rect 5942 19768 5954 19771
rect 6362 19768 6368 19780
rect 5942 19740 6368 19768
rect 5942 19737 5954 19740
rect 5896 19731 5954 19737
rect 6362 19728 6368 19740
rect 6420 19728 6426 19780
rect 8588 19768 8616 19876
rect 10410 19864 10416 19876
rect 10468 19864 10474 19916
rect 11701 19907 11759 19913
rect 11701 19904 11713 19907
rect 10612 19876 11713 19904
rect 9122 19796 9128 19848
rect 9180 19836 9186 19848
rect 9401 19839 9459 19845
rect 9401 19836 9413 19839
rect 9180 19808 9413 19836
rect 9180 19796 9186 19808
rect 9401 19805 9413 19808
rect 9447 19805 9459 19839
rect 9950 19836 9956 19848
rect 9911 19808 9956 19836
rect 9401 19799 9459 19805
rect 9950 19796 9956 19808
rect 10008 19796 10014 19848
rect 10045 19839 10103 19845
rect 10045 19805 10057 19839
rect 10091 19805 10103 19839
rect 10502 19836 10508 19848
rect 10463 19808 10508 19836
rect 10045 19799 10103 19805
rect 6472 19740 8616 19768
rect 3602 19700 3608 19712
rect 2332 19672 3608 19700
rect 3602 19660 3608 19672
rect 3660 19660 3666 19712
rect 4338 19660 4344 19712
rect 4396 19700 4402 19712
rect 6472 19700 6500 19740
rect 9766 19728 9772 19780
rect 9824 19768 9830 19780
rect 10060 19768 10088 19799
rect 10502 19796 10508 19808
rect 10560 19796 10566 19848
rect 9824 19740 10088 19768
rect 9824 19728 9830 19740
rect 10134 19728 10140 19780
rect 10192 19768 10198 19780
rect 10612 19768 10640 19876
rect 11701 19873 11713 19876
rect 11747 19873 11759 19907
rect 12084 19904 12112 19944
rect 14274 19932 14280 19984
rect 14332 19972 14338 19984
rect 15105 19975 15163 19981
rect 15105 19972 15117 19975
rect 14332 19944 15117 19972
rect 14332 19932 14338 19944
rect 15105 19941 15117 19944
rect 15151 19941 15163 19975
rect 17696 19972 17724 20012
rect 17773 20009 17785 20043
rect 17819 20040 17831 20043
rect 18046 20040 18052 20052
rect 17819 20012 18052 20040
rect 17819 20009 17831 20012
rect 17773 20003 17831 20009
rect 18046 20000 18052 20012
rect 18104 20000 18110 20052
rect 18230 20000 18236 20052
rect 18288 20040 18294 20052
rect 19613 20043 19671 20049
rect 19613 20040 19625 20043
rect 18288 20012 19625 20040
rect 18288 20000 18294 20012
rect 19613 20009 19625 20012
rect 19659 20009 19671 20043
rect 19613 20003 19671 20009
rect 19978 20000 19984 20052
rect 20036 20040 20042 20052
rect 21266 20040 21272 20052
rect 20036 20012 21272 20040
rect 20036 20000 20042 20012
rect 21266 20000 21272 20012
rect 21324 20000 21330 20052
rect 21634 20000 21640 20052
rect 21692 20040 21698 20052
rect 22278 20040 22284 20052
rect 21692 20012 22284 20040
rect 21692 20000 21698 20012
rect 22278 20000 22284 20012
rect 22336 20040 22342 20052
rect 22336 20012 23428 20040
rect 22336 20000 22342 20012
rect 18322 19972 18328 19984
rect 17696 19944 18328 19972
rect 15105 19935 15163 19941
rect 18322 19932 18328 19944
rect 18380 19932 18386 19984
rect 18598 19932 18604 19984
rect 18656 19972 18662 19984
rect 19242 19972 19248 19984
rect 18656 19944 19248 19972
rect 18656 19932 18662 19944
rect 19242 19932 19248 19944
rect 19300 19972 19306 19984
rect 21545 19975 21603 19981
rect 21545 19972 21557 19975
rect 19300 19944 21557 19972
rect 19300 19932 19306 19944
rect 21545 19941 21557 19944
rect 21591 19972 21603 19975
rect 21910 19972 21916 19984
rect 21591 19944 21916 19972
rect 21591 19941 21603 19944
rect 21545 19935 21603 19941
rect 21910 19932 21916 19944
rect 21968 19972 21974 19984
rect 23400 19972 23428 20012
rect 23474 20000 23480 20052
rect 23532 20040 23538 20052
rect 23845 20043 23903 20049
rect 23845 20040 23857 20043
rect 23532 20012 23857 20040
rect 23532 20000 23538 20012
rect 23845 20009 23857 20012
rect 23891 20009 23903 20043
rect 23845 20003 23903 20009
rect 24213 20043 24271 20049
rect 24213 20009 24225 20043
rect 24259 20040 24271 20043
rect 24762 20040 24768 20052
rect 24259 20012 24624 20040
rect 24723 20012 24768 20040
rect 24259 20009 24271 20012
rect 24213 20003 24271 20009
rect 24596 19972 24624 20012
rect 24762 20000 24768 20012
rect 24820 20000 24826 20052
rect 25041 20043 25099 20049
rect 25041 20009 25053 20043
rect 25087 20040 25099 20043
rect 26234 20040 26240 20052
rect 25087 20012 26240 20040
rect 25087 20009 25099 20012
rect 25041 20003 25099 20009
rect 26234 20000 26240 20012
rect 26292 20040 26298 20052
rect 27249 20043 27307 20049
rect 26292 20012 27200 20040
rect 26292 20000 26298 20012
rect 25222 19972 25228 19984
rect 21968 19944 22094 19972
rect 23400 19944 24512 19972
rect 24596 19944 25228 19972
rect 21968 19932 21974 19944
rect 14093 19907 14151 19913
rect 14093 19904 14105 19907
rect 11701 19867 11759 19873
rect 11788 19876 12112 19904
rect 12912 19876 14105 19904
rect 11238 19836 11244 19848
rect 11199 19808 11244 19836
rect 11238 19796 11244 19808
rect 11296 19796 11302 19848
rect 11514 19796 11520 19848
rect 11572 19836 11578 19848
rect 11788 19836 11816 19876
rect 11572 19808 11816 19836
rect 11885 19839 11943 19845
rect 11572 19796 11578 19808
rect 11885 19805 11897 19839
rect 11931 19805 11943 19839
rect 11885 19799 11943 19805
rect 12069 19839 12127 19845
rect 12069 19805 12081 19839
rect 12115 19836 12127 19839
rect 12342 19836 12348 19848
rect 12115 19808 12348 19836
rect 12115 19805 12127 19808
rect 12069 19799 12127 19805
rect 10192 19740 10640 19768
rect 10192 19728 10198 19740
rect 11054 19728 11060 19780
rect 11112 19768 11118 19780
rect 11900 19768 11928 19799
rect 12342 19796 12348 19808
rect 12400 19796 12406 19848
rect 12912 19845 12940 19876
rect 14093 19873 14105 19876
rect 14139 19873 14151 19907
rect 14093 19867 14151 19873
rect 14182 19864 14188 19916
rect 14240 19904 14246 19916
rect 15749 19907 15807 19913
rect 14240 19876 15608 19904
rect 14240 19864 14246 19876
rect 12897 19839 12955 19845
rect 12897 19805 12909 19839
rect 12943 19805 12955 19839
rect 13078 19836 13084 19848
rect 13039 19808 13084 19836
rect 12897 19799 12955 19805
rect 13078 19796 13084 19808
rect 13136 19796 13142 19848
rect 13173 19839 13231 19845
rect 13173 19805 13185 19839
rect 13219 19805 13231 19839
rect 13173 19799 13231 19805
rect 13299 19839 13357 19845
rect 13299 19805 13311 19839
rect 13345 19836 13357 19839
rect 13541 19839 13599 19845
rect 13345 19808 13492 19836
rect 13345 19805 13357 19808
rect 13299 19799 13357 19805
rect 11112 19740 11928 19768
rect 11112 19728 11118 19740
rect 11974 19728 11980 19780
rect 12032 19768 12038 19780
rect 12032 19740 12198 19768
rect 12032 19728 12038 19740
rect 4396 19672 6500 19700
rect 4396 19660 4402 19672
rect 7650 19660 7656 19712
rect 7708 19700 7714 19712
rect 8021 19703 8079 19709
rect 8021 19700 8033 19703
rect 7708 19672 8033 19700
rect 7708 19660 7714 19672
rect 8021 19669 8033 19672
rect 8067 19669 8079 19703
rect 8021 19663 8079 19669
rect 8110 19660 8116 19712
rect 8168 19700 8174 19712
rect 8168 19672 8213 19700
rect 8168 19660 8174 19672
rect 8570 19660 8576 19712
rect 8628 19700 8634 19712
rect 12066 19700 12072 19712
rect 8628 19672 12072 19700
rect 8628 19660 8634 19672
rect 12066 19660 12072 19672
rect 12124 19660 12130 19712
rect 12170 19700 12198 19740
rect 12986 19728 12992 19780
rect 13044 19768 13050 19780
rect 13188 19768 13216 19799
rect 13044 19740 13216 19768
rect 13464 19768 13492 19808
rect 13541 19805 13553 19839
rect 13587 19836 13599 19839
rect 13633 19839 13691 19845
rect 13633 19836 13645 19839
rect 13587 19808 13645 19836
rect 13587 19805 13599 19808
rect 13541 19799 13599 19805
rect 13633 19805 13645 19808
rect 13679 19805 13691 19839
rect 13633 19799 13691 19805
rect 13998 19796 14004 19848
rect 14056 19836 14062 19848
rect 14277 19839 14335 19845
rect 14277 19836 14289 19839
rect 14056 19808 14289 19836
rect 14056 19796 14062 19808
rect 14277 19805 14289 19808
rect 14323 19836 14335 19839
rect 14366 19836 14372 19848
rect 14323 19808 14372 19836
rect 14323 19805 14335 19808
rect 14277 19799 14335 19805
rect 14366 19796 14372 19808
rect 14424 19796 14430 19848
rect 14458 19796 14464 19848
rect 14516 19836 14522 19848
rect 14553 19839 14611 19845
rect 14553 19836 14565 19839
rect 14516 19808 14565 19836
rect 14516 19796 14522 19808
rect 14553 19805 14565 19808
rect 14599 19805 14611 19839
rect 14553 19799 14611 19805
rect 14918 19796 14924 19848
rect 14976 19836 14982 19848
rect 15286 19836 15292 19848
rect 14976 19808 15292 19836
rect 14976 19796 14982 19808
rect 15286 19796 15292 19808
rect 15344 19796 15350 19848
rect 15470 19836 15476 19848
rect 15431 19808 15476 19836
rect 15470 19796 15476 19808
rect 15528 19796 15534 19848
rect 15580 19836 15608 19876
rect 15749 19873 15761 19907
rect 15795 19904 15807 19907
rect 16022 19904 16028 19916
rect 15795 19876 16028 19904
rect 15795 19873 15807 19876
rect 15749 19867 15807 19873
rect 16022 19864 16028 19876
rect 16080 19864 16086 19916
rect 16850 19904 16856 19916
rect 16811 19876 16856 19904
rect 16850 19864 16856 19876
rect 16908 19864 16914 19916
rect 17218 19904 17224 19916
rect 17179 19876 17224 19904
rect 17218 19864 17224 19876
rect 17276 19864 17282 19916
rect 17494 19864 17500 19916
rect 17552 19904 17558 19916
rect 17552 19876 17908 19904
rect 17552 19864 17558 19876
rect 17880 19848 17908 19876
rect 18046 19864 18052 19916
rect 18104 19904 18110 19916
rect 18874 19904 18880 19916
rect 18104 19876 18880 19904
rect 18104 19864 18110 19876
rect 18874 19864 18880 19876
rect 18932 19864 18938 19916
rect 18966 19864 18972 19916
rect 19024 19904 19030 19916
rect 19150 19904 19156 19916
rect 19024 19876 19156 19904
rect 19024 19864 19030 19876
rect 19150 19864 19156 19876
rect 19208 19864 19214 19916
rect 22066 19904 22094 19944
rect 22465 19907 22523 19913
rect 22465 19904 22477 19907
rect 22066 19876 22477 19904
rect 22465 19873 22477 19876
rect 22511 19873 22523 19907
rect 22465 19867 22523 19873
rect 15580 19830 17639 19836
rect 17770 19830 17776 19848
rect 15580 19808 17776 19830
rect 17611 19802 17776 19808
rect 17770 19796 17776 19802
rect 17828 19796 17834 19848
rect 17862 19796 17868 19848
rect 17920 19836 17926 19848
rect 17957 19839 18015 19845
rect 17957 19836 17969 19839
rect 17920 19808 17969 19836
rect 17920 19796 17926 19808
rect 17957 19805 17969 19808
rect 18003 19805 18015 19839
rect 19978 19836 19984 19848
rect 17957 19799 18015 19805
rect 18156 19808 19984 19836
rect 14090 19768 14096 19780
rect 13464 19740 14096 19768
rect 13044 19728 13050 19740
rect 14090 19728 14096 19740
rect 14148 19768 14154 19780
rect 14148 19740 14504 19768
rect 14148 19728 14154 19740
rect 14182 19700 14188 19712
rect 12170 19672 14188 19700
rect 14182 19660 14188 19672
rect 14240 19660 14246 19712
rect 14476 19709 14504 19740
rect 15102 19728 15108 19780
rect 15160 19768 15166 19780
rect 18156 19777 18184 19808
rect 19978 19796 19984 19808
rect 20036 19796 20042 19848
rect 20346 19796 20352 19848
rect 20404 19836 20410 19848
rect 20404 19808 20760 19836
rect 20404 19796 20410 19808
rect 18141 19771 18199 19777
rect 18141 19768 18153 19771
rect 15160 19740 17816 19768
rect 15160 19728 15166 19740
rect 14461 19703 14519 19709
rect 14461 19669 14473 19703
rect 14507 19700 14519 19703
rect 14734 19700 14740 19712
rect 14507 19672 14740 19700
rect 14507 19669 14519 19672
rect 14461 19663 14519 19669
rect 14734 19660 14740 19672
rect 14792 19660 14798 19712
rect 15562 19660 15568 19712
rect 15620 19700 15626 19712
rect 17037 19703 17095 19709
rect 15620 19672 15665 19700
rect 15620 19660 15626 19672
rect 17037 19669 17049 19703
rect 17083 19700 17095 19703
rect 17681 19703 17739 19709
rect 17681 19700 17693 19703
rect 17083 19672 17693 19700
rect 17083 19669 17095 19672
rect 17037 19663 17095 19669
rect 17681 19669 17693 19672
rect 17727 19669 17739 19703
rect 17788 19700 17816 19740
rect 17984 19740 18153 19768
rect 17984 19700 18012 19740
rect 18141 19737 18153 19740
rect 18187 19737 18199 19771
rect 18141 19731 18199 19737
rect 19429 19771 19487 19777
rect 19429 19737 19441 19771
rect 19475 19768 19487 19771
rect 20070 19768 20076 19780
rect 19475 19740 20076 19768
rect 19475 19737 19487 19740
rect 19429 19731 19487 19737
rect 20070 19728 20076 19740
rect 20128 19728 20134 19780
rect 20257 19771 20315 19777
rect 20257 19737 20269 19771
rect 20303 19768 20315 19771
rect 20622 19768 20628 19780
rect 20303 19740 20628 19768
rect 20303 19737 20315 19740
rect 20257 19731 20315 19737
rect 20622 19728 20628 19740
rect 20680 19728 20686 19780
rect 20732 19768 20760 19808
rect 22002 19796 22008 19848
rect 22060 19836 22066 19848
rect 22721 19839 22779 19845
rect 22721 19836 22733 19839
rect 22060 19808 22733 19836
rect 22060 19796 22066 19808
rect 22721 19805 22733 19808
rect 22767 19805 22779 19839
rect 22721 19799 22779 19805
rect 24213 19839 24271 19845
rect 24213 19805 24225 19839
rect 24259 19836 24271 19839
rect 24397 19839 24455 19845
rect 24397 19836 24409 19839
rect 24259 19808 24409 19836
rect 24259 19805 24271 19808
rect 24213 19799 24271 19805
rect 24397 19805 24409 19808
rect 24443 19805 24455 19839
rect 24484 19836 24512 19944
rect 25222 19932 25228 19944
rect 25280 19932 25286 19984
rect 27172 19972 27200 20012
rect 27249 20009 27261 20043
rect 27295 20040 27307 20043
rect 27798 20040 27804 20052
rect 27295 20012 27804 20040
rect 27295 20009 27307 20012
rect 27249 20003 27307 20009
rect 27798 20000 27804 20012
rect 27856 20000 27862 20052
rect 28258 20000 28264 20052
rect 28316 20040 28322 20052
rect 28353 20043 28411 20049
rect 28353 20040 28365 20043
rect 28316 20012 28365 20040
rect 28316 20000 28322 20012
rect 28353 20009 28365 20012
rect 28399 20009 28411 20043
rect 29454 20040 29460 20052
rect 28353 20003 28411 20009
rect 28552 20012 29460 20040
rect 27430 19972 27436 19984
rect 27172 19944 27436 19972
rect 27430 19932 27436 19944
rect 27488 19932 27494 19984
rect 27522 19932 27528 19984
rect 27580 19972 27586 19984
rect 27709 19975 27767 19981
rect 27709 19972 27721 19975
rect 27580 19944 27721 19972
rect 27580 19932 27586 19944
rect 27709 19941 27721 19944
rect 27755 19941 27767 19975
rect 27709 19935 27767 19941
rect 24854 19864 24860 19916
rect 24912 19904 24918 19916
rect 24912 19876 25452 19904
rect 24912 19864 24918 19876
rect 25424 19845 25452 19876
rect 27614 19864 27620 19916
rect 27672 19864 27678 19916
rect 27724 19904 27752 19935
rect 28552 19904 28580 20012
rect 29454 20000 29460 20012
rect 29512 20000 29518 20052
rect 29546 20000 29552 20052
rect 29604 20040 29610 20052
rect 30558 20040 30564 20052
rect 29604 20012 30564 20040
rect 29604 20000 29610 20012
rect 30558 20000 30564 20012
rect 30616 20000 30622 20052
rect 28902 19972 28908 19984
rect 27724 19876 28580 19904
rect 24581 19839 24639 19845
rect 24581 19836 24593 19839
rect 24484 19808 24593 19836
rect 24397 19799 24455 19805
rect 24581 19805 24593 19808
rect 24627 19805 24639 19839
rect 24581 19799 24639 19805
rect 25041 19839 25099 19845
rect 25041 19805 25053 19839
rect 25087 19836 25099 19839
rect 25225 19839 25283 19845
rect 25225 19836 25237 19839
rect 25087 19808 25237 19836
rect 25087 19805 25099 19808
rect 25041 19799 25099 19805
rect 25225 19805 25237 19808
rect 25271 19805 25283 19839
rect 25225 19799 25283 19805
rect 25409 19839 25467 19845
rect 25409 19805 25421 19839
rect 25455 19805 25467 19839
rect 25409 19799 25467 19805
rect 25774 19796 25780 19848
rect 25832 19836 25838 19848
rect 26142 19845 26148 19848
rect 25869 19839 25927 19845
rect 25869 19836 25881 19839
rect 25832 19808 25881 19836
rect 25832 19796 25838 19808
rect 25869 19805 25881 19808
rect 25915 19805 25927 19839
rect 26136 19836 26148 19845
rect 26103 19808 26148 19836
rect 25869 19799 25927 19805
rect 26136 19799 26148 19808
rect 26142 19796 26148 19799
rect 26200 19796 26206 19848
rect 27632 19836 27660 19864
rect 28552 19845 28580 19876
rect 28828 19944 28908 19972
rect 27709 19839 27767 19845
rect 27709 19836 27721 19839
rect 27586 19808 27721 19836
rect 22094 19768 22100 19780
rect 20732 19740 22100 19768
rect 22094 19728 22100 19740
rect 22152 19728 22158 19780
rect 24670 19768 24676 19780
rect 23400 19740 24676 19768
rect 17788 19672 18012 19700
rect 17681 19663 17739 19669
rect 18598 19660 18604 19712
rect 18656 19700 18662 19712
rect 19629 19703 19687 19709
rect 19629 19700 19641 19703
rect 18656 19672 19641 19700
rect 18656 19660 18662 19672
rect 19629 19669 19641 19672
rect 19675 19669 19687 19703
rect 19629 19663 19687 19669
rect 19797 19703 19855 19709
rect 19797 19669 19809 19703
rect 19843 19700 19855 19703
rect 23400 19700 23428 19740
rect 24670 19728 24676 19740
rect 24728 19728 24734 19780
rect 25130 19728 25136 19780
rect 25188 19768 25194 19780
rect 27586 19768 27614 19808
rect 27709 19805 27721 19808
rect 27755 19805 27767 19839
rect 27893 19839 27951 19845
rect 27893 19836 27905 19839
rect 27709 19799 27767 19805
rect 27816 19808 27905 19836
rect 27816 19780 27844 19808
rect 27893 19805 27905 19808
rect 27939 19805 27951 19839
rect 27893 19799 27951 19805
rect 28537 19839 28595 19845
rect 28537 19805 28549 19839
rect 28583 19805 28595 19839
rect 28537 19799 28595 19805
rect 28629 19839 28687 19845
rect 28629 19805 28641 19839
rect 28675 19836 28687 19839
rect 28718 19836 28724 19848
rect 28675 19808 28724 19836
rect 28675 19805 28687 19808
rect 28629 19799 28687 19805
rect 28718 19796 28724 19808
rect 28776 19796 28782 19848
rect 28828 19845 28856 19944
rect 28902 19932 28908 19944
rect 28960 19932 28966 19984
rect 29914 19904 29920 19916
rect 29875 19876 29920 19904
rect 29914 19864 29920 19876
rect 29972 19864 29978 19916
rect 28813 19839 28871 19845
rect 28813 19805 28825 19839
rect 28859 19805 28871 19839
rect 28813 19799 28871 19805
rect 28902 19796 28908 19848
rect 28960 19836 28966 19848
rect 30184 19839 30242 19845
rect 28960 19808 29005 19836
rect 28960 19796 28966 19808
rect 30184 19805 30196 19839
rect 30230 19836 30242 19839
rect 30742 19836 30748 19848
rect 30230 19808 30748 19836
rect 30230 19805 30242 19808
rect 30184 19799 30242 19805
rect 30742 19796 30748 19808
rect 30800 19796 30806 19848
rect 25188 19740 27614 19768
rect 25188 19728 25194 19740
rect 27798 19728 27804 19780
rect 27856 19728 27862 19780
rect 28350 19728 28356 19780
rect 28408 19768 28414 19780
rect 30374 19768 30380 19780
rect 28408 19740 30380 19768
rect 28408 19728 28414 19740
rect 30374 19728 30380 19740
rect 30432 19768 30438 19780
rect 31202 19768 31208 19780
rect 30432 19740 31208 19768
rect 30432 19728 30438 19740
rect 31202 19728 31208 19740
rect 31260 19728 31266 19780
rect 19843 19672 23428 19700
rect 19843 19669 19855 19672
rect 19797 19663 19855 19669
rect 23474 19660 23480 19712
rect 23532 19700 23538 19712
rect 25317 19703 25375 19709
rect 25317 19700 25329 19703
rect 23532 19672 25329 19700
rect 23532 19660 23538 19672
rect 25317 19669 25329 19672
rect 25363 19669 25375 19703
rect 25317 19663 25375 19669
rect 28166 19660 28172 19712
rect 28224 19700 28230 19712
rect 29362 19700 29368 19712
rect 28224 19672 29368 19700
rect 28224 19660 28230 19672
rect 29362 19660 29368 19672
rect 29420 19660 29426 19712
rect 29822 19660 29828 19712
rect 29880 19700 29886 19712
rect 30558 19700 30564 19712
rect 29880 19672 30564 19700
rect 29880 19660 29886 19672
rect 30558 19660 30564 19672
rect 30616 19660 30622 19712
rect 31110 19660 31116 19712
rect 31168 19700 31174 19712
rect 31297 19703 31355 19709
rect 31297 19700 31309 19703
rect 31168 19672 31309 19700
rect 31168 19660 31174 19672
rect 31297 19669 31309 19672
rect 31343 19669 31355 19703
rect 31297 19663 31355 19669
rect 1104 19610 32016 19632
rect 1104 19558 7288 19610
rect 7340 19558 17592 19610
rect 17644 19558 27896 19610
rect 27948 19558 32016 19610
rect 1104 19536 32016 19558
rect 2774 19496 2780 19508
rect 1412 19468 2780 19496
rect 1412 19369 1440 19468
rect 2774 19456 2780 19468
rect 2832 19496 2838 19508
rect 3878 19496 3884 19508
rect 2832 19468 3884 19496
rect 2832 19456 2838 19468
rect 3878 19456 3884 19468
rect 3936 19456 3942 19508
rect 4338 19496 4344 19508
rect 4299 19468 4344 19496
rect 4338 19456 4344 19468
rect 4396 19456 4402 19508
rect 6086 19456 6092 19508
rect 6144 19496 6150 19508
rect 6822 19496 6828 19508
rect 6144 19468 6828 19496
rect 6144 19456 6150 19468
rect 6822 19456 6828 19468
rect 6880 19456 6886 19508
rect 7006 19496 7012 19508
rect 6967 19468 7012 19496
rect 7006 19456 7012 19468
rect 7064 19456 7070 19508
rect 7193 19499 7251 19505
rect 7193 19465 7205 19499
rect 7239 19496 7251 19499
rect 8202 19496 8208 19508
rect 7239 19468 8208 19496
rect 7239 19465 7251 19468
rect 7193 19459 7251 19465
rect 8202 19456 8208 19468
rect 8260 19456 8266 19508
rect 8754 19456 8760 19508
rect 8812 19496 8818 19508
rect 11974 19496 11980 19508
rect 8812 19468 10548 19496
rect 8812 19456 8818 19468
rect 1578 19388 1584 19440
rect 1636 19428 1642 19440
rect 1854 19428 1860 19440
rect 1636 19400 1860 19428
rect 1636 19388 1642 19400
rect 1854 19388 1860 19400
rect 1912 19388 1918 19440
rect 7558 19428 7564 19440
rect 4540 19400 7564 19428
rect 1670 19369 1676 19372
rect 1397 19363 1455 19369
rect 1397 19329 1409 19363
rect 1443 19329 1455 19363
rect 1397 19323 1455 19329
rect 1664 19323 1676 19369
rect 1728 19360 1734 19372
rect 1728 19332 1764 19360
rect 1670 19320 1676 19323
rect 1728 19320 1734 19332
rect 1946 19320 1952 19372
rect 2004 19360 2010 19372
rect 2682 19360 2688 19372
rect 2004 19332 2688 19360
rect 2004 19320 2010 19332
rect 2682 19320 2688 19332
rect 2740 19360 2746 19372
rect 3421 19363 3479 19369
rect 3421 19360 3433 19363
rect 2740 19332 3433 19360
rect 2740 19320 2746 19332
rect 3421 19329 3433 19332
rect 3467 19329 3479 19363
rect 3421 19323 3479 19329
rect 3510 19320 3516 19372
rect 3568 19360 3574 19372
rect 3697 19363 3755 19369
rect 3697 19360 3709 19363
rect 3568 19332 3709 19360
rect 3568 19320 3574 19332
rect 3697 19329 3709 19332
rect 3743 19329 3755 19363
rect 3697 19323 3755 19329
rect 3712 19292 3740 19323
rect 3786 19320 3792 19372
rect 3844 19360 3850 19372
rect 4540 19369 4568 19400
rect 7558 19388 7564 19400
rect 7616 19388 7622 19440
rect 8938 19428 8944 19440
rect 7668 19400 8944 19428
rect 3881 19363 3939 19369
rect 3881 19360 3893 19363
rect 3844 19332 3893 19360
rect 3844 19320 3850 19332
rect 3881 19329 3893 19332
rect 3927 19329 3939 19363
rect 3881 19323 3939 19329
rect 4525 19363 4583 19369
rect 4525 19329 4537 19363
rect 4571 19329 4583 19363
rect 4525 19323 4583 19329
rect 4985 19363 5043 19369
rect 4985 19329 4997 19363
rect 5031 19360 5043 19363
rect 5166 19360 5172 19372
rect 5031 19332 5172 19360
rect 5031 19329 5043 19332
rect 4985 19323 5043 19329
rect 5166 19320 5172 19332
rect 5224 19320 5230 19372
rect 5261 19363 5319 19369
rect 5261 19329 5273 19363
rect 5307 19329 5319 19363
rect 5261 19323 5319 19329
rect 3970 19292 3976 19304
rect 3712 19264 3976 19292
rect 3970 19252 3976 19264
rect 4028 19252 4034 19304
rect 4430 19252 4436 19304
rect 4488 19292 4494 19304
rect 5276 19292 5304 19323
rect 5626 19320 5632 19372
rect 5684 19360 5690 19372
rect 7668 19369 7696 19400
rect 8938 19388 8944 19400
rect 8996 19388 9002 19440
rect 7653 19363 7711 19369
rect 7653 19360 7665 19363
rect 5684 19332 7665 19360
rect 5684 19320 5690 19332
rect 7653 19329 7665 19332
rect 7699 19329 7711 19363
rect 7653 19323 7711 19329
rect 7920 19363 7978 19369
rect 7920 19329 7932 19363
rect 7966 19360 7978 19363
rect 7966 19332 8708 19360
rect 7966 19329 7978 19332
rect 7920 19323 7978 19329
rect 6638 19292 6644 19304
rect 4488 19264 6644 19292
rect 4488 19252 4494 19264
rect 6638 19252 6644 19264
rect 6696 19252 6702 19304
rect 8680 19292 8708 19332
rect 8754 19320 8760 19372
rect 8812 19360 8818 19372
rect 9493 19363 9551 19369
rect 9493 19360 9505 19363
rect 8812 19332 9505 19360
rect 8812 19320 8818 19332
rect 9493 19329 9505 19332
rect 9539 19329 9551 19363
rect 9493 19323 9551 19329
rect 9677 19363 9735 19369
rect 9677 19329 9689 19363
rect 9723 19360 9735 19363
rect 9950 19360 9956 19372
rect 9723 19332 9956 19360
rect 9723 19329 9735 19332
rect 9677 19323 9735 19329
rect 9950 19320 9956 19332
rect 10008 19320 10014 19372
rect 10520 19369 10548 19468
rect 11072 19468 11980 19496
rect 10778 19388 10784 19440
rect 10836 19428 10842 19440
rect 10873 19431 10931 19437
rect 10873 19428 10885 19431
rect 10836 19400 10885 19428
rect 10836 19388 10842 19400
rect 10873 19397 10885 19400
rect 10919 19397 10931 19431
rect 10873 19391 10931 19397
rect 10505 19363 10563 19369
rect 10505 19329 10517 19363
rect 10551 19360 10563 19363
rect 11072 19360 11100 19468
rect 11974 19456 11980 19468
rect 12032 19456 12038 19508
rect 12894 19496 12900 19508
rect 12855 19468 12900 19496
rect 12894 19456 12900 19468
rect 12952 19456 12958 19508
rect 13078 19456 13084 19508
rect 13136 19496 13142 19508
rect 13357 19499 13415 19505
rect 13357 19496 13369 19499
rect 13136 19468 13369 19496
rect 13136 19456 13142 19468
rect 13357 19465 13369 19468
rect 13403 19465 13415 19499
rect 13357 19459 13415 19465
rect 14277 19499 14335 19505
rect 14277 19465 14289 19499
rect 14323 19496 14335 19499
rect 14826 19496 14832 19508
rect 14323 19468 14832 19496
rect 14323 19465 14335 19468
rect 14277 19459 14335 19465
rect 14826 19456 14832 19468
rect 14884 19456 14890 19508
rect 15381 19499 15439 19505
rect 15381 19465 15393 19499
rect 15427 19496 15439 19499
rect 15562 19496 15568 19508
rect 15427 19468 15568 19496
rect 15427 19465 15439 19468
rect 15381 19459 15439 19465
rect 15562 19456 15568 19468
rect 15620 19456 15626 19508
rect 15746 19496 15752 19508
rect 15707 19468 15752 19496
rect 15746 19456 15752 19468
rect 15804 19456 15810 19508
rect 16482 19496 16488 19508
rect 16443 19468 16488 19496
rect 16482 19456 16488 19468
rect 16540 19456 16546 19508
rect 16853 19499 16911 19505
rect 16853 19465 16865 19499
rect 16899 19496 16911 19499
rect 16942 19496 16948 19508
rect 16899 19468 16948 19496
rect 16899 19465 16911 19468
rect 16853 19459 16911 19465
rect 16942 19456 16948 19468
rect 17000 19456 17006 19508
rect 17129 19499 17187 19505
rect 17129 19465 17141 19499
rect 17175 19496 17187 19499
rect 18233 19499 18291 19505
rect 18233 19496 18245 19499
rect 17175 19468 18245 19496
rect 17175 19465 17187 19468
rect 17129 19459 17187 19465
rect 18233 19465 18245 19468
rect 18279 19465 18291 19499
rect 18233 19459 18291 19465
rect 18322 19456 18328 19508
rect 18380 19496 18386 19508
rect 19153 19499 19211 19505
rect 19153 19496 19165 19499
rect 18380 19468 19165 19496
rect 18380 19456 18386 19468
rect 19153 19465 19165 19468
rect 19199 19496 19211 19499
rect 19610 19496 19616 19508
rect 19199 19468 19616 19496
rect 19199 19465 19211 19468
rect 19153 19459 19211 19465
rect 19610 19456 19616 19468
rect 19668 19456 19674 19508
rect 21818 19496 21824 19508
rect 21779 19468 21824 19496
rect 21818 19456 21824 19468
rect 21876 19456 21882 19508
rect 23201 19499 23259 19505
rect 23201 19465 23213 19499
rect 23247 19465 23259 19499
rect 23201 19459 23259 19465
rect 11606 19388 11612 19440
rect 11664 19428 11670 19440
rect 11762 19431 11820 19437
rect 11762 19428 11774 19431
rect 11664 19400 11774 19428
rect 11664 19388 11670 19400
rect 11762 19397 11774 19400
rect 11808 19397 11820 19431
rect 11762 19391 11820 19397
rect 12066 19388 12072 19440
rect 12124 19428 12130 19440
rect 18138 19428 18144 19440
rect 12124 19400 16804 19428
rect 12124 19388 12130 19400
rect 11330 19360 11336 19372
rect 10551 19358 10824 19360
rect 10980 19358 11100 19360
rect 10551 19332 11100 19358
rect 11164 19332 11336 19360
rect 10551 19329 10563 19332
rect 10796 19330 11008 19332
rect 10505 19323 10563 19329
rect 9585 19295 9643 19301
rect 9585 19292 9597 19295
rect 8680 19264 9597 19292
rect 9585 19261 9597 19264
rect 9631 19261 9643 19295
rect 10689 19295 10747 19301
rect 9585 19255 9643 19261
rect 9683 19264 10640 19292
rect 6454 19184 6460 19236
rect 6512 19224 6518 19236
rect 9683 19224 9711 19264
rect 10612 19236 10640 19264
rect 10689 19261 10701 19295
rect 10735 19292 10747 19295
rect 11164 19292 11192 19332
rect 11330 19320 11336 19332
rect 11388 19320 11394 19372
rect 11514 19360 11520 19372
rect 11475 19332 11520 19360
rect 11514 19320 11520 19332
rect 11572 19320 11578 19372
rect 11624 19332 12572 19360
rect 11624 19292 11652 19332
rect 10735 19264 11192 19292
rect 11348 19264 11652 19292
rect 12544 19292 12572 19332
rect 12618 19320 12624 19372
rect 12676 19360 12682 19372
rect 13078 19360 13084 19372
rect 12676 19332 13084 19360
rect 12676 19320 12682 19332
rect 13078 19320 13084 19332
rect 13136 19360 13142 19372
rect 13541 19363 13599 19369
rect 13541 19360 13553 19363
rect 13136 19332 13553 19360
rect 13136 19320 13142 19332
rect 13541 19329 13553 19332
rect 13587 19329 13599 19363
rect 13722 19360 13728 19372
rect 13683 19332 13728 19360
rect 13541 19323 13599 19329
rect 13722 19320 13728 19332
rect 13780 19320 13786 19372
rect 14458 19360 14464 19372
rect 14419 19332 14464 19360
rect 14458 19320 14464 19332
rect 14516 19320 14522 19372
rect 14737 19363 14795 19369
rect 14737 19329 14749 19363
rect 14783 19329 14795 19363
rect 14737 19323 14795 19329
rect 14921 19363 14979 19369
rect 14921 19329 14933 19363
rect 14967 19360 14979 19363
rect 15378 19360 15384 19372
rect 14967 19332 15384 19360
rect 14967 19329 14979 19332
rect 14921 19323 14979 19329
rect 13354 19292 13360 19304
rect 12544 19264 13360 19292
rect 10735 19261 10747 19264
rect 10689 19255 10747 19261
rect 6512 19196 7144 19224
rect 6512 19184 6518 19196
rect 1302 19156 1308 19168
rect 860 19128 1308 19156
rect 0 19020 800 19034
rect 860 19020 888 19128
rect 1302 19116 1308 19128
rect 1360 19116 1366 19168
rect 2590 19116 2596 19168
rect 2648 19156 2654 19168
rect 2777 19159 2835 19165
rect 2777 19156 2789 19159
rect 2648 19128 2789 19156
rect 2648 19116 2654 19128
rect 2777 19125 2789 19128
rect 2823 19125 2835 19159
rect 2777 19119 2835 19125
rect 2958 19116 2964 19168
rect 3016 19156 3022 19168
rect 3237 19159 3295 19165
rect 3237 19156 3249 19159
rect 3016 19128 3249 19156
rect 3016 19116 3022 19128
rect 3237 19125 3249 19128
rect 3283 19125 3295 19159
rect 3237 19119 3295 19125
rect 4614 19116 4620 19168
rect 4672 19156 4678 19168
rect 7009 19159 7067 19165
rect 7009 19156 7021 19159
rect 4672 19128 7021 19156
rect 4672 19116 4678 19128
rect 7009 19125 7021 19128
rect 7055 19125 7067 19159
rect 7116 19156 7144 19196
rect 8864 19196 9711 19224
rect 8864 19156 8892 19196
rect 10594 19184 10600 19236
rect 10652 19184 10658 19236
rect 10781 19227 10839 19233
rect 10781 19193 10793 19227
rect 10827 19224 10839 19227
rect 11238 19224 11244 19236
rect 10827 19196 11244 19224
rect 10827 19193 10839 19196
rect 10781 19187 10839 19193
rect 11238 19184 11244 19196
rect 11296 19184 11302 19236
rect 11348 19233 11376 19264
rect 13354 19252 13360 19264
rect 13412 19252 13418 19304
rect 13817 19295 13875 19301
rect 13817 19261 13829 19295
rect 13863 19292 13875 19295
rect 14642 19292 14648 19304
rect 13863 19264 14648 19292
rect 13863 19261 13875 19264
rect 13817 19255 13875 19261
rect 14642 19252 14648 19264
rect 14700 19252 14706 19304
rect 14752 19292 14780 19323
rect 15378 19320 15384 19332
rect 15436 19320 15442 19372
rect 15841 19363 15899 19369
rect 15841 19329 15853 19363
rect 15887 19360 15899 19363
rect 16482 19360 16488 19372
rect 15887 19332 16488 19360
rect 15887 19329 15899 19332
rect 15841 19323 15899 19329
rect 16482 19320 16488 19332
rect 16540 19320 16546 19372
rect 16666 19360 16672 19372
rect 16627 19332 16672 19360
rect 16666 19320 16672 19332
rect 16724 19320 16730 19372
rect 15286 19292 15292 19304
rect 14752 19264 15292 19292
rect 15286 19252 15292 19264
rect 15344 19252 15350 19304
rect 15396 19292 15424 19320
rect 15933 19295 15991 19301
rect 15933 19292 15945 19295
rect 15396 19264 15945 19292
rect 15933 19261 15945 19264
rect 15979 19261 15991 19295
rect 16776 19292 16804 19400
rect 17696 19400 18144 19428
rect 16853 19363 16911 19369
rect 16853 19329 16865 19363
rect 16899 19360 16911 19363
rect 17037 19363 17095 19369
rect 17037 19360 17049 19363
rect 16899 19332 17049 19360
rect 16899 19329 16911 19332
rect 16853 19323 16911 19329
rect 17037 19329 17049 19332
rect 17083 19329 17095 19363
rect 17037 19323 17095 19329
rect 17126 19320 17132 19372
rect 17184 19360 17190 19372
rect 17497 19363 17555 19369
rect 17497 19360 17509 19363
rect 17184 19332 17509 19360
rect 17184 19320 17190 19332
rect 17497 19329 17509 19332
rect 17543 19329 17555 19363
rect 17696 19358 17724 19400
rect 18138 19388 18144 19400
rect 18196 19428 18202 19440
rect 18506 19428 18512 19440
rect 18196 19400 18512 19428
rect 18196 19388 18202 19400
rect 18506 19388 18512 19400
rect 18564 19388 18570 19440
rect 23216 19428 23244 19459
rect 23290 19456 23296 19508
rect 23348 19496 23354 19508
rect 25038 19496 25044 19508
rect 23348 19468 25044 19496
rect 23348 19456 23354 19468
rect 18691 19400 23244 19428
rect 17773 19363 17831 19369
rect 17773 19358 17785 19363
rect 17696 19330 17785 19358
rect 17497 19323 17555 19329
rect 17773 19329 17785 19330
rect 17819 19329 17831 19363
rect 17773 19323 17831 19329
rect 17957 19366 18015 19369
rect 18049 19366 18107 19369
rect 17957 19363 18107 19366
rect 17957 19329 17969 19363
rect 18003 19338 18061 19363
rect 18003 19329 18015 19338
rect 17957 19323 18015 19329
rect 18049 19329 18061 19338
rect 18095 19329 18107 19363
rect 18049 19323 18107 19329
rect 18414 19320 18420 19372
rect 18472 19360 18478 19372
rect 18601 19363 18659 19369
rect 18601 19360 18613 19363
rect 18472 19332 18613 19360
rect 18472 19320 18478 19332
rect 18601 19329 18613 19332
rect 18647 19329 18659 19363
rect 18601 19323 18659 19329
rect 18691 19292 18719 19400
rect 23382 19388 23388 19440
rect 23440 19388 23446 19440
rect 18877 19363 18935 19369
rect 18877 19360 18889 19363
rect 16776 19264 17877 19292
rect 15933 19255 15991 19261
rect 11333 19227 11391 19233
rect 11333 19193 11345 19227
rect 11379 19193 11391 19227
rect 15010 19224 15016 19236
rect 11333 19187 11391 19193
rect 13556 19196 15016 19224
rect 9030 19156 9036 19168
rect 7116 19128 8892 19156
rect 8991 19128 9036 19156
rect 7009 19119 7067 19125
rect 9030 19116 9036 19128
rect 9088 19116 9094 19168
rect 9214 19116 9220 19168
rect 9272 19156 9278 19168
rect 10965 19159 11023 19165
rect 10965 19156 10977 19159
rect 9272 19128 10977 19156
rect 9272 19116 9278 19128
rect 10965 19125 10977 19128
rect 11011 19125 11023 19159
rect 10965 19119 11023 19125
rect 11054 19116 11060 19168
rect 11112 19156 11118 19168
rect 11698 19156 11704 19168
rect 11112 19128 11704 19156
rect 11112 19116 11118 19128
rect 11698 19116 11704 19128
rect 11756 19156 11762 19168
rect 13556 19156 13584 19196
rect 15010 19184 15016 19196
rect 15068 19184 15074 19236
rect 17129 19227 17187 19233
rect 17129 19224 17141 19227
rect 15120 19196 17141 19224
rect 11756 19128 13584 19156
rect 11756 19116 11762 19128
rect 13630 19116 13636 19168
rect 13688 19156 13694 19168
rect 15120 19156 15148 19196
rect 17129 19193 17141 19196
rect 17175 19193 17187 19227
rect 17849 19224 17877 19264
rect 18064 19264 18719 19292
rect 18800 19332 18889 19360
rect 18064 19224 18092 19264
rect 18414 19224 18420 19236
rect 17849 19196 18092 19224
rect 18375 19196 18420 19224
rect 17129 19187 17187 19193
rect 18414 19184 18420 19196
rect 18472 19184 18478 19236
rect 18506 19184 18512 19236
rect 18564 19224 18570 19236
rect 18800 19224 18828 19332
rect 18877 19329 18889 19332
rect 18923 19329 18935 19363
rect 18877 19323 18935 19329
rect 19061 19363 19119 19369
rect 19061 19329 19073 19363
rect 19107 19360 19119 19363
rect 19150 19360 19156 19372
rect 19107 19332 19156 19360
rect 19107 19329 19119 19332
rect 19061 19323 19119 19329
rect 19150 19320 19156 19332
rect 19208 19320 19214 19372
rect 19426 19320 19432 19372
rect 19484 19360 19490 19372
rect 19797 19363 19855 19369
rect 19797 19360 19809 19363
rect 19484 19332 19809 19360
rect 19484 19320 19490 19332
rect 19797 19329 19809 19332
rect 19843 19360 19855 19363
rect 20346 19360 20352 19372
rect 19843 19332 20352 19360
rect 19843 19329 19855 19332
rect 19797 19323 19855 19329
rect 20346 19320 20352 19332
rect 20404 19320 20410 19372
rect 20993 19363 21051 19369
rect 20993 19360 21005 19363
rect 20456 19332 21005 19360
rect 19518 19292 19524 19304
rect 19431 19264 19524 19292
rect 19518 19252 19524 19264
rect 19576 19252 19582 19304
rect 20162 19252 20168 19304
rect 20220 19292 20226 19304
rect 20456 19292 20484 19332
rect 20993 19329 21005 19332
rect 21039 19329 21051 19363
rect 21174 19360 21180 19372
rect 21135 19332 21180 19360
rect 20993 19323 21051 19329
rect 21174 19320 21180 19332
rect 21232 19320 21238 19372
rect 22005 19363 22063 19369
rect 22005 19329 22017 19363
rect 22051 19360 22063 19363
rect 22094 19360 22100 19372
rect 22051 19332 22100 19360
rect 22051 19329 22063 19332
rect 22005 19323 22063 19329
rect 22094 19320 22100 19332
rect 22152 19320 22158 19372
rect 22281 19363 22339 19369
rect 22281 19329 22293 19363
rect 22327 19360 22339 19363
rect 22465 19363 22523 19369
rect 22327 19332 22361 19360
rect 22327 19329 22339 19332
rect 22281 19323 22339 19329
rect 22465 19329 22477 19363
rect 22511 19360 22523 19363
rect 23400 19360 23428 19388
rect 22511 19332 23428 19360
rect 22511 19329 22523 19332
rect 22465 19323 22523 19329
rect 20220 19264 20484 19292
rect 20809 19295 20867 19301
rect 20220 19252 20226 19264
rect 20809 19261 20821 19295
rect 20855 19292 20867 19295
rect 21542 19292 21548 19304
rect 20855 19264 21548 19292
rect 20855 19261 20867 19264
rect 20809 19255 20867 19261
rect 21542 19252 21548 19264
rect 21600 19252 21606 19304
rect 22296 19292 22324 19323
rect 22554 19292 22560 19304
rect 22296 19264 22560 19292
rect 22554 19252 22560 19264
rect 22612 19252 22618 19304
rect 23382 19292 23388 19304
rect 23343 19264 23388 19292
rect 23382 19252 23388 19264
rect 23440 19252 23446 19304
rect 23584 19301 23612 19468
rect 25038 19456 25044 19468
rect 25096 19496 25102 19508
rect 25590 19496 25596 19508
rect 25096 19468 25596 19496
rect 25096 19456 25102 19468
rect 25590 19456 25596 19468
rect 25648 19456 25654 19508
rect 25682 19456 25688 19508
rect 25740 19496 25746 19508
rect 27985 19499 28043 19505
rect 25740 19468 26188 19496
rect 25740 19456 25746 19468
rect 25774 19428 25780 19440
rect 24228 19400 25780 19428
rect 24228 19369 24256 19400
rect 25774 19388 25780 19400
rect 25832 19388 25838 19440
rect 24213 19363 24271 19369
rect 24213 19329 24225 19363
rect 24259 19329 24271 19363
rect 24213 19323 24271 19329
rect 24302 19320 24308 19372
rect 24360 19360 24366 19372
rect 24469 19363 24527 19369
rect 24469 19360 24481 19363
rect 24360 19332 24481 19360
rect 24360 19320 24366 19332
rect 24469 19329 24481 19332
rect 24515 19329 24527 19363
rect 24469 19323 24527 19329
rect 24946 19320 24952 19372
rect 25004 19360 25010 19372
rect 26053 19363 26111 19369
rect 26053 19360 26065 19363
rect 25004 19332 26065 19360
rect 25004 19320 25010 19332
rect 26053 19329 26065 19332
rect 26099 19329 26111 19363
rect 26160 19360 26188 19468
rect 27985 19465 27997 19499
rect 28031 19496 28043 19499
rect 28350 19496 28356 19508
rect 28031 19468 28356 19496
rect 28031 19465 28043 19468
rect 27985 19459 28043 19465
rect 28350 19456 28356 19468
rect 28408 19456 28414 19508
rect 28534 19496 28540 19508
rect 28495 19468 28540 19496
rect 28534 19456 28540 19468
rect 28592 19456 28598 19508
rect 29546 19496 29552 19508
rect 28966 19468 29552 19496
rect 28629 19431 28687 19437
rect 28629 19397 28641 19431
rect 28675 19428 28687 19431
rect 28966 19428 28994 19468
rect 29546 19456 29552 19468
rect 29604 19456 29610 19508
rect 30101 19499 30159 19505
rect 30101 19465 30113 19499
rect 30147 19496 30159 19499
rect 30147 19468 31156 19496
rect 30147 19465 30159 19468
rect 30101 19459 30159 19465
rect 28675 19400 28994 19428
rect 28675 19397 28687 19400
rect 28629 19391 28687 19397
rect 29178 19388 29184 19440
rect 29236 19428 29242 19440
rect 29236 19400 29776 19428
rect 29236 19388 29242 19400
rect 26237 19363 26295 19369
rect 26237 19360 26249 19363
rect 26160 19332 26249 19360
rect 26053 19323 26111 19329
rect 26237 19329 26249 19332
rect 26283 19329 26295 19363
rect 26237 19323 26295 19329
rect 27433 19363 27491 19369
rect 27433 19329 27445 19363
rect 27479 19360 27491 19363
rect 28442 19360 28448 19372
rect 27479 19332 28448 19360
rect 27479 19329 27491 19332
rect 27433 19323 27491 19329
rect 28442 19320 28448 19332
rect 28500 19320 28506 19372
rect 28552 19332 28856 19360
rect 23477 19295 23535 19301
rect 23477 19261 23489 19295
rect 23523 19261 23535 19295
rect 23477 19255 23535 19261
rect 23569 19295 23627 19301
rect 23569 19261 23581 19295
rect 23615 19261 23627 19295
rect 23569 19255 23627 19261
rect 23661 19295 23719 19301
rect 23661 19261 23673 19295
rect 23707 19292 23719 19295
rect 23842 19292 23848 19304
rect 23707 19264 23848 19292
rect 23707 19261 23719 19264
rect 23661 19255 23719 19261
rect 18564 19196 18828 19224
rect 18564 19184 18570 19196
rect 18874 19184 18880 19236
rect 18932 19224 18938 19236
rect 19536 19224 19564 19252
rect 18932 19196 19564 19224
rect 23492 19224 23520 19255
rect 23842 19252 23848 19264
rect 23900 19252 23906 19304
rect 25866 19252 25872 19304
rect 25924 19292 25930 19304
rect 27338 19292 27344 19304
rect 25924 19264 27344 19292
rect 25924 19252 25930 19264
rect 27338 19252 27344 19264
rect 27396 19252 27402 19304
rect 27709 19295 27767 19301
rect 27709 19261 27721 19295
rect 27755 19292 27767 19295
rect 28552 19292 28580 19332
rect 27755 19264 28580 19292
rect 27755 19261 27767 19264
rect 27709 19255 27767 19261
rect 28626 19252 28632 19304
rect 28684 19292 28690 19304
rect 28721 19295 28779 19301
rect 28721 19292 28733 19295
rect 28684 19264 28733 19292
rect 28684 19252 28690 19264
rect 28721 19261 28733 19264
rect 28767 19261 28779 19295
rect 28828 19292 28856 19332
rect 29362 19320 29368 19372
rect 29420 19360 29426 19372
rect 29748 19369 29776 19400
rect 30466 19388 30472 19440
rect 30524 19428 30530 19440
rect 30561 19431 30619 19437
rect 30561 19428 30573 19431
rect 30524 19400 30573 19428
rect 30524 19388 30530 19400
rect 30561 19397 30573 19400
rect 30607 19397 30619 19431
rect 30561 19391 30619 19397
rect 29549 19363 29607 19369
rect 29549 19360 29561 19363
rect 29420 19332 29561 19360
rect 29420 19320 29426 19332
rect 29549 19329 29561 19332
rect 29595 19329 29607 19363
rect 29549 19323 29607 19329
rect 29733 19363 29791 19369
rect 29733 19329 29745 19363
rect 29779 19329 29791 19363
rect 29733 19323 29791 19329
rect 29821 19363 29879 19369
rect 29821 19346 29833 19363
rect 29867 19346 29879 19363
rect 29917 19363 29975 19369
rect 29821 19323 29828 19346
rect 29822 19294 29828 19323
rect 29880 19294 29886 19346
rect 29917 19329 29929 19363
rect 29963 19360 29975 19363
rect 30098 19360 30104 19372
rect 29963 19332 30104 19360
rect 29963 19329 29975 19332
rect 29917 19323 29975 19329
rect 30098 19320 30104 19332
rect 30156 19320 30162 19372
rect 30282 19320 30288 19372
rect 30340 19360 30346 19372
rect 30745 19363 30803 19369
rect 30745 19360 30757 19363
rect 30340 19332 30757 19360
rect 30340 19320 30346 19332
rect 30745 19329 30757 19332
rect 30791 19329 30803 19363
rect 30745 19323 30803 19329
rect 30837 19363 30895 19369
rect 30837 19329 30849 19363
rect 30883 19329 30895 19363
rect 31018 19360 31024 19372
rect 30979 19332 31024 19360
rect 30837 19323 30895 19329
rect 28828 19264 29776 19292
rect 28721 19255 28779 19261
rect 28902 19224 28908 19236
rect 23492 19196 23612 19224
rect 18932 19184 18938 19196
rect 13688 19128 15148 19156
rect 13688 19116 13694 19128
rect 15562 19116 15568 19168
rect 15620 19156 15626 19168
rect 16485 19159 16543 19165
rect 16485 19156 16497 19159
rect 15620 19128 16497 19156
rect 15620 19116 15626 19128
rect 16485 19125 16497 19128
rect 16531 19125 16543 19159
rect 17034 19156 17040 19168
rect 16995 19128 17040 19156
rect 16485 19119 16543 19125
rect 17034 19116 17040 19128
rect 17092 19116 17098 19168
rect 17218 19116 17224 19168
rect 17276 19156 17282 19168
rect 17313 19159 17371 19165
rect 17313 19156 17325 19159
rect 17276 19128 17325 19156
rect 17276 19116 17282 19128
rect 17313 19125 17325 19128
rect 17359 19125 17371 19159
rect 17313 19119 17371 19125
rect 17954 19116 17960 19168
rect 18012 19156 18018 19168
rect 18141 19159 18199 19165
rect 18141 19156 18153 19159
rect 18012 19128 18153 19156
rect 18012 19116 18018 19128
rect 18141 19125 18153 19128
rect 18187 19125 18199 19159
rect 18141 19119 18199 19125
rect 18233 19159 18291 19165
rect 18233 19125 18245 19159
rect 18279 19156 18291 19159
rect 21818 19156 21824 19168
rect 18279 19128 21824 19156
rect 18279 19125 18291 19128
rect 18233 19119 18291 19125
rect 21818 19116 21824 19128
rect 21876 19116 21882 19168
rect 22002 19116 22008 19168
rect 22060 19156 22066 19168
rect 23584 19156 23612 19196
rect 25148 19196 28908 19224
rect 25148 19156 25176 19196
rect 28902 19184 28908 19196
rect 28960 19184 28966 19236
rect 29748 19224 29776 19264
rect 30852 19224 30880 19323
rect 31018 19320 31024 19332
rect 31076 19320 31082 19372
rect 31128 19369 31156 19468
rect 31113 19363 31171 19369
rect 31113 19329 31125 19363
rect 31159 19329 31171 19363
rect 31113 19323 31171 19329
rect 31294 19224 31300 19236
rect 29748 19196 31300 19224
rect 31294 19184 31300 19196
rect 31352 19184 31358 19236
rect 26142 19156 26148 19168
rect 22060 19128 25176 19156
rect 26103 19128 26148 19156
rect 22060 19116 22066 19128
rect 26142 19116 26148 19128
rect 26200 19116 26206 19168
rect 27246 19156 27252 19168
rect 27207 19128 27252 19156
rect 27246 19116 27252 19128
rect 27304 19116 27310 19168
rect 27617 19159 27675 19165
rect 27617 19125 27629 19159
rect 27663 19156 27675 19159
rect 27985 19159 28043 19165
rect 27985 19156 27997 19159
rect 27663 19128 27997 19156
rect 27663 19125 27675 19128
rect 27617 19119 27675 19125
rect 27985 19125 27997 19128
rect 28031 19125 28043 19159
rect 27985 19119 28043 19125
rect 28074 19116 28080 19168
rect 28132 19156 28138 19168
rect 28169 19159 28227 19165
rect 28169 19156 28181 19159
rect 28132 19128 28181 19156
rect 28132 19116 28138 19128
rect 28169 19125 28181 19128
rect 28215 19125 28227 19159
rect 28169 19119 28227 19125
rect 0 18992 888 19020
rect 1104 19066 32016 19088
rect 1104 19014 2136 19066
rect 2188 19014 12440 19066
rect 12492 19014 22744 19066
rect 22796 19014 32016 19066
rect 32320 19020 33120 19034
rect 1104 18992 32016 19014
rect 32048 18992 33120 19020
rect 0 18978 800 18992
rect 5442 18912 5448 18964
rect 5500 18952 5506 18964
rect 6638 18952 6644 18964
rect 5500 18924 6316 18952
rect 6599 18924 6644 18952
rect 5500 18912 5506 18924
rect 1397 18887 1455 18893
rect 1397 18853 1409 18887
rect 1443 18884 1455 18887
rect 6288 18884 6316 18924
rect 6638 18912 6644 18924
rect 6696 18912 6702 18964
rect 9677 18955 9735 18961
rect 9677 18952 9689 18955
rect 6748 18924 9689 18952
rect 6748 18884 6776 18924
rect 9677 18921 9689 18924
rect 9723 18921 9735 18955
rect 9677 18915 9735 18921
rect 9769 18955 9827 18961
rect 9769 18921 9781 18955
rect 9815 18952 9827 18955
rect 10502 18952 10508 18964
rect 9815 18924 10508 18952
rect 9815 18921 9827 18924
rect 9769 18915 9827 18921
rect 10502 18912 10508 18924
rect 10560 18912 10566 18964
rect 10594 18912 10600 18964
rect 10652 18952 10658 18964
rect 13817 18955 13875 18961
rect 13817 18952 13829 18955
rect 10652 18924 13829 18952
rect 10652 18912 10658 18924
rect 13817 18921 13829 18924
rect 13863 18921 13875 18955
rect 13817 18915 13875 18921
rect 13906 18912 13912 18964
rect 13964 18952 13970 18964
rect 14277 18955 14335 18961
rect 14277 18952 14289 18955
rect 13964 18924 14289 18952
rect 13964 18912 13970 18924
rect 14277 18921 14289 18924
rect 14323 18921 14335 18955
rect 14277 18915 14335 18921
rect 17681 18955 17739 18961
rect 17681 18921 17693 18955
rect 17727 18952 17739 18955
rect 21174 18952 21180 18964
rect 17727 18924 20760 18952
rect 21087 18924 21180 18952
rect 17727 18921 17739 18924
rect 17681 18915 17739 18921
rect 1443 18856 6224 18884
rect 6288 18856 6776 18884
rect 1443 18853 1455 18856
rect 1397 18847 1455 18853
rect 1946 18776 1952 18828
rect 2004 18816 2010 18828
rect 3970 18816 3976 18828
rect 2004 18788 2268 18816
rect 2004 18776 2010 18788
rect 2240 18757 2268 18788
rect 2516 18788 3976 18816
rect 2516 18757 2544 18788
rect 3970 18776 3976 18788
rect 4028 18776 4034 18828
rect 1581 18751 1639 18757
rect 1581 18717 1593 18751
rect 1627 18717 1639 18751
rect 1581 18711 1639 18717
rect 2225 18751 2283 18757
rect 2225 18717 2237 18751
rect 2271 18717 2283 18751
rect 2225 18711 2283 18717
rect 2501 18751 2559 18757
rect 2501 18717 2513 18751
rect 2547 18717 2559 18751
rect 2501 18711 2559 18717
rect 2685 18751 2743 18757
rect 2685 18717 2697 18751
rect 2731 18717 2743 18751
rect 2685 18711 2743 18717
rect 4525 18751 4583 18757
rect 4525 18717 4537 18751
rect 4571 18748 4583 18751
rect 4706 18748 4712 18760
rect 4571 18720 4712 18748
rect 4571 18717 4583 18720
rect 4525 18711 4583 18717
rect 1596 18680 1624 18711
rect 1596 18652 2544 18680
rect 1946 18572 1952 18624
rect 2004 18612 2010 18624
rect 2041 18615 2099 18621
rect 2041 18612 2053 18615
rect 2004 18584 2053 18612
rect 2004 18572 2010 18584
rect 2041 18581 2053 18584
rect 2087 18581 2099 18615
rect 2516 18612 2544 18652
rect 2590 18640 2596 18692
rect 2648 18680 2654 18692
rect 2700 18680 2728 18711
rect 4706 18708 4712 18720
rect 4764 18708 4770 18760
rect 4801 18751 4859 18757
rect 4801 18717 4813 18751
rect 4847 18748 4859 18751
rect 4890 18748 4896 18760
rect 4847 18720 4896 18748
rect 4847 18717 4859 18720
rect 4801 18711 4859 18717
rect 4890 18708 4896 18720
rect 4948 18708 4954 18760
rect 2648 18652 2728 18680
rect 2648 18640 2654 18652
rect 2866 18640 2872 18692
rect 2924 18680 2930 18692
rect 3881 18683 3939 18689
rect 3881 18680 3893 18683
rect 2924 18652 3893 18680
rect 2924 18640 2930 18652
rect 3881 18649 3893 18652
rect 3927 18649 3939 18683
rect 3881 18643 3939 18649
rect 4065 18683 4123 18689
rect 4065 18649 4077 18683
rect 4111 18680 4123 18683
rect 5166 18680 5172 18692
rect 4111 18652 5172 18680
rect 4111 18649 4123 18652
rect 4065 18643 4123 18649
rect 5166 18640 5172 18652
rect 5224 18640 5230 18692
rect 6196 18680 6224 18856
rect 7190 18844 7196 18896
rect 7248 18884 7254 18896
rect 8113 18887 8171 18893
rect 8113 18884 8125 18887
rect 7248 18856 8125 18884
rect 7248 18844 7254 18856
rect 8113 18853 8125 18856
rect 8159 18853 8171 18887
rect 8113 18847 8171 18853
rect 8570 18844 8576 18896
rect 8628 18884 8634 18896
rect 8941 18887 8999 18893
rect 8941 18884 8953 18887
rect 8628 18856 8953 18884
rect 8628 18844 8634 18856
rect 8941 18853 8953 18856
rect 8987 18853 8999 18887
rect 9950 18884 9956 18896
rect 8941 18847 8999 18853
rect 9232 18856 9956 18884
rect 6273 18819 6331 18825
rect 6273 18785 6285 18819
rect 6319 18816 6331 18819
rect 7006 18816 7012 18828
rect 6319 18788 7012 18816
rect 6319 18785 6331 18788
rect 6273 18779 6331 18785
rect 7006 18776 7012 18788
rect 7064 18776 7070 18828
rect 8662 18776 8668 18828
rect 8720 18816 8726 18828
rect 8720 18788 9168 18816
rect 8720 18776 8726 18788
rect 7024 18748 7052 18776
rect 7377 18751 7435 18757
rect 7377 18748 7389 18751
rect 7024 18720 7389 18748
rect 7377 18717 7389 18720
rect 7423 18717 7435 18751
rect 7377 18711 7435 18717
rect 7469 18751 7527 18757
rect 7469 18717 7481 18751
rect 7515 18748 7527 18751
rect 8018 18748 8024 18760
rect 7515 18720 8024 18748
rect 7515 18717 7527 18720
rect 7469 18711 7527 18717
rect 8018 18708 8024 18720
rect 8076 18748 8082 18760
rect 8297 18751 8355 18757
rect 8297 18748 8309 18751
rect 8076 18720 8309 18748
rect 8076 18708 8082 18720
rect 8297 18717 8309 18720
rect 8343 18717 8355 18751
rect 8297 18711 8355 18717
rect 8389 18751 8447 18757
rect 8389 18717 8401 18751
rect 8435 18748 8447 18751
rect 8754 18748 8760 18760
rect 8435 18720 8760 18748
rect 8435 18717 8447 18720
rect 8389 18711 8447 18717
rect 8754 18708 8760 18720
rect 8812 18708 8818 18760
rect 7558 18680 7564 18692
rect 6196 18652 7564 18680
rect 7558 18640 7564 18652
rect 7616 18640 7622 18692
rect 8113 18683 8171 18689
rect 8113 18649 8125 18683
rect 8159 18680 8171 18683
rect 8941 18683 8999 18689
rect 8941 18680 8953 18683
rect 8159 18652 8953 18680
rect 8159 18649 8171 18652
rect 8113 18643 8171 18649
rect 8941 18649 8953 18652
rect 8987 18680 8999 18683
rect 9030 18680 9036 18692
rect 8987 18652 9036 18680
rect 8987 18649 8999 18652
rect 8941 18643 8999 18649
rect 9030 18640 9036 18652
rect 9088 18640 9094 18692
rect 9140 18680 9168 18788
rect 9232 18757 9260 18856
rect 9950 18844 9956 18856
rect 10008 18884 10014 18896
rect 10008 18856 11836 18884
rect 10008 18844 10014 18856
rect 9398 18776 9404 18828
rect 9456 18816 9462 18828
rect 9456 18788 10180 18816
rect 9456 18776 9462 18788
rect 9217 18751 9275 18757
rect 9217 18717 9229 18751
rect 9263 18748 9275 18751
rect 9306 18748 9312 18760
rect 9263 18720 9312 18748
rect 9263 18717 9275 18720
rect 9217 18711 9275 18717
rect 9306 18708 9312 18720
rect 9364 18708 9370 18760
rect 9674 18708 9680 18760
rect 9732 18748 9738 18760
rect 9953 18751 10011 18757
rect 9953 18748 9965 18751
rect 9732 18720 9965 18748
rect 9732 18708 9738 18720
rect 9953 18717 9965 18720
rect 9999 18717 10011 18751
rect 10152 18748 10180 18788
rect 10594 18776 10600 18828
rect 10652 18816 10658 18828
rect 10652 18788 11192 18816
rect 10652 18776 10658 18788
rect 10226 18761 10284 18767
rect 10226 18748 10238 18761
rect 10152 18727 10238 18748
rect 10272 18727 10284 18761
rect 10152 18721 10284 18727
rect 10965 18751 11023 18757
rect 10152 18720 10272 18721
rect 9953 18711 10011 18717
rect 10965 18717 10977 18751
rect 11011 18748 11023 18751
rect 11054 18748 11060 18760
rect 11011 18720 11060 18748
rect 11011 18717 11023 18720
rect 10965 18711 11023 18717
rect 11054 18708 11060 18720
rect 11112 18708 11118 18760
rect 11164 18748 11192 18788
rect 11422 18776 11428 18828
rect 11480 18816 11486 18828
rect 11698 18816 11704 18828
rect 11480 18788 11704 18816
rect 11480 18776 11486 18788
rect 11698 18776 11704 18788
rect 11756 18776 11762 18828
rect 11330 18748 11336 18760
rect 11164 18720 11336 18748
rect 11330 18708 11336 18720
rect 11388 18748 11394 18760
rect 11808 18757 11836 18856
rect 12250 18844 12256 18896
rect 12308 18884 12314 18896
rect 12618 18884 12624 18896
rect 12308 18856 12624 18884
rect 12308 18844 12314 18856
rect 12618 18844 12624 18856
rect 12676 18884 12682 18896
rect 12713 18887 12771 18893
rect 12713 18884 12725 18887
rect 12676 18856 12725 18884
rect 12676 18844 12682 18856
rect 12713 18853 12725 18856
rect 12759 18853 12771 18887
rect 12713 18847 12771 18853
rect 12802 18844 12808 18896
rect 12860 18884 12866 18896
rect 17313 18887 17371 18893
rect 12860 18856 16804 18884
rect 12860 18844 12866 18856
rect 11977 18819 12035 18825
rect 11977 18785 11989 18819
rect 12023 18816 12035 18819
rect 13725 18819 13783 18825
rect 13725 18816 13737 18819
rect 12023 18788 13737 18816
rect 12023 18785 12035 18788
rect 11977 18779 12035 18785
rect 13725 18785 13737 18788
rect 13771 18785 13783 18819
rect 13725 18779 13783 18785
rect 13817 18819 13875 18825
rect 13817 18785 13829 18819
rect 13863 18816 13875 18819
rect 16666 18816 16672 18828
rect 13863 18788 16672 18816
rect 13863 18785 13875 18788
rect 13817 18779 13875 18785
rect 16666 18776 16672 18788
rect 16724 18776 16730 18828
rect 16776 18816 16804 18856
rect 17313 18853 17325 18887
rect 17359 18884 17371 18887
rect 18966 18884 18972 18896
rect 17359 18856 18972 18884
rect 17359 18853 17371 18856
rect 17313 18847 17371 18853
rect 18966 18844 18972 18856
rect 19024 18844 19030 18896
rect 20732 18884 20760 18924
rect 21174 18912 21180 18924
rect 21232 18952 21238 18964
rect 22186 18952 22192 18964
rect 21232 18924 22192 18952
rect 21232 18912 21238 18924
rect 22186 18912 22192 18924
rect 22244 18952 22250 18964
rect 22281 18955 22339 18961
rect 22281 18952 22293 18955
rect 22244 18924 22293 18952
rect 22244 18912 22250 18924
rect 22281 18921 22293 18924
rect 22327 18952 22339 18955
rect 23014 18952 23020 18964
rect 22327 18924 23020 18952
rect 22327 18921 22339 18924
rect 22281 18915 22339 18921
rect 23014 18912 23020 18924
rect 23072 18912 23078 18964
rect 23842 18952 23848 18964
rect 23803 18924 23848 18952
rect 23842 18912 23848 18924
rect 23900 18912 23906 18964
rect 24486 18912 24492 18964
rect 24544 18952 24550 18964
rect 25682 18952 25688 18964
rect 24544 18924 25688 18952
rect 24544 18912 24550 18924
rect 25682 18912 25688 18924
rect 25740 18912 25746 18964
rect 32048 18952 32076 18992
rect 32320 18978 33120 18992
rect 25792 18924 32076 18952
rect 25792 18884 25820 18924
rect 20732 18856 25820 18884
rect 27338 18844 27344 18896
rect 27396 18884 27402 18896
rect 28902 18884 28908 18896
rect 27396 18856 28304 18884
rect 28863 18856 28908 18884
rect 27396 18844 27402 18856
rect 17681 18819 17739 18825
rect 17681 18816 17693 18819
rect 16776 18788 17693 18816
rect 17681 18785 17693 18788
rect 17727 18785 17739 18819
rect 18230 18816 18236 18828
rect 18191 18788 18236 18816
rect 17681 18779 17739 18785
rect 18230 18776 18236 18788
rect 18288 18776 18294 18828
rect 18506 18776 18512 18828
rect 18564 18816 18570 18828
rect 18782 18816 18788 18828
rect 18564 18788 18788 18816
rect 18564 18776 18570 18788
rect 11609 18751 11667 18757
rect 11609 18748 11621 18751
rect 11388 18720 11621 18748
rect 11388 18708 11394 18720
rect 11609 18717 11621 18720
rect 11655 18717 11667 18751
rect 11609 18711 11667 18717
rect 11793 18751 11851 18757
rect 11793 18717 11805 18751
rect 11839 18717 11851 18751
rect 13170 18748 13176 18760
rect 13131 18720 13176 18748
rect 11793 18711 11851 18717
rect 13170 18708 13176 18720
rect 13228 18708 13234 18760
rect 13446 18708 13452 18760
rect 13504 18748 13510 18760
rect 14093 18751 14151 18757
rect 14093 18748 14105 18751
rect 13504 18720 14105 18748
rect 13504 18708 13510 18720
rect 14093 18717 14105 18720
rect 14139 18748 14151 18751
rect 14182 18748 14188 18760
rect 14139 18720 14188 18748
rect 14139 18717 14151 18720
rect 14093 18711 14151 18717
rect 14182 18708 14188 18720
rect 14240 18708 14246 18760
rect 15102 18708 15108 18760
rect 15160 18748 15166 18760
rect 15289 18751 15347 18757
rect 15289 18748 15301 18751
rect 15160 18720 15301 18748
rect 15160 18708 15166 18720
rect 15289 18717 15301 18720
rect 15335 18717 15347 18751
rect 15289 18711 15347 18717
rect 15378 18708 15384 18760
rect 15436 18748 15442 18760
rect 15565 18751 15623 18757
rect 15565 18748 15577 18751
rect 15436 18720 15577 18748
rect 15436 18708 15442 18720
rect 15565 18717 15577 18720
rect 15611 18717 15623 18751
rect 15565 18711 15623 18717
rect 16758 18708 16764 18760
rect 16816 18748 16822 18760
rect 16945 18751 17003 18757
rect 16945 18748 16957 18751
rect 16816 18720 16957 18748
rect 16816 18708 16822 18720
rect 16945 18717 16957 18720
rect 16991 18717 17003 18751
rect 16945 18711 17003 18717
rect 17129 18751 17187 18757
rect 17129 18717 17141 18751
rect 17175 18748 17187 18751
rect 17218 18748 17224 18760
rect 17175 18720 17224 18748
rect 17175 18717 17187 18720
rect 17129 18711 17187 18717
rect 17218 18708 17224 18720
rect 17276 18708 17282 18760
rect 17405 18751 17463 18757
rect 17405 18717 17417 18751
rect 17451 18748 17463 18751
rect 17451 18720 17724 18748
rect 17451 18717 17463 18720
rect 17405 18711 17463 18717
rect 10134 18680 10140 18692
rect 9140 18652 10140 18680
rect 10134 18640 10140 18652
rect 10192 18640 10198 18692
rect 11149 18683 11207 18689
rect 10704 18652 11100 18680
rect 5442 18612 5448 18624
rect 2516 18584 5448 18612
rect 2041 18575 2099 18581
rect 5442 18572 5448 18584
rect 5500 18572 5506 18624
rect 5994 18572 6000 18624
rect 6052 18612 6058 18624
rect 6454 18612 6460 18624
rect 6052 18584 6460 18612
rect 6052 18572 6058 18584
rect 6454 18572 6460 18584
rect 6512 18612 6518 18624
rect 6641 18615 6699 18621
rect 6641 18612 6653 18615
rect 6512 18584 6653 18612
rect 6512 18572 6518 18584
rect 6641 18581 6653 18584
rect 6687 18581 6699 18615
rect 6641 18575 6699 18581
rect 6730 18572 6736 18624
rect 6788 18612 6794 18624
rect 6825 18615 6883 18621
rect 6825 18612 6837 18615
rect 6788 18584 6837 18612
rect 6788 18572 6794 18584
rect 6825 18581 6837 18584
rect 6871 18581 6883 18615
rect 6825 18575 6883 18581
rect 7742 18572 7748 18624
rect 7800 18612 7806 18624
rect 9125 18615 9183 18621
rect 9125 18612 9137 18615
rect 7800 18584 9137 18612
rect 7800 18572 7806 18584
rect 9125 18581 9137 18584
rect 9171 18581 9183 18615
rect 9125 18575 9183 18581
rect 9677 18615 9735 18621
rect 9677 18581 9689 18615
rect 9723 18612 9735 18615
rect 10704 18612 10732 18652
rect 9723 18584 10732 18612
rect 9723 18581 9735 18584
rect 9677 18575 9735 18581
rect 10778 18572 10784 18624
rect 10836 18612 10842 18624
rect 10962 18612 10968 18624
rect 10836 18584 10968 18612
rect 10836 18572 10842 18584
rect 10962 18572 10968 18584
rect 11020 18572 11026 18624
rect 11072 18612 11100 18652
rect 11149 18649 11161 18683
rect 11195 18680 11207 18683
rect 12529 18683 12587 18689
rect 11195 18652 12434 18680
rect 11195 18649 11207 18652
rect 11149 18643 11207 18649
rect 12158 18612 12164 18624
rect 11072 18584 12164 18612
rect 12158 18572 12164 18584
rect 12216 18572 12222 18624
rect 12406 18612 12434 18652
rect 12529 18649 12541 18683
rect 12575 18680 12587 18683
rect 12894 18680 12900 18692
rect 12575 18652 12900 18680
rect 12575 18649 12587 18652
rect 12529 18643 12587 18649
rect 12894 18640 12900 18652
rect 12952 18640 12958 18692
rect 15930 18680 15936 18692
rect 13188 18652 15936 18680
rect 13188 18612 13216 18652
rect 15930 18640 15936 18652
rect 15988 18640 15994 18692
rect 17034 18640 17040 18692
rect 17092 18680 17098 18692
rect 17420 18680 17448 18711
rect 17696 18692 17724 18720
rect 18322 18708 18328 18760
rect 18380 18748 18386 18760
rect 18709 18757 18737 18788
rect 18782 18776 18788 18788
rect 18840 18776 18846 18828
rect 19242 18776 19248 18828
rect 19300 18816 19306 18828
rect 19797 18819 19855 18825
rect 19797 18816 19809 18819
rect 19300 18788 19809 18816
rect 19300 18776 19306 18788
rect 19797 18785 19809 18788
rect 19843 18785 19855 18819
rect 19797 18779 19855 18785
rect 20990 18776 20996 18828
rect 21048 18816 21054 18828
rect 23750 18816 23756 18828
rect 21048 18788 23756 18816
rect 21048 18776 21054 18788
rect 23750 18776 23756 18788
rect 23808 18816 23814 18828
rect 24489 18819 24547 18825
rect 24489 18816 24501 18819
rect 23808 18788 24501 18816
rect 23808 18776 23814 18788
rect 24489 18785 24501 18788
rect 24535 18785 24547 18819
rect 24489 18779 24547 18785
rect 27249 18819 27307 18825
rect 27249 18785 27261 18819
rect 27295 18816 27307 18819
rect 28169 18819 28227 18825
rect 28169 18816 28181 18819
rect 27295 18788 28181 18816
rect 27295 18785 27307 18788
rect 27249 18779 27307 18785
rect 28169 18785 28181 18788
rect 28215 18785 28227 18819
rect 28276 18816 28304 18856
rect 28902 18844 28908 18856
rect 28960 18844 28966 18896
rect 29549 18887 29607 18893
rect 29549 18853 29561 18887
rect 29595 18853 29607 18887
rect 30190 18884 30196 18896
rect 30151 18856 30196 18884
rect 29549 18847 29607 18853
rect 29564 18816 29592 18847
rect 30190 18844 30196 18856
rect 30248 18844 30254 18896
rect 28276 18788 29592 18816
rect 28169 18779 28227 18785
rect 18417 18751 18475 18757
rect 18417 18748 18429 18751
rect 18380 18720 18429 18748
rect 18380 18708 18386 18720
rect 18417 18717 18429 18720
rect 18463 18717 18475 18751
rect 18417 18711 18475 18717
rect 18693 18751 18751 18757
rect 18693 18717 18705 18751
rect 18739 18717 18751 18751
rect 20898 18748 20904 18760
rect 18693 18711 18751 18717
rect 18800 18720 20904 18748
rect 17092 18652 17448 18680
rect 17092 18640 17098 18652
rect 17678 18640 17684 18692
rect 17736 18640 17742 18692
rect 18800 18680 18828 18720
rect 20898 18708 20904 18720
rect 20956 18708 20962 18760
rect 21726 18708 21732 18760
rect 21784 18748 21790 18760
rect 21913 18751 21971 18757
rect 21913 18748 21925 18751
rect 21784 18720 21925 18748
rect 21784 18708 21790 18720
rect 21913 18717 21925 18720
rect 21959 18717 21971 18751
rect 21913 18711 21971 18717
rect 23201 18751 23259 18757
rect 23201 18717 23213 18751
rect 23247 18748 23259 18751
rect 23290 18748 23296 18760
rect 23247 18720 23296 18748
rect 23247 18717 23259 18720
rect 23201 18711 23259 18717
rect 23290 18708 23296 18720
rect 23348 18708 23354 18760
rect 23477 18751 23535 18757
rect 23477 18717 23489 18751
rect 23523 18748 23535 18751
rect 24026 18748 24032 18760
rect 23523 18720 24032 18748
rect 23523 18717 23535 18720
rect 23477 18711 23535 18717
rect 24026 18708 24032 18720
rect 24084 18708 24090 18760
rect 24578 18708 24584 18760
rect 24636 18748 24642 18760
rect 24765 18751 24823 18757
rect 24765 18748 24777 18751
rect 24636 18720 24777 18748
rect 24636 18708 24642 18720
rect 24765 18717 24777 18720
rect 24811 18717 24823 18751
rect 25774 18748 25780 18760
rect 25735 18720 25780 18748
rect 24765 18711 24823 18717
rect 25774 18708 25780 18720
rect 25832 18708 25838 18760
rect 26050 18757 26056 18760
rect 26044 18748 26056 18757
rect 26011 18720 26056 18748
rect 26044 18711 26056 18720
rect 26050 18708 26056 18711
rect 26108 18708 26114 18760
rect 28074 18708 28080 18760
rect 28132 18748 28138 18760
rect 28132 18720 28177 18748
rect 28132 18708 28138 18720
rect 28534 18708 28540 18760
rect 28592 18748 28598 18760
rect 28813 18751 28871 18757
rect 28813 18748 28825 18751
rect 28592 18720 28825 18748
rect 28592 18708 28598 18720
rect 28813 18717 28825 18720
rect 28859 18717 28871 18751
rect 28813 18711 28871 18717
rect 29733 18751 29791 18757
rect 29733 18717 29745 18751
rect 29779 18717 29791 18751
rect 29733 18711 29791 18717
rect 30377 18751 30435 18757
rect 30377 18717 30389 18751
rect 30423 18717 30435 18751
rect 30377 18711 30435 18717
rect 17788 18652 18828 18680
rect 13354 18612 13360 18624
rect 12406 18584 13216 18612
rect 13315 18584 13360 18612
rect 13354 18572 13360 18584
rect 13412 18572 13418 18624
rect 13725 18615 13783 18621
rect 13725 18581 13737 18615
rect 13771 18612 13783 18615
rect 13814 18612 13820 18624
rect 13771 18584 13820 18612
rect 13771 18581 13783 18584
rect 13725 18575 13783 18581
rect 13814 18572 13820 18584
rect 13872 18572 13878 18624
rect 17218 18572 17224 18624
rect 17276 18612 17282 18624
rect 17788 18612 17816 18652
rect 19518 18640 19524 18692
rect 19576 18680 19582 18692
rect 20042 18683 20100 18689
rect 20042 18680 20054 18683
rect 19576 18652 20054 18680
rect 19576 18640 19582 18652
rect 20042 18649 20054 18652
rect 20088 18649 20100 18683
rect 20042 18643 20100 18649
rect 21634 18640 21640 18692
rect 21692 18680 21698 18692
rect 23686 18683 23744 18689
rect 23686 18680 23698 18683
rect 21692 18652 23698 18680
rect 21692 18640 21698 18652
rect 23686 18649 23698 18652
rect 23732 18649 23744 18683
rect 23686 18643 23744 18649
rect 24670 18640 24676 18692
rect 24728 18680 24734 18692
rect 27249 18683 27307 18689
rect 27249 18680 27261 18683
rect 24728 18652 27261 18680
rect 24728 18640 24734 18652
rect 27249 18649 27261 18652
rect 27295 18649 27307 18683
rect 27982 18680 27988 18692
rect 27943 18652 27988 18680
rect 27249 18643 27307 18649
rect 27982 18640 27988 18652
rect 28040 18640 28046 18692
rect 28626 18640 28632 18692
rect 28684 18680 28690 18692
rect 29748 18680 29776 18711
rect 30190 18680 30196 18692
rect 28684 18652 30196 18680
rect 28684 18640 28690 18652
rect 30190 18640 30196 18652
rect 30248 18640 30254 18692
rect 30392 18680 30420 18711
rect 30466 18708 30472 18760
rect 30524 18748 30530 18760
rect 30650 18748 30656 18760
rect 30524 18720 30656 18748
rect 30524 18708 30530 18720
rect 30650 18708 30656 18720
rect 30708 18708 30714 18760
rect 30837 18751 30895 18757
rect 30837 18717 30849 18751
rect 30883 18748 30895 18751
rect 31110 18748 31116 18760
rect 30883 18720 31116 18748
rect 30883 18717 30895 18720
rect 30837 18711 30895 18717
rect 31110 18708 31116 18720
rect 31168 18708 31174 18760
rect 30742 18680 30748 18692
rect 30392 18652 30748 18680
rect 30742 18640 30748 18652
rect 30800 18640 30806 18692
rect 17276 18584 17816 18612
rect 17276 18572 17282 18584
rect 17954 18572 17960 18624
rect 18012 18612 18018 18624
rect 18601 18615 18659 18621
rect 18601 18612 18613 18615
rect 18012 18584 18613 18612
rect 18012 18572 18018 18584
rect 18601 18581 18613 18584
rect 18647 18612 18659 18615
rect 19334 18612 19340 18624
rect 18647 18584 19340 18612
rect 18647 18581 18659 18584
rect 18601 18575 18659 18581
rect 19334 18572 19340 18584
rect 19392 18612 19398 18624
rect 20714 18612 20720 18624
rect 19392 18584 20720 18612
rect 19392 18572 19398 18584
rect 20714 18572 20720 18584
rect 20772 18572 20778 18624
rect 22281 18615 22339 18621
rect 22281 18581 22293 18615
rect 22327 18612 22339 18615
rect 22370 18612 22376 18624
rect 22327 18584 22376 18612
rect 22327 18581 22339 18584
rect 22281 18575 22339 18581
rect 22370 18572 22376 18584
rect 22428 18572 22434 18624
rect 22465 18615 22523 18621
rect 22465 18581 22477 18615
rect 22511 18612 22523 18615
rect 23014 18612 23020 18624
rect 22511 18584 23020 18612
rect 22511 18581 22523 18584
rect 22465 18575 22523 18581
rect 23014 18572 23020 18584
rect 23072 18572 23078 18624
rect 23569 18615 23627 18621
rect 23569 18581 23581 18615
rect 23615 18612 23627 18615
rect 23842 18612 23848 18624
rect 23615 18584 23848 18612
rect 23615 18581 23627 18584
rect 23569 18575 23627 18581
rect 23842 18572 23848 18584
rect 23900 18612 23906 18624
rect 24118 18612 24124 18624
rect 23900 18584 24124 18612
rect 23900 18572 23906 18584
rect 24118 18572 24124 18584
rect 24176 18572 24182 18624
rect 24486 18572 24492 18624
rect 24544 18612 24550 18624
rect 27062 18612 27068 18624
rect 24544 18584 27068 18612
rect 24544 18572 24550 18584
rect 27062 18572 27068 18584
rect 27120 18572 27126 18624
rect 27157 18615 27215 18621
rect 27157 18581 27169 18615
rect 27203 18612 27215 18615
rect 27522 18612 27528 18624
rect 27203 18584 27528 18612
rect 27203 18581 27215 18584
rect 27157 18575 27215 18581
rect 27522 18572 27528 18584
rect 27580 18572 27586 18624
rect 27617 18615 27675 18621
rect 27617 18581 27629 18615
rect 27663 18612 27675 18615
rect 28810 18612 28816 18624
rect 27663 18584 28816 18612
rect 27663 18581 27675 18584
rect 27617 18575 27675 18581
rect 28810 18572 28816 18584
rect 28868 18572 28874 18624
rect 28994 18572 29000 18624
rect 29052 18612 29058 18624
rect 30834 18612 30840 18624
rect 29052 18584 30840 18612
rect 29052 18572 29058 18584
rect 30834 18572 30840 18584
rect 30892 18572 30898 18624
rect 1104 18522 32016 18544
rect 1104 18470 7288 18522
rect 7340 18470 17592 18522
rect 17644 18470 27896 18522
rect 27948 18470 32016 18522
rect 1104 18448 32016 18470
rect 1670 18368 1676 18420
rect 1728 18408 1734 18420
rect 1765 18411 1823 18417
rect 1765 18408 1777 18411
rect 1728 18380 1777 18408
rect 1728 18368 1734 18380
rect 1765 18377 1777 18380
rect 1811 18377 1823 18411
rect 1765 18371 1823 18377
rect 3697 18411 3755 18417
rect 3697 18377 3709 18411
rect 3743 18408 3755 18411
rect 6086 18408 6092 18420
rect 3743 18380 6092 18408
rect 3743 18377 3755 18380
rect 3697 18371 3755 18377
rect 6086 18368 6092 18380
rect 6144 18368 6150 18420
rect 6362 18408 6368 18420
rect 6323 18380 6368 18408
rect 6362 18368 6368 18380
rect 6420 18368 6426 18420
rect 6917 18411 6975 18417
rect 6917 18377 6929 18411
rect 6963 18408 6975 18411
rect 7190 18408 7196 18420
rect 6963 18380 7196 18408
rect 6963 18377 6975 18380
rect 6917 18371 6975 18377
rect 7190 18368 7196 18380
rect 7248 18368 7254 18420
rect 7466 18408 7472 18420
rect 7427 18380 7472 18408
rect 7466 18368 7472 18380
rect 7524 18368 7530 18420
rect 7558 18368 7564 18420
rect 7616 18408 7622 18420
rect 14458 18408 14464 18420
rect 7616 18380 14464 18408
rect 7616 18368 7622 18380
rect 14458 18368 14464 18380
rect 14516 18368 14522 18420
rect 15010 18368 15016 18420
rect 15068 18408 15074 18420
rect 15068 18380 17356 18408
rect 15068 18368 15074 18380
rect 2222 18340 2228 18352
rect 2148 18312 2228 18340
rect 1946 18272 1952 18284
rect 1907 18244 1952 18272
rect 1946 18232 1952 18244
rect 2004 18232 2010 18284
rect 2148 18145 2176 18312
rect 2222 18300 2228 18312
rect 2280 18300 2286 18352
rect 3786 18340 3792 18352
rect 2792 18312 3792 18340
rect 2225 18207 2283 18213
rect 2225 18173 2237 18207
rect 2271 18204 2283 18207
rect 2682 18204 2688 18216
rect 2271 18176 2688 18204
rect 2271 18173 2283 18176
rect 2225 18167 2283 18173
rect 2682 18164 2688 18176
rect 2740 18204 2746 18216
rect 2792 18204 2820 18312
rect 3786 18300 3792 18312
rect 3844 18300 3850 18352
rect 4154 18349 4160 18352
rect 4148 18340 4160 18349
rect 4115 18312 4160 18340
rect 4148 18303 4160 18312
rect 4154 18300 4160 18303
rect 4212 18300 4218 18352
rect 5442 18300 5448 18352
rect 5500 18340 5506 18352
rect 5500 18312 7052 18340
rect 5500 18300 5506 18312
rect 2958 18272 2964 18284
rect 2919 18244 2964 18272
rect 2958 18232 2964 18244
rect 3016 18232 3022 18284
rect 3142 18232 3148 18284
rect 3200 18272 3206 18284
rect 6609 18275 6667 18281
rect 3200 18244 4936 18272
rect 3200 18232 3206 18244
rect 4908 18216 4936 18244
rect 6609 18241 6621 18275
rect 6655 18272 6667 18275
rect 6917 18275 6975 18281
rect 6917 18272 6929 18275
rect 6655 18244 6929 18272
rect 6655 18241 6667 18244
rect 6609 18235 6667 18241
rect 6917 18241 6929 18244
rect 6963 18241 6975 18275
rect 6917 18235 6975 18241
rect 2740 18176 2820 18204
rect 3237 18207 3295 18213
rect 2740 18164 2746 18176
rect 3237 18173 3249 18207
rect 3283 18204 3295 18207
rect 3697 18207 3755 18213
rect 3697 18204 3709 18207
rect 3283 18176 3709 18204
rect 3283 18173 3295 18176
rect 3237 18167 3295 18173
rect 3697 18173 3709 18176
rect 3743 18173 3755 18207
rect 3878 18204 3884 18216
rect 3839 18176 3884 18204
rect 3697 18167 3755 18173
rect 3878 18164 3884 18176
rect 3936 18164 3942 18216
rect 4890 18164 4896 18216
rect 4948 18204 4954 18216
rect 6733 18207 6791 18213
rect 6733 18204 6745 18207
rect 4948 18176 6745 18204
rect 4948 18164 4954 18176
rect 6733 18173 6745 18176
rect 6779 18173 6791 18207
rect 6733 18167 6791 18173
rect 6825 18207 6883 18213
rect 6825 18173 6837 18207
rect 6871 18173 6883 18207
rect 7024 18204 7052 18312
rect 7098 18300 7104 18352
rect 7156 18340 7162 18352
rect 8665 18343 8723 18349
rect 8665 18340 8677 18343
rect 7156 18312 8677 18340
rect 7156 18300 7162 18312
rect 8665 18309 8677 18312
rect 8711 18309 8723 18343
rect 8665 18303 8723 18309
rect 8754 18300 8760 18352
rect 8812 18340 8818 18352
rect 8849 18343 8907 18349
rect 8849 18340 8861 18343
rect 8812 18312 8861 18340
rect 8812 18300 8818 18312
rect 8849 18309 8861 18312
rect 8895 18309 8907 18343
rect 8849 18303 8907 18309
rect 7650 18272 7656 18284
rect 7611 18244 7656 18272
rect 7650 18232 7656 18244
rect 7708 18232 7714 18284
rect 7742 18232 7748 18284
rect 7800 18272 7806 18284
rect 7926 18272 7932 18284
rect 7800 18244 7845 18272
rect 7887 18244 7932 18272
rect 7800 18232 7806 18244
rect 7926 18232 7932 18244
rect 7984 18232 7990 18284
rect 8018 18232 8024 18284
rect 8076 18272 8082 18284
rect 8864 18272 8892 18303
rect 9030 18300 9036 18352
rect 9088 18340 9094 18352
rect 13630 18340 13636 18352
rect 9088 18312 13636 18340
rect 9088 18300 9094 18312
rect 13630 18300 13636 18312
rect 13688 18300 13694 18352
rect 13814 18340 13820 18352
rect 13740 18312 13820 18340
rect 9306 18272 9312 18284
rect 8076 18244 8121 18272
rect 8864 18244 9312 18272
rect 8076 18232 8082 18244
rect 9306 18232 9312 18244
rect 9364 18232 9370 18284
rect 9493 18275 9551 18281
rect 9493 18241 9505 18275
rect 9539 18272 9551 18275
rect 10229 18275 10287 18281
rect 10229 18272 10241 18275
rect 9539 18244 10241 18272
rect 9539 18241 9551 18244
rect 9493 18235 9551 18241
rect 10229 18241 10241 18244
rect 10275 18241 10287 18275
rect 10410 18272 10416 18284
rect 10371 18244 10416 18272
rect 10229 18235 10287 18241
rect 10410 18232 10416 18244
rect 10468 18232 10474 18284
rect 10689 18275 10747 18281
rect 10689 18241 10701 18275
rect 10735 18241 10747 18275
rect 10870 18272 10876 18284
rect 10831 18244 10876 18272
rect 10689 18235 10747 18241
rect 9214 18204 9220 18216
rect 7024 18176 9220 18204
rect 6825 18167 6883 18173
rect 2133 18139 2191 18145
rect 2133 18105 2145 18139
rect 2179 18136 2191 18139
rect 3142 18136 3148 18148
rect 2179 18108 3148 18136
rect 2179 18105 2191 18108
rect 2133 18099 2191 18105
rect 3142 18096 3148 18108
rect 3200 18096 3206 18148
rect 6638 18096 6644 18148
rect 6696 18136 6702 18148
rect 6840 18136 6868 18167
rect 9214 18164 9220 18176
rect 9272 18164 9278 18216
rect 9582 18164 9588 18216
rect 9640 18204 9646 18216
rect 9769 18207 9827 18213
rect 9769 18204 9781 18207
rect 9640 18176 9781 18204
rect 9640 18164 9646 18176
rect 9769 18173 9781 18176
rect 9815 18173 9827 18207
rect 9769 18167 9827 18173
rect 10042 18164 10048 18216
rect 10100 18204 10106 18216
rect 10594 18204 10600 18216
rect 10100 18176 10600 18204
rect 10100 18164 10106 18176
rect 10594 18164 10600 18176
rect 10652 18164 10658 18216
rect 10704 18204 10732 18235
rect 10870 18232 10876 18244
rect 10928 18232 10934 18284
rect 11698 18272 11704 18284
rect 11624 18244 11704 18272
rect 11624 18204 11652 18244
rect 11698 18232 11704 18244
rect 11756 18232 11762 18284
rect 11793 18275 11851 18281
rect 11793 18241 11805 18275
rect 11839 18272 11851 18275
rect 11882 18272 11888 18284
rect 11839 18244 11888 18272
rect 11839 18241 11851 18244
rect 11793 18235 11851 18241
rect 11882 18232 11888 18244
rect 11940 18232 11946 18284
rect 12069 18275 12127 18281
rect 12069 18241 12081 18275
rect 12115 18272 12127 18275
rect 12250 18272 12256 18284
rect 12115 18244 12256 18272
rect 12115 18241 12127 18244
rect 12069 18235 12127 18241
rect 12250 18232 12256 18244
rect 12308 18232 12314 18284
rect 12526 18232 12532 18284
rect 12584 18272 12590 18284
rect 12989 18275 13047 18281
rect 12989 18272 13001 18275
rect 12584 18244 13001 18272
rect 12584 18232 12590 18244
rect 12989 18241 13001 18244
rect 13035 18272 13047 18275
rect 13170 18272 13176 18284
rect 13035 18244 13176 18272
rect 13035 18241 13047 18244
rect 12989 18235 13047 18241
rect 13170 18232 13176 18244
rect 13228 18232 13234 18284
rect 13740 18281 13768 18312
rect 13814 18300 13820 18312
rect 13872 18340 13878 18352
rect 17328 18340 17356 18380
rect 17402 18368 17408 18420
rect 17460 18408 17466 18420
rect 17770 18408 17776 18420
rect 17460 18380 17776 18408
rect 17460 18368 17466 18380
rect 17770 18368 17776 18380
rect 17828 18368 17834 18420
rect 17954 18368 17960 18420
rect 18012 18408 18018 18420
rect 18049 18411 18107 18417
rect 18049 18408 18061 18411
rect 18012 18380 18061 18408
rect 18012 18368 18018 18380
rect 18049 18377 18061 18380
rect 18095 18408 18107 18411
rect 18230 18408 18236 18420
rect 18095 18380 18236 18408
rect 18095 18377 18107 18380
rect 18049 18371 18107 18377
rect 18230 18368 18236 18380
rect 18288 18368 18294 18420
rect 18322 18368 18328 18420
rect 18380 18408 18386 18420
rect 19242 18408 19248 18420
rect 18380 18380 19248 18408
rect 18380 18368 18386 18380
rect 19242 18368 19248 18380
rect 19300 18368 19306 18420
rect 19518 18408 19524 18420
rect 19479 18380 19524 18408
rect 19518 18368 19524 18380
rect 19576 18368 19582 18420
rect 22002 18408 22008 18420
rect 21963 18380 22008 18408
rect 22002 18368 22008 18380
rect 22060 18368 22066 18420
rect 22094 18368 22100 18420
rect 22152 18408 22158 18420
rect 22370 18408 22376 18420
rect 22152 18380 22376 18408
rect 22152 18368 22158 18380
rect 22370 18368 22376 18380
rect 22428 18368 22434 18420
rect 23382 18368 23388 18420
rect 23440 18408 23446 18420
rect 24210 18408 24216 18420
rect 23440 18380 24216 18408
rect 23440 18368 23446 18380
rect 24210 18368 24216 18380
rect 24268 18368 24274 18420
rect 24305 18411 24363 18417
rect 24305 18377 24317 18411
rect 24351 18408 24363 18411
rect 26142 18408 26148 18420
rect 24351 18380 26148 18408
rect 24351 18377 24363 18380
rect 24305 18371 24363 18377
rect 26142 18368 26148 18380
rect 26200 18408 26206 18420
rect 26789 18411 26847 18417
rect 26789 18408 26801 18411
rect 26200 18380 26801 18408
rect 26200 18368 26206 18380
rect 26789 18377 26801 18380
rect 26835 18377 26847 18411
rect 26970 18408 26976 18420
rect 26931 18380 26976 18408
rect 26789 18371 26847 18377
rect 26970 18368 26976 18380
rect 27028 18368 27034 18420
rect 27706 18368 27712 18420
rect 27764 18408 27770 18420
rect 28277 18411 28335 18417
rect 28277 18408 28289 18411
rect 27764 18380 28289 18408
rect 27764 18368 27770 18380
rect 28277 18377 28289 18380
rect 28323 18377 28335 18411
rect 28277 18371 28335 18377
rect 28442 18368 28448 18420
rect 28500 18408 28506 18420
rect 28905 18411 28963 18417
rect 28905 18408 28917 18411
rect 28500 18380 28917 18408
rect 28500 18368 28506 18380
rect 28905 18377 28917 18380
rect 28951 18377 28963 18411
rect 29178 18408 29184 18420
rect 28905 18371 28963 18377
rect 29012 18380 29184 18408
rect 18509 18343 18567 18349
rect 13872 18312 16712 18340
rect 17328 18312 18000 18340
rect 13872 18300 13878 18312
rect 13725 18275 13783 18281
rect 13725 18241 13737 18275
rect 13771 18241 13783 18275
rect 13725 18235 13783 18241
rect 13992 18275 14050 18281
rect 13992 18241 14004 18275
rect 14038 18272 14050 18275
rect 15565 18275 15623 18281
rect 15565 18272 15577 18275
rect 14038 18244 15577 18272
rect 14038 18241 14050 18244
rect 13992 18235 14050 18241
rect 15565 18241 15577 18244
rect 15611 18241 15623 18275
rect 15565 18235 15623 18241
rect 15749 18275 15807 18281
rect 15749 18241 15761 18275
rect 15795 18241 15807 18275
rect 16022 18272 16028 18284
rect 15983 18244 16028 18272
rect 15749 18235 15807 18241
rect 10704 18176 11652 18204
rect 11716 18176 12020 18204
rect 6696 18108 6868 18136
rect 9140 18108 10180 18136
rect 6696 18096 6702 18108
rect 2222 18028 2228 18080
rect 2280 18068 2286 18080
rect 2777 18071 2835 18077
rect 2777 18068 2789 18071
rect 2280 18040 2789 18068
rect 2280 18028 2286 18040
rect 2777 18037 2789 18040
rect 2823 18037 2835 18071
rect 2777 18031 2835 18037
rect 5074 18028 5080 18080
rect 5132 18068 5138 18080
rect 5261 18071 5319 18077
rect 5261 18068 5273 18071
rect 5132 18040 5273 18068
rect 5132 18028 5138 18040
rect 5261 18037 5273 18040
rect 5307 18037 5319 18071
rect 5261 18031 5319 18037
rect 5902 18028 5908 18080
rect 5960 18068 5966 18080
rect 9140 18068 9168 18108
rect 5960 18040 9168 18068
rect 5960 18028 5966 18040
rect 9214 18028 9220 18080
rect 9272 18068 9278 18080
rect 9309 18071 9367 18077
rect 9309 18068 9321 18071
rect 9272 18040 9321 18068
rect 9272 18028 9278 18040
rect 9309 18037 9321 18040
rect 9355 18037 9367 18071
rect 9309 18031 9367 18037
rect 9677 18071 9735 18077
rect 9677 18037 9689 18071
rect 9723 18068 9735 18071
rect 10042 18068 10048 18080
rect 9723 18040 10048 18068
rect 9723 18037 9735 18040
rect 9677 18031 9735 18037
rect 10042 18028 10048 18040
rect 10100 18028 10106 18080
rect 10152 18068 10180 18108
rect 10318 18096 10324 18148
rect 10376 18136 10382 18148
rect 10962 18136 10968 18148
rect 10376 18108 10968 18136
rect 10376 18096 10382 18108
rect 10962 18096 10968 18108
rect 11020 18096 11026 18148
rect 11054 18096 11060 18148
rect 11112 18136 11118 18148
rect 11609 18139 11667 18145
rect 11609 18136 11621 18139
rect 11112 18108 11621 18136
rect 11112 18096 11118 18108
rect 11609 18105 11621 18108
rect 11655 18105 11667 18139
rect 11609 18099 11667 18105
rect 11716 18068 11744 18176
rect 11992 18136 12020 18176
rect 12158 18164 12164 18216
rect 12216 18204 12222 18216
rect 12216 18176 13216 18204
rect 12216 18164 12222 18176
rect 12802 18136 12808 18148
rect 11992 18108 12808 18136
rect 12802 18096 12808 18108
rect 12860 18096 12866 18148
rect 13188 18145 13216 18176
rect 14826 18164 14832 18216
rect 14884 18204 14890 18216
rect 15764 18204 15792 18235
rect 16022 18232 16028 18244
rect 16080 18232 16086 18284
rect 16684 18281 16712 18312
rect 17972 18284 18000 18312
rect 18509 18309 18521 18343
rect 18555 18340 18567 18343
rect 18598 18340 18604 18352
rect 18555 18312 18604 18340
rect 18555 18309 18567 18312
rect 18509 18303 18567 18309
rect 18598 18300 18604 18312
rect 18656 18300 18662 18352
rect 20254 18340 20260 18352
rect 18708 18312 20260 18340
rect 16669 18275 16727 18281
rect 16669 18241 16681 18275
rect 16715 18241 16727 18275
rect 16669 18235 16727 18241
rect 16758 18232 16764 18284
rect 16816 18272 16822 18284
rect 16925 18275 16983 18281
rect 16925 18272 16937 18275
rect 16816 18244 16937 18272
rect 16816 18232 16822 18244
rect 16925 18241 16937 18244
rect 16971 18241 16983 18275
rect 16925 18235 16983 18241
rect 17402 18232 17408 18284
rect 17460 18278 17466 18284
rect 17460 18272 17522 18278
rect 17460 18250 17715 18272
rect 17460 18232 17466 18250
rect 17494 18244 17715 18250
rect 15930 18204 15936 18216
rect 14884 18176 15792 18204
rect 15891 18176 15936 18204
rect 14884 18164 14890 18176
rect 15930 18164 15936 18176
rect 15988 18164 15994 18216
rect 17687 18204 17715 18244
rect 17954 18232 17960 18284
rect 18012 18232 18018 18284
rect 18138 18232 18144 18284
rect 18196 18272 18202 18284
rect 18414 18272 18420 18284
rect 18196 18244 18420 18272
rect 18196 18232 18202 18244
rect 18414 18232 18420 18244
rect 18472 18232 18478 18284
rect 18708 18281 18736 18312
rect 20254 18300 20260 18312
rect 20312 18300 20318 18352
rect 21818 18340 21824 18352
rect 21779 18312 21824 18340
rect 21818 18300 21824 18312
rect 21876 18300 21882 18352
rect 24118 18340 24124 18352
rect 21928 18312 24124 18340
rect 18694 18275 18752 18281
rect 18694 18241 18706 18275
rect 18740 18241 18752 18275
rect 18694 18235 18752 18241
rect 18785 18275 18843 18281
rect 18785 18241 18797 18275
rect 18831 18241 18843 18275
rect 18785 18235 18843 18241
rect 19061 18275 19119 18281
rect 19061 18241 19073 18275
rect 19107 18272 19119 18275
rect 19334 18272 19340 18284
rect 19107 18244 19340 18272
rect 19107 18241 19119 18244
rect 19061 18235 19119 18241
rect 18800 18204 18828 18235
rect 19334 18232 19340 18244
rect 19392 18232 19398 18284
rect 19705 18275 19763 18281
rect 19705 18241 19717 18275
rect 19751 18272 19763 18275
rect 20441 18275 20499 18281
rect 20441 18272 20453 18275
rect 19751 18244 20453 18272
rect 19751 18241 19763 18244
rect 19705 18235 19763 18241
rect 20441 18241 20453 18244
rect 20487 18241 20499 18275
rect 20441 18235 20499 18241
rect 20625 18275 20683 18281
rect 20625 18241 20637 18275
rect 20671 18241 20683 18275
rect 20625 18235 20683 18241
rect 20901 18275 20959 18281
rect 20901 18241 20913 18275
rect 20947 18241 20959 18275
rect 20901 18235 20959 18241
rect 17687 18176 18828 18204
rect 13173 18139 13231 18145
rect 13173 18105 13185 18139
rect 13219 18105 13231 18139
rect 13173 18099 13231 18105
rect 15028 18108 16712 18136
rect 10152 18040 11744 18068
rect 11977 18071 12035 18077
rect 11977 18037 11989 18071
rect 12023 18068 12035 18071
rect 12158 18068 12164 18080
rect 12023 18040 12164 18068
rect 12023 18037 12035 18040
rect 11977 18031 12035 18037
rect 12158 18028 12164 18040
rect 12216 18028 12222 18080
rect 12342 18028 12348 18080
rect 12400 18068 12406 18080
rect 12894 18068 12900 18080
rect 12400 18040 12900 18068
rect 12400 18028 12406 18040
rect 12894 18028 12900 18040
rect 12952 18028 12958 18080
rect 13188 18068 13216 18099
rect 15028 18068 15056 18108
rect 13188 18040 15056 18068
rect 15105 18071 15163 18077
rect 15105 18037 15117 18071
rect 15151 18068 15163 18071
rect 15470 18068 15476 18080
rect 15151 18040 15476 18068
rect 15151 18037 15163 18040
rect 15105 18031 15163 18037
rect 15470 18028 15476 18040
rect 15528 18028 15534 18080
rect 15838 18028 15844 18080
rect 15896 18068 15902 18080
rect 16022 18068 16028 18080
rect 15896 18040 16028 18068
rect 15896 18028 15902 18040
rect 16022 18028 16028 18040
rect 16080 18028 16086 18080
rect 16684 18068 16712 18108
rect 17862 18096 17868 18148
rect 17920 18136 17926 18148
rect 18322 18136 18328 18148
rect 17920 18108 18328 18136
rect 17920 18096 17926 18108
rect 18322 18096 18328 18108
rect 18380 18096 18386 18148
rect 18800 18136 18828 18176
rect 19981 18207 20039 18213
rect 19981 18173 19993 18207
rect 20027 18204 20039 18207
rect 20254 18204 20260 18216
rect 20027 18176 20260 18204
rect 20027 18173 20039 18176
rect 19981 18167 20039 18173
rect 20254 18164 20260 18176
rect 20312 18164 20318 18216
rect 20346 18164 20352 18216
rect 20404 18204 20410 18216
rect 20640 18204 20668 18235
rect 20404 18176 20668 18204
rect 20404 18164 20410 18176
rect 20916 18136 20944 18235
rect 20990 18232 20996 18284
rect 21048 18272 21054 18284
rect 21085 18275 21143 18281
rect 21085 18272 21097 18275
rect 21048 18244 21097 18272
rect 21048 18232 21054 18244
rect 21085 18241 21097 18244
rect 21131 18272 21143 18275
rect 21174 18272 21180 18284
rect 21131 18244 21180 18272
rect 21131 18241 21143 18244
rect 21085 18235 21143 18241
rect 21174 18232 21180 18244
rect 21232 18232 21238 18284
rect 21358 18232 21364 18284
rect 21416 18272 21422 18284
rect 21928 18272 21956 18312
rect 24118 18300 24124 18312
rect 24176 18300 24182 18352
rect 24397 18343 24455 18349
rect 24397 18309 24409 18343
rect 24443 18340 24455 18343
rect 24486 18340 24492 18352
rect 24443 18312 24492 18340
rect 24443 18309 24455 18312
rect 24397 18303 24455 18309
rect 24486 18300 24492 18312
rect 24544 18300 24550 18352
rect 24613 18343 24671 18349
rect 24613 18309 24625 18343
rect 24659 18340 24671 18343
rect 25130 18340 25136 18352
rect 24659 18312 25136 18340
rect 24659 18309 24671 18312
rect 24613 18303 24671 18309
rect 25130 18300 25136 18312
rect 25188 18300 25194 18352
rect 27062 18300 27068 18352
rect 27120 18340 27126 18352
rect 28077 18343 28135 18349
rect 27120 18312 28028 18340
rect 27120 18300 27126 18312
rect 22094 18272 22100 18284
rect 21416 18244 21956 18272
rect 22055 18244 22100 18272
rect 21416 18232 21422 18244
rect 22094 18232 22100 18244
rect 22152 18232 22158 18284
rect 22824 18275 22882 18281
rect 22824 18241 22836 18275
rect 22870 18272 22882 18275
rect 23106 18272 23112 18284
rect 22870 18244 23112 18272
rect 22870 18241 22882 18244
rect 22824 18235 22882 18241
rect 23106 18232 23112 18244
rect 23164 18232 23170 18284
rect 23750 18232 23756 18284
rect 23808 18272 23814 18284
rect 25225 18275 25283 18281
rect 25225 18272 25237 18275
rect 23808 18244 25237 18272
rect 23808 18232 23814 18244
rect 25225 18241 25237 18244
rect 25271 18241 25283 18275
rect 25225 18235 25283 18241
rect 25501 18275 25559 18281
rect 25501 18241 25513 18275
rect 25547 18272 25559 18275
rect 25866 18272 25872 18284
rect 25547 18244 25872 18272
rect 25547 18241 25559 18244
rect 25501 18235 25559 18241
rect 25866 18232 25872 18244
rect 25924 18272 25930 18284
rect 27157 18275 27215 18281
rect 27157 18272 27169 18275
rect 25924 18244 27169 18272
rect 25924 18232 25930 18244
rect 27157 18241 27169 18244
rect 27203 18241 27215 18275
rect 27157 18235 27215 18241
rect 27338 18232 27344 18284
rect 27396 18272 27402 18284
rect 27433 18275 27491 18281
rect 27433 18272 27445 18275
rect 27396 18244 27445 18272
rect 27396 18232 27402 18244
rect 27433 18241 27445 18244
rect 27479 18241 27491 18275
rect 27433 18235 27491 18241
rect 27522 18232 27528 18284
rect 27580 18272 27586 18284
rect 27617 18275 27675 18281
rect 27617 18272 27629 18275
rect 27580 18244 27629 18272
rect 27580 18232 27586 18244
rect 27617 18241 27629 18244
rect 27663 18241 27675 18275
rect 28000 18272 28028 18312
rect 28077 18309 28089 18343
rect 28123 18340 28135 18343
rect 29012 18340 29040 18380
rect 29178 18368 29184 18380
rect 29236 18368 29242 18420
rect 29641 18411 29699 18417
rect 29641 18408 29653 18411
rect 29380 18380 29653 18408
rect 28123 18312 29040 18340
rect 28123 18309 28135 18312
rect 28077 18303 28135 18309
rect 28994 18272 29000 18284
rect 28000 18244 29000 18272
rect 27617 18235 27675 18241
rect 28994 18232 29000 18244
rect 29052 18232 29058 18284
rect 29086 18232 29092 18284
rect 29144 18272 29150 18284
rect 29380 18281 29408 18380
rect 29641 18377 29653 18380
rect 29687 18377 29699 18411
rect 30006 18408 30012 18420
rect 29967 18380 30012 18408
rect 29641 18371 29699 18377
rect 30006 18368 30012 18380
rect 30064 18368 30070 18420
rect 29365 18275 29423 18281
rect 29144 18244 29189 18272
rect 29144 18232 29150 18244
rect 29365 18241 29377 18275
rect 29411 18241 29423 18275
rect 29503 18275 29561 18281
rect 29503 18272 29515 18275
rect 29365 18235 29423 18241
rect 29481 18241 29515 18272
rect 29549 18241 29561 18275
rect 29481 18235 29561 18241
rect 21910 18164 21916 18216
rect 21968 18204 21974 18216
rect 22557 18207 22615 18213
rect 22557 18204 22569 18207
rect 21968 18176 22569 18204
rect 21968 18164 21974 18176
rect 22557 18173 22569 18176
rect 22603 18173 22615 18207
rect 28166 18204 28172 18216
rect 22557 18167 22615 18173
rect 25148 18176 28172 18204
rect 23937 18139 23995 18145
rect 18800 18108 20300 18136
rect 20916 18108 22094 18136
rect 18874 18068 18880 18080
rect 16684 18040 18880 18068
rect 18874 18028 18880 18040
rect 18932 18028 18938 18080
rect 18969 18071 19027 18077
rect 18969 18037 18981 18071
rect 19015 18068 19027 18071
rect 19242 18068 19248 18080
rect 19015 18040 19248 18068
rect 19015 18037 19027 18040
rect 18969 18031 19027 18037
rect 19242 18028 19248 18040
rect 19300 18028 19306 18080
rect 19334 18028 19340 18080
rect 19392 18068 19398 18080
rect 19794 18068 19800 18080
rect 19392 18040 19800 18068
rect 19392 18028 19398 18040
rect 19794 18028 19800 18040
rect 19852 18028 19858 18080
rect 19889 18071 19947 18077
rect 19889 18037 19901 18071
rect 19935 18068 19947 18071
rect 20162 18068 20168 18080
rect 19935 18040 20168 18068
rect 19935 18037 19947 18040
rect 19889 18031 19947 18037
rect 20162 18028 20168 18040
rect 20220 18028 20226 18080
rect 20272 18068 20300 18108
rect 21634 18068 21640 18080
rect 20272 18040 21640 18068
rect 21634 18028 21640 18040
rect 21692 18028 21698 18080
rect 21818 18068 21824 18080
rect 21779 18040 21824 18068
rect 21818 18028 21824 18040
rect 21876 18028 21882 18080
rect 22066 18068 22094 18108
rect 23937 18105 23949 18139
rect 23983 18136 23995 18139
rect 24026 18136 24032 18148
rect 23983 18108 24032 18136
rect 23983 18105 23995 18108
rect 23937 18099 23995 18105
rect 24026 18096 24032 18108
rect 24084 18136 24090 18148
rect 24486 18136 24492 18148
rect 24084 18108 24492 18136
rect 24084 18096 24090 18108
rect 24486 18096 24492 18108
rect 24544 18136 24550 18148
rect 24765 18139 24823 18145
rect 24544 18108 24716 18136
rect 24544 18096 24550 18108
rect 22554 18068 22560 18080
rect 22066 18040 22560 18068
rect 22554 18028 22560 18040
rect 22612 18068 22618 18080
rect 23198 18068 23204 18080
rect 22612 18040 23204 18068
rect 22612 18028 22618 18040
rect 23198 18028 23204 18040
rect 23256 18028 23262 18080
rect 24305 18071 24363 18077
rect 24305 18037 24317 18071
rect 24351 18068 24363 18071
rect 24581 18071 24639 18077
rect 24581 18068 24593 18071
rect 24351 18040 24593 18068
rect 24351 18037 24363 18040
rect 24305 18031 24363 18037
rect 24581 18037 24593 18040
rect 24627 18037 24639 18071
rect 24688 18068 24716 18108
rect 24765 18105 24777 18139
rect 24811 18136 24823 18139
rect 25148 18136 25176 18176
rect 28166 18164 28172 18176
rect 28224 18164 28230 18216
rect 28534 18204 28540 18216
rect 28276 18176 28540 18204
rect 28276 18136 28304 18176
rect 28534 18164 28540 18176
rect 28592 18164 28598 18216
rect 29178 18164 29184 18216
rect 29236 18204 29242 18216
rect 29481 18204 29509 18235
rect 30181 18232 30187 18284
rect 30239 18281 30245 18284
rect 30239 18272 30251 18281
rect 30834 18272 30840 18284
rect 30239 18244 30284 18272
rect 30795 18244 30840 18272
rect 30239 18235 30251 18244
rect 30239 18232 30245 18235
rect 30834 18232 30840 18244
rect 30892 18232 30898 18284
rect 31113 18275 31171 18281
rect 31113 18241 31125 18275
rect 31159 18241 31171 18275
rect 31294 18272 31300 18284
rect 31255 18244 31300 18272
rect 31113 18235 31171 18241
rect 29236 18176 29509 18204
rect 29641 18207 29699 18213
rect 29236 18164 29242 18176
rect 29641 18173 29653 18207
rect 29687 18204 29699 18207
rect 30466 18204 30472 18216
rect 29687 18176 30472 18204
rect 29687 18173 29699 18176
rect 29641 18167 29699 18173
rect 30466 18164 30472 18176
rect 30524 18204 30530 18216
rect 31128 18204 31156 18235
rect 31294 18232 31300 18244
rect 31352 18232 31358 18284
rect 30524 18176 31156 18204
rect 30524 18164 30530 18176
rect 24811 18108 25176 18136
rect 25220 18108 28304 18136
rect 28445 18139 28503 18145
rect 24811 18105 24823 18108
rect 24765 18099 24823 18105
rect 25220 18068 25248 18108
rect 28445 18105 28457 18139
rect 28491 18136 28503 18139
rect 31018 18136 31024 18148
rect 28491 18108 31024 18136
rect 28491 18105 28503 18108
rect 28445 18099 28503 18105
rect 31018 18096 31024 18108
rect 31076 18096 31082 18148
rect 24688 18040 25248 18068
rect 24581 18031 24639 18037
rect 25498 18028 25504 18080
rect 25556 18068 25562 18080
rect 26142 18068 26148 18080
rect 25556 18040 26148 18068
rect 25556 18028 25562 18040
rect 26142 18028 26148 18040
rect 26200 18028 26206 18080
rect 26789 18071 26847 18077
rect 26789 18037 26801 18071
rect 26835 18068 26847 18071
rect 27798 18068 27804 18080
rect 26835 18040 27804 18068
rect 26835 18037 26847 18040
rect 26789 18031 26847 18037
rect 27798 18028 27804 18040
rect 27856 18068 27862 18080
rect 28261 18071 28319 18077
rect 28261 18068 28273 18071
rect 27856 18040 28273 18068
rect 27856 18028 27862 18040
rect 28261 18037 28273 18040
rect 28307 18037 28319 18071
rect 28261 18031 28319 18037
rect 30653 18071 30711 18077
rect 30653 18037 30665 18071
rect 30699 18068 30711 18071
rect 30742 18068 30748 18080
rect 30699 18040 30748 18068
rect 30699 18037 30711 18040
rect 30653 18031 30711 18037
rect 30742 18028 30748 18040
rect 30800 18028 30806 18080
rect 1104 17978 32016 18000
rect 1104 17926 2136 17978
rect 2188 17926 12440 17978
rect 12492 17926 22744 17978
rect 22796 17926 32016 17978
rect 1104 17904 32016 17926
rect 2777 17867 2835 17873
rect 2777 17833 2789 17867
rect 2823 17864 2835 17867
rect 3050 17864 3056 17876
rect 2823 17836 3056 17864
rect 2823 17833 2835 17836
rect 2777 17827 2835 17833
rect 3050 17824 3056 17836
rect 3108 17824 3114 17876
rect 3142 17824 3148 17876
rect 3200 17864 3206 17876
rect 3200 17836 3245 17864
rect 3200 17824 3206 17836
rect 4062 17824 4068 17876
rect 4120 17864 4126 17876
rect 4982 17864 4988 17876
rect 4120 17836 4988 17864
rect 4120 17824 4126 17836
rect 4982 17824 4988 17836
rect 5040 17864 5046 17876
rect 5169 17867 5227 17873
rect 5169 17864 5181 17867
rect 5040 17836 5181 17864
rect 5040 17824 5046 17836
rect 5169 17833 5181 17836
rect 5215 17833 5227 17867
rect 5169 17827 5227 17833
rect 5534 17824 5540 17876
rect 5592 17864 5598 17876
rect 6822 17864 6828 17876
rect 5592 17836 6828 17864
rect 5592 17824 5598 17836
rect 6822 17824 6828 17836
rect 6880 17864 6886 17876
rect 7374 17864 7380 17876
rect 6880 17836 7380 17864
rect 6880 17824 6886 17836
rect 7374 17824 7380 17836
rect 7432 17824 7438 17876
rect 7561 17867 7619 17873
rect 7561 17833 7573 17867
rect 7607 17864 7619 17867
rect 7650 17864 7656 17876
rect 7607 17836 7656 17864
rect 7607 17833 7619 17836
rect 7561 17827 7619 17833
rect 7650 17824 7656 17836
rect 7708 17824 7714 17876
rect 10134 17824 10140 17876
rect 10192 17864 10198 17876
rect 14182 17864 14188 17876
rect 10192 17836 14188 17864
rect 10192 17824 10198 17836
rect 14182 17824 14188 17836
rect 14240 17824 14246 17876
rect 14277 17867 14335 17873
rect 14277 17833 14289 17867
rect 14323 17864 14335 17867
rect 18141 17867 18199 17873
rect 14323 17836 18092 17864
rect 14323 17833 14335 17836
rect 14277 17827 14335 17833
rect 934 17756 940 17808
rect 992 17796 998 17808
rect 2041 17799 2099 17805
rect 2041 17796 2053 17799
rect 992 17768 2053 17796
rect 992 17756 998 17768
rect 2041 17765 2053 17768
rect 2087 17796 2099 17799
rect 4614 17796 4620 17808
rect 2087 17768 4620 17796
rect 2087 17765 2099 17768
rect 2041 17759 2099 17765
rect 4614 17756 4620 17768
rect 4672 17756 4678 17808
rect 8202 17756 8208 17808
rect 8260 17796 8266 17808
rect 8260 17768 9996 17796
rect 8260 17756 8266 17768
rect 1673 17731 1731 17737
rect 1673 17697 1685 17731
rect 1719 17728 1731 17731
rect 2682 17728 2688 17740
rect 1719 17700 2688 17728
rect 1719 17697 1731 17700
rect 1673 17691 1731 17697
rect 2682 17688 2688 17700
rect 2740 17688 2746 17740
rect 3050 17688 3056 17740
rect 3108 17728 3114 17740
rect 3237 17731 3295 17737
rect 3237 17728 3249 17731
rect 3108 17700 3249 17728
rect 3108 17688 3114 17700
rect 3237 17697 3249 17700
rect 3283 17697 3295 17731
rect 3237 17691 3295 17697
rect 5626 17688 5632 17740
rect 5684 17728 5690 17740
rect 5721 17731 5779 17737
rect 5721 17728 5733 17731
rect 5684 17700 5733 17728
rect 5684 17688 5690 17700
rect 5721 17697 5733 17700
rect 5767 17697 5779 17731
rect 5721 17691 5779 17697
rect 8113 17731 8171 17737
rect 8113 17697 8125 17731
rect 8159 17728 8171 17731
rect 8386 17728 8392 17740
rect 8159 17700 8392 17728
rect 8159 17697 8171 17700
rect 8113 17691 8171 17697
rect 8386 17688 8392 17700
rect 8444 17688 8450 17740
rect 9968 17728 9996 17768
rect 10042 17756 10048 17808
rect 10100 17796 10106 17808
rect 10778 17796 10784 17808
rect 10100 17768 10784 17796
rect 10100 17756 10106 17768
rect 10778 17756 10784 17768
rect 10836 17756 10842 17808
rect 11425 17799 11483 17805
rect 11425 17765 11437 17799
rect 11471 17796 11483 17799
rect 11514 17796 11520 17808
rect 11471 17768 11520 17796
rect 11471 17765 11483 17768
rect 11425 17759 11483 17765
rect 11514 17756 11520 17768
rect 11572 17756 11578 17808
rect 12253 17799 12311 17805
rect 12253 17796 12265 17799
rect 11624 17768 12265 17796
rect 11238 17728 11244 17740
rect 9968 17700 11244 17728
rect 11238 17688 11244 17700
rect 11296 17688 11302 17740
rect 11333 17731 11391 17737
rect 11333 17697 11345 17731
rect 11379 17728 11391 17731
rect 11624 17728 11652 17768
rect 12253 17765 12265 17768
rect 12299 17765 12311 17799
rect 12253 17759 12311 17765
rect 12345 17799 12403 17805
rect 12345 17765 12357 17799
rect 12391 17796 12403 17799
rect 12618 17796 12624 17808
rect 12391 17768 12624 17796
rect 12391 17765 12403 17768
rect 12345 17759 12403 17765
rect 12618 17756 12624 17768
rect 12676 17756 12682 17808
rect 12986 17756 12992 17808
rect 13044 17796 13050 17808
rect 17218 17796 17224 17808
rect 13044 17768 17224 17796
rect 13044 17756 13050 17768
rect 17218 17756 17224 17768
rect 17276 17756 17282 17808
rect 17494 17756 17500 17808
rect 17552 17796 17558 17808
rect 17954 17796 17960 17808
rect 17552 17768 17960 17796
rect 17552 17756 17558 17768
rect 17954 17756 17960 17768
rect 18012 17756 18018 17808
rect 11379 17700 11652 17728
rect 11992 17700 13124 17728
rect 11379 17697 11391 17700
rect 11333 17691 11391 17697
rect 11992 17672 12020 17700
rect 2866 17660 2872 17672
rect 768 17632 2872 17660
rect 768 17388 796 17632
rect 2866 17620 2872 17632
rect 2924 17620 2930 17672
rect 2961 17663 3019 17669
rect 2961 17629 2973 17663
rect 3007 17629 3019 17663
rect 2961 17623 3019 17629
rect 1486 17552 1492 17604
rect 1544 17592 1550 17604
rect 2976 17592 3004 17623
rect 3602 17620 3608 17672
rect 3660 17660 3666 17672
rect 3973 17663 4031 17669
rect 3973 17660 3985 17663
rect 3660 17632 3985 17660
rect 3660 17620 3666 17632
rect 3973 17629 3985 17632
rect 4019 17629 4031 17663
rect 3973 17623 4031 17629
rect 4062 17620 4068 17672
rect 4120 17660 4126 17672
rect 4249 17663 4307 17669
rect 4249 17660 4261 17663
rect 4120 17632 4261 17660
rect 4120 17620 4126 17632
rect 4249 17629 4261 17632
rect 4295 17629 4307 17663
rect 4430 17660 4436 17672
rect 4391 17632 4436 17660
rect 4249 17623 4307 17629
rect 4430 17620 4436 17632
rect 4488 17620 4494 17672
rect 6546 17620 6552 17672
rect 6604 17660 6610 17672
rect 8021 17663 8079 17669
rect 8021 17660 8033 17663
rect 6604 17632 8033 17660
rect 6604 17620 6610 17632
rect 8021 17629 8033 17632
rect 8067 17660 8079 17663
rect 8202 17660 8208 17672
rect 8067 17632 8208 17660
rect 8067 17629 8079 17632
rect 8021 17623 8079 17629
rect 8202 17620 8208 17632
rect 8260 17620 8266 17672
rect 10410 17620 10416 17672
rect 10468 17660 10474 17672
rect 11514 17660 11520 17672
rect 10468 17632 11520 17660
rect 10468 17620 10474 17632
rect 11514 17620 11520 17632
rect 11572 17660 11578 17672
rect 11701 17663 11759 17669
rect 11701 17660 11713 17663
rect 11572 17632 11713 17660
rect 11572 17620 11578 17632
rect 11701 17629 11713 17632
rect 11747 17629 11759 17663
rect 11974 17660 11980 17672
rect 11935 17632 11980 17660
rect 11701 17623 11759 17629
rect 3789 17595 3847 17601
rect 3789 17592 3801 17595
rect 1544 17564 2820 17592
rect 2976 17564 3801 17592
rect 1544 17552 1550 17564
rect 2038 17484 2044 17536
rect 2096 17524 2102 17536
rect 2133 17527 2191 17533
rect 2133 17524 2145 17527
rect 2096 17496 2145 17524
rect 2096 17484 2102 17496
rect 2133 17493 2145 17496
rect 2179 17493 2191 17527
rect 2792 17524 2820 17564
rect 3789 17561 3801 17564
rect 3835 17561 3847 17595
rect 5074 17592 5080 17604
rect 5035 17564 5080 17592
rect 3789 17555 3847 17561
rect 5074 17552 5080 17564
rect 5132 17552 5138 17604
rect 5988 17595 6046 17601
rect 5988 17561 6000 17595
rect 6034 17592 6046 17595
rect 6914 17592 6920 17604
rect 6034 17564 6920 17592
rect 6034 17561 6046 17564
rect 5988 17555 6046 17561
rect 6914 17552 6920 17564
rect 6972 17552 6978 17604
rect 9309 17595 9367 17601
rect 9309 17592 9321 17595
rect 7024 17564 9321 17592
rect 2866 17524 2872 17536
rect 2792 17496 2872 17524
rect 2133 17487 2191 17493
rect 2866 17484 2872 17496
rect 2924 17484 2930 17536
rect 3510 17484 3516 17536
rect 3568 17524 3574 17536
rect 7024 17524 7052 17564
rect 9309 17561 9321 17564
rect 9355 17592 9367 17595
rect 11333 17595 11391 17601
rect 11333 17592 11345 17595
rect 9355 17564 11345 17592
rect 9355 17561 9367 17564
rect 9309 17555 9367 17561
rect 11333 17561 11345 17564
rect 11379 17561 11391 17595
rect 11716 17592 11744 17623
rect 11974 17620 11980 17632
rect 12032 17620 12038 17672
rect 13096 17669 13124 17700
rect 13354 17688 13360 17740
rect 13412 17728 13418 17740
rect 16485 17731 16543 17737
rect 16485 17728 16497 17731
rect 13412 17700 16497 17728
rect 13412 17688 13418 17700
rect 16485 17697 16497 17700
rect 16531 17697 16543 17731
rect 16485 17691 16543 17697
rect 17773 17731 17831 17737
rect 17773 17697 17785 17731
rect 17819 17728 17831 17731
rect 17862 17728 17868 17740
rect 17819 17700 17868 17728
rect 17819 17697 17831 17700
rect 17773 17691 17831 17697
rect 17862 17688 17868 17700
rect 17920 17688 17926 17740
rect 18064 17728 18092 17836
rect 18141 17833 18153 17867
rect 18187 17864 18199 17867
rect 18966 17864 18972 17876
rect 18187 17836 18972 17864
rect 18187 17833 18199 17836
rect 18141 17827 18199 17833
rect 18966 17824 18972 17836
rect 19024 17824 19030 17876
rect 20990 17864 20996 17876
rect 20732 17836 20996 17864
rect 19794 17796 19800 17808
rect 18340 17768 19800 17796
rect 18340 17728 18368 17768
rect 19794 17756 19800 17768
rect 19852 17756 19858 17808
rect 18064 17700 18368 17728
rect 20257 17731 20315 17737
rect 20257 17697 20269 17731
rect 20303 17728 20315 17731
rect 20732 17728 20760 17836
rect 20990 17824 20996 17836
rect 21048 17824 21054 17876
rect 21726 17824 21732 17876
rect 21784 17864 21790 17876
rect 22097 17867 22155 17873
rect 22097 17864 22109 17867
rect 21784 17836 22109 17864
rect 21784 17824 21790 17836
rect 22097 17833 22109 17836
rect 22143 17864 22155 17867
rect 23201 17867 23259 17873
rect 23201 17864 23213 17867
rect 22143 17836 23213 17864
rect 22143 17833 22155 17836
rect 22097 17827 22155 17833
rect 23201 17833 23213 17836
rect 23247 17833 23259 17867
rect 23750 17864 23756 17876
rect 23711 17836 23756 17864
rect 23201 17827 23259 17833
rect 23750 17824 23756 17836
rect 23808 17824 23814 17876
rect 24118 17824 24124 17876
rect 24176 17864 24182 17876
rect 25590 17864 25596 17876
rect 24176 17836 25596 17864
rect 24176 17824 24182 17836
rect 25590 17824 25596 17836
rect 25648 17824 25654 17876
rect 25958 17824 25964 17876
rect 26016 17824 26022 17876
rect 26142 17824 26148 17876
rect 26200 17864 26206 17876
rect 27338 17864 27344 17876
rect 26200 17836 27344 17864
rect 26200 17824 26206 17836
rect 27338 17824 27344 17836
rect 27396 17824 27402 17876
rect 27430 17824 27436 17876
rect 27488 17864 27494 17876
rect 27801 17867 27859 17873
rect 27801 17864 27813 17867
rect 27488 17836 27813 17864
rect 27488 17824 27494 17836
rect 27801 17833 27813 17836
rect 27847 17833 27859 17867
rect 27801 17827 27859 17833
rect 30558 17824 30564 17876
rect 30616 17864 30622 17876
rect 31297 17867 31355 17873
rect 31297 17864 31309 17867
rect 30616 17836 31309 17864
rect 30616 17824 30622 17836
rect 31297 17833 31309 17836
rect 31343 17833 31355 17867
rect 31297 17827 31355 17833
rect 23474 17796 23480 17808
rect 22848 17768 23480 17796
rect 22848 17737 22876 17768
rect 23474 17756 23480 17768
rect 23532 17756 23538 17808
rect 24026 17796 24032 17808
rect 23584 17768 24032 17796
rect 20303 17700 20760 17728
rect 22833 17731 22891 17737
rect 20303 17697 20315 17700
rect 20257 17691 20315 17697
rect 22833 17697 22845 17731
rect 22879 17697 22891 17731
rect 23014 17728 23020 17740
rect 22975 17700 23020 17728
rect 22833 17691 22891 17697
rect 23014 17688 23020 17700
rect 23072 17688 23078 17740
rect 12161 17663 12219 17669
rect 12161 17629 12173 17663
rect 12207 17660 12219 17663
rect 12345 17663 12403 17669
rect 12345 17660 12357 17663
rect 12207 17632 12357 17660
rect 12207 17629 12219 17632
rect 12161 17623 12219 17629
rect 12345 17629 12357 17632
rect 12391 17629 12403 17663
rect 12345 17623 12403 17629
rect 12529 17663 12587 17669
rect 12529 17629 12541 17663
rect 12575 17660 12587 17663
rect 12805 17663 12863 17669
rect 12805 17660 12817 17663
rect 12575 17632 12817 17660
rect 12575 17629 12587 17632
rect 12529 17623 12587 17629
rect 12805 17629 12817 17632
rect 12851 17629 12863 17663
rect 12805 17623 12863 17629
rect 13081 17663 13139 17669
rect 13081 17629 13093 17663
rect 13127 17629 13139 17663
rect 13081 17623 13139 17629
rect 13265 17663 13323 17669
rect 13265 17629 13277 17663
rect 13311 17660 13323 17663
rect 13906 17660 13912 17672
rect 13311 17632 13912 17660
rect 13311 17629 13323 17632
rect 13265 17623 13323 17629
rect 13906 17620 13912 17632
rect 13964 17620 13970 17672
rect 14458 17620 14464 17672
rect 14516 17660 14522 17672
rect 15010 17660 15016 17672
rect 14516 17632 15016 17660
rect 14516 17620 14522 17632
rect 15010 17620 15016 17632
rect 15068 17620 15074 17672
rect 15289 17663 15347 17669
rect 15289 17629 15301 17663
rect 15335 17629 15347 17663
rect 15470 17660 15476 17672
rect 15431 17632 15476 17660
rect 15289 17623 15347 17629
rect 12253 17595 12311 17601
rect 11716 17564 11836 17592
rect 11333 17555 11391 17561
rect 3568 17496 7052 17524
rect 7101 17527 7159 17533
rect 3568 17484 3574 17496
rect 7101 17493 7113 17527
rect 7147 17524 7159 17527
rect 7190 17524 7196 17536
rect 7147 17496 7196 17524
rect 7147 17493 7159 17496
rect 7101 17487 7159 17493
rect 7190 17484 7196 17496
rect 7248 17484 7254 17536
rect 7929 17527 7987 17533
rect 7929 17493 7941 17527
rect 7975 17524 7987 17527
rect 8662 17524 8668 17536
rect 7975 17496 8668 17524
rect 7975 17493 7987 17496
rect 7929 17487 7987 17493
rect 8662 17484 8668 17496
rect 8720 17484 8726 17536
rect 8938 17484 8944 17536
rect 8996 17524 9002 17536
rect 10597 17527 10655 17533
rect 10597 17524 10609 17527
rect 8996 17496 10609 17524
rect 8996 17484 9002 17496
rect 10597 17493 10609 17496
rect 10643 17524 10655 17527
rect 11425 17527 11483 17533
rect 11425 17524 11437 17527
rect 10643 17496 11437 17524
rect 10643 17493 10655 17496
rect 10597 17487 10655 17493
rect 11425 17493 11437 17496
rect 11471 17493 11483 17527
rect 11425 17487 11483 17493
rect 11517 17527 11575 17533
rect 11517 17493 11529 17527
rect 11563 17524 11575 17527
rect 11698 17524 11704 17536
rect 11563 17496 11704 17524
rect 11563 17493 11575 17496
rect 11517 17487 11575 17493
rect 11698 17484 11704 17496
rect 11756 17484 11762 17536
rect 11808 17524 11836 17564
rect 12253 17561 12265 17595
rect 12299 17592 12311 17595
rect 14090 17592 14096 17604
rect 12299 17564 14096 17592
rect 12299 17561 12311 17564
rect 12253 17555 12311 17561
rect 14090 17552 14096 17564
rect 14148 17552 14154 17604
rect 14185 17595 14243 17601
rect 14185 17561 14197 17595
rect 14231 17561 14243 17595
rect 14826 17592 14832 17604
rect 14787 17564 14832 17592
rect 14185 17555 14243 17561
rect 12529 17527 12587 17533
rect 12529 17524 12541 17527
rect 11808 17496 12541 17524
rect 12529 17493 12541 17496
rect 12575 17493 12587 17527
rect 12529 17487 12587 17493
rect 12621 17527 12679 17533
rect 12621 17493 12633 17527
rect 12667 17524 12679 17527
rect 13998 17524 14004 17536
rect 12667 17496 14004 17524
rect 12667 17493 12679 17496
rect 12621 17487 12679 17493
rect 13998 17484 14004 17496
rect 14056 17484 14062 17536
rect 14200 17524 14228 17555
rect 14826 17552 14832 17564
rect 14884 17552 14890 17604
rect 15304 17592 15332 17623
rect 15470 17620 15476 17632
rect 15528 17660 15534 17672
rect 16666 17660 16672 17672
rect 15528 17632 16672 17660
rect 15528 17620 15534 17632
rect 16666 17620 16672 17632
rect 16724 17620 16730 17672
rect 16761 17663 16819 17669
rect 16761 17629 16773 17663
rect 16807 17660 16819 17663
rect 17611 17660 17724 17670
rect 17957 17663 18015 17669
rect 16807 17642 17917 17660
rect 16807 17632 17639 17642
rect 17696 17632 17917 17642
rect 16807 17629 16819 17632
rect 16761 17623 16819 17629
rect 15378 17592 15384 17604
rect 15291 17564 15384 17592
rect 15378 17552 15384 17564
rect 15436 17592 15442 17604
rect 15838 17592 15844 17604
rect 15436 17564 15844 17592
rect 15436 17552 15442 17564
rect 15838 17552 15844 17564
rect 15896 17552 15902 17604
rect 15930 17552 15936 17604
rect 15988 17592 15994 17604
rect 16942 17592 16948 17604
rect 15988 17564 16948 17592
rect 15988 17552 15994 17564
rect 16942 17552 16948 17564
rect 17000 17552 17006 17604
rect 17889 17592 17917 17632
rect 17957 17629 17969 17663
rect 18003 17660 18015 17663
rect 18046 17660 18052 17672
rect 18003 17632 18052 17660
rect 18003 17629 18015 17632
rect 17957 17623 18015 17629
rect 18046 17620 18052 17632
rect 18104 17620 18110 17672
rect 18230 17660 18236 17672
rect 18191 17632 18236 17660
rect 18230 17620 18236 17632
rect 18288 17620 18294 17672
rect 19978 17660 19984 17672
rect 19939 17632 19984 17660
rect 19978 17620 19984 17632
rect 20036 17620 20042 17672
rect 20162 17660 20168 17672
rect 20123 17632 20168 17660
rect 20162 17620 20168 17632
rect 20220 17620 20226 17672
rect 20717 17663 20775 17669
rect 20717 17629 20729 17663
rect 20763 17660 20775 17663
rect 21910 17660 21916 17672
rect 20763 17632 21916 17660
rect 20763 17629 20775 17632
rect 20717 17623 20775 17629
rect 21910 17620 21916 17632
rect 21968 17620 21974 17672
rect 22554 17620 22560 17672
rect 22612 17660 22618 17672
rect 23584 17669 23612 17768
rect 24026 17756 24032 17768
rect 24084 17796 24090 17808
rect 25976 17796 26004 17824
rect 24084 17768 26004 17796
rect 24084 17756 24090 17768
rect 26602 17756 26608 17808
rect 26660 17796 26666 17808
rect 28626 17796 28632 17808
rect 26660 17768 28632 17796
rect 26660 17756 26666 17768
rect 28626 17756 28632 17768
rect 28684 17756 28690 17808
rect 25498 17728 25504 17740
rect 24872 17700 25504 17728
rect 22741 17663 22799 17669
rect 22741 17660 22753 17663
rect 22612 17632 22753 17660
rect 22612 17620 22618 17632
rect 22741 17629 22753 17632
rect 22787 17629 22799 17663
rect 22741 17623 22799 17629
rect 22925 17663 22983 17669
rect 22925 17629 22937 17663
rect 22971 17660 22983 17663
rect 23201 17663 23259 17669
rect 23201 17660 23213 17663
rect 22971 17632 23213 17660
rect 22971 17629 22983 17632
rect 22925 17623 22983 17629
rect 23201 17629 23213 17632
rect 23247 17629 23259 17663
rect 23201 17623 23259 17629
rect 23569 17663 23627 17669
rect 23569 17629 23581 17663
rect 23615 17629 23627 17663
rect 24578 17660 24584 17672
rect 24539 17632 24584 17660
rect 23569 17623 23627 17629
rect 24578 17620 24584 17632
rect 24636 17620 24642 17672
rect 24872 17669 24900 17700
rect 25498 17688 25504 17700
rect 25556 17688 25562 17740
rect 26694 17688 26700 17740
rect 26752 17728 26758 17740
rect 27985 17731 28043 17737
rect 27985 17728 27997 17731
rect 26752 17700 27997 17728
rect 26752 17688 26758 17700
rect 27985 17697 27997 17700
rect 28031 17697 28043 17731
rect 29914 17728 29920 17740
rect 29875 17700 29920 17728
rect 27985 17691 28043 17697
rect 29914 17688 29920 17700
rect 29972 17688 29978 17740
rect 24857 17663 24915 17669
rect 24857 17629 24869 17663
rect 24903 17629 24915 17663
rect 25038 17660 25044 17672
rect 24999 17632 25044 17660
rect 24857 17623 24915 17629
rect 25038 17620 25044 17632
rect 25096 17620 25102 17672
rect 26050 17620 26056 17672
rect 26108 17660 26114 17672
rect 27709 17663 27767 17669
rect 27709 17660 27721 17663
rect 26108 17632 27721 17660
rect 26108 17620 26114 17632
rect 27709 17629 27721 17632
rect 27755 17629 27767 17663
rect 27709 17623 27767 17629
rect 19797 17595 19855 17601
rect 17889 17564 19748 17592
rect 15102 17524 15108 17536
rect 14200 17496 15108 17524
rect 15102 17484 15108 17496
rect 15160 17484 15166 17536
rect 17126 17484 17132 17536
rect 17184 17524 17190 17536
rect 17589 17527 17647 17533
rect 17589 17524 17601 17527
rect 17184 17496 17601 17524
rect 17184 17484 17190 17496
rect 17589 17493 17601 17496
rect 17635 17493 17647 17527
rect 17589 17487 17647 17493
rect 17678 17484 17684 17536
rect 17736 17524 17742 17536
rect 17736 17496 17781 17524
rect 17736 17484 17742 17496
rect 18966 17484 18972 17536
rect 19024 17524 19030 17536
rect 19334 17524 19340 17536
rect 19024 17496 19340 17524
rect 19024 17484 19030 17496
rect 19334 17484 19340 17496
rect 19392 17484 19398 17536
rect 19720 17524 19748 17564
rect 19797 17561 19809 17595
rect 19843 17592 19855 17595
rect 20962 17595 21020 17601
rect 20962 17592 20974 17595
rect 19843 17564 20974 17592
rect 19843 17561 19855 17564
rect 19797 17555 19855 17561
rect 20962 17561 20974 17564
rect 21008 17561 21020 17595
rect 25501 17595 25559 17601
rect 25501 17592 25513 17595
rect 20962 17555 21020 17561
rect 22066 17564 25513 17592
rect 20346 17524 20352 17536
rect 19720 17496 20352 17524
rect 20346 17484 20352 17496
rect 20404 17484 20410 17536
rect 20622 17484 20628 17536
rect 20680 17524 20686 17536
rect 22066 17524 22094 17564
rect 25501 17561 25513 17564
rect 25547 17592 25559 17595
rect 26142 17592 26148 17604
rect 25547 17564 26148 17592
rect 25547 17561 25559 17564
rect 25501 17555 25559 17561
rect 26142 17552 26148 17564
rect 26200 17552 26206 17604
rect 27798 17552 27804 17604
rect 27856 17592 27862 17604
rect 28813 17595 28871 17601
rect 28813 17592 28825 17595
rect 27856 17564 28825 17592
rect 27856 17552 27862 17564
rect 28813 17561 28825 17564
rect 28859 17561 28871 17595
rect 28813 17555 28871 17561
rect 28997 17595 29055 17601
rect 28997 17561 29009 17595
rect 29043 17592 29055 17595
rect 29270 17592 29276 17604
rect 29043 17564 29276 17592
rect 29043 17561 29055 17564
rect 28997 17555 29055 17561
rect 29270 17552 29276 17564
rect 29328 17552 29334 17604
rect 30184 17595 30242 17601
rect 30184 17561 30196 17595
rect 30230 17592 30242 17595
rect 30558 17592 30564 17604
rect 30230 17564 30564 17592
rect 30230 17561 30242 17564
rect 30184 17555 30242 17561
rect 30558 17552 30564 17564
rect 30616 17552 30622 17604
rect 20680 17496 22094 17524
rect 22557 17527 22615 17533
rect 20680 17484 20686 17496
rect 22557 17493 22569 17527
rect 22603 17524 22615 17527
rect 23014 17524 23020 17536
rect 22603 17496 23020 17524
rect 22603 17493 22615 17496
rect 22557 17487 22615 17493
rect 23014 17484 23020 17496
rect 23072 17484 23078 17536
rect 24210 17484 24216 17536
rect 24268 17524 24274 17536
rect 24397 17527 24455 17533
rect 24397 17524 24409 17527
rect 24268 17496 24409 17524
rect 24268 17484 24274 17496
rect 24397 17493 24409 17496
rect 24443 17493 24455 17527
rect 24397 17487 24455 17493
rect 24946 17484 24952 17536
rect 25004 17524 25010 17536
rect 25774 17524 25780 17536
rect 25004 17496 25780 17524
rect 25004 17484 25010 17496
rect 25774 17484 25780 17496
rect 25832 17524 25838 17536
rect 26789 17527 26847 17533
rect 26789 17524 26801 17527
rect 25832 17496 26801 17524
rect 25832 17484 25838 17496
rect 26789 17493 26801 17496
rect 26835 17524 26847 17527
rect 27614 17524 27620 17536
rect 26835 17496 27620 17524
rect 26835 17493 26847 17496
rect 26789 17487 26847 17493
rect 27614 17484 27620 17496
rect 27672 17484 27678 17536
rect 28258 17524 28264 17536
rect 28219 17496 28264 17524
rect 28258 17484 28264 17496
rect 28316 17484 28322 17536
rect 1104 17434 32016 17456
rect 768 17360 888 17388
rect 1104 17382 7288 17434
rect 7340 17382 17592 17434
rect 17644 17382 27896 17434
rect 27948 17382 32016 17434
rect 1104 17360 32016 17382
rect 0 17252 800 17266
rect 860 17252 888 17360
rect 0 17224 888 17252
rect 1504 17292 3832 17320
rect 0 17210 800 17224
rect 1504 17193 1532 17292
rect 2777 17255 2835 17261
rect 1688 17224 2360 17252
rect 1688 17193 1716 17224
rect 2332 17193 2360 17224
rect 2777 17221 2789 17255
rect 2823 17252 2835 17255
rect 3510 17252 3516 17264
rect 2823 17224 3516 17252
rect 2823 17221 2835 17224
rect 2777 17215 2835 17221
rect 3510 17212 3516 17224
rect 3568 17212 3574 17264
rect 1489 17187 1547 17193
rect 1489 17153 1501 17187
rect 1535 17153 1547 17187
rect 1489 17147 1547 17153
rect 1673 17187 1731 17193
rect 1673 17153 1685 17187
rect 1719 17153 1731 17187
rect 1673 17147 1731 17153
rect 2133 17187 2191 17193
rect 2133 17153 2145 17187
rect 2179 17153 2191 17187
rect 2133 17147 2191 17153
rect 2317 17187 2375 17193
rect 2317 17153 2329 17187
rect 2363 17184 2375 17187
rect 2682 17184 2688 17196
rect 2363 17156 2688 17184
rect 2363 17153 2375 17156
rect 2317 17147 2375 17153
rect 2148 17116 2176 17147
rect 2682 17144 2688 17156
rect 2740 17144 2746 17196
rect 3804 17184 3832 17292
rect 3878 17280 3884 17332
rect 3936 17320 3942 17332
rect 4065 17323 4123 17329
rect 4065 17320 4077 17323
rect 3936 17292 4077 17320
rect 3936 17280 3942 17292
rect 4065 17289 4077 17292
rect 4111 17289 4123 17323
rect 5442 17320 5448 17332
rect 5403 17292 5448 17320
rect 4065 17283 4123 17289
rect 5442 17280 5448 17292
rect 5500 17280 5506 17332
rect 7101 17323 7159 17329
rect 7101 17289 7113 17323
rect 7147 17320 7159 17323
rect 7190 17320 7196 17332
rect 7147 17292 7196 17320
rect 7147 17289 7159 17292
rect 7101 17283 7159 17289
rect 7190 17280 7196 17292
rect 7248 17280 7254 17332
rect 7285 17323 7343 17329
rect 7285 17289 7297 17323
rect 7331 17320 7343 17323
rect 7926 17320 7932 17332
rect 7331 17292 7932 17320
rect 7331 17289 7343 17292
rect 7285 17283 7343 17289
rect 7926 17280 7932 17292
rect 7984 17280 7990 17332
rect 8018 17280 8024 17332
rect 8076 17320 8082 17332
rect 8113 17323 8171 17329
rect 8113 17320 8125 17323
rect 8076 17292 8125 17320
rect 8076 17280 8082 17292
rect 8113 17289 8125 17292
rect 8159 17320 8171 17323
rect 10873 17323 10931 17329
rect 10873 17320 10885 17323
rect 8159 17292 10885 17320
rect 8159 17289 8171 17292
rect 8113 17283 8171 17289
rect 10873 17289 10885 17292
rect 10919 17289 10931 17323
rect 10873 17283 10931 17289
rect 11517 17323 11575 17329
rect 11517 17289 11529 17323
rect 11563 17320 11575 17323
rect 11606 17320 11612 17332
rect 11563 17292 11612 17320
rect 11563 17289 11575 17292
rect 11517 17283 11575 17289
rect 11606 17280 11612 17292
rect 11664 17280 11670 17332
rect 17221 17323 17279 17329
rect 17221 17320 17233 17323
rect 12406 17292 17233 17320
rect 4982 17252 4988 17264
rect 4943 17224 4988 17252
rect 4982 17212 4988 17224
rect 5040 17212 5046 17264
rect 12406 17252 12434 17292
rect 17221 17289 17233 17292
rect 17267 17289 17279 17323
rect 17221 17283 17279 17289
rect 17678 17280 17684 17332
rect 17736 17320 17742 17332
rect 18046 17320 18052 17332
rect 17736 17292 18052 17320
rect 17736 17280 17742 17292
rect 18046 17280 18052 17292
rect 18104 17280 18110 17332
rect 18138 17280 18144 17332
rect 18196 17320 18202 17332
rect 18690 17320 18696 17332
rect 18196 17292 18696 17320
rect 18196 17280 18202 17292
rect 18690 17280 18696 17292
rect 18748 17280 18754 17332
rect 18969 17323 19027 17329
rect 18969 17289 18981 17323
rect 19015 17320 19027 17323
rect 19150 17320 19156 17332
rect 19015 17292 19156 17320
rect 19015 17289 19027 17292
rect 18969 17283 19027 17289
rect 19150 17280 19156 17292
rect 19208 17280 19214 17332
rect 19978 17280 19984 17332
rect 20036 17320 20042 17332
rect 20165 17323 20223 17329
rect 20165 17320 20177 17323
rect 20036 17292 20177 17320
rect 20036 17280 20042 17292
rect 20165 17289 20177 17292
rect 20211 17289 20223 17323
rect 20165 17283 20223 17289
rect 22373 17323 22431 17329
rect 22373 17289 22385 17323
rect 22419 17320 22431 17323
rect 22554 17320 22560 17332
rect 22419 17292 22560 17320
rect 22419 17289 22431 17292
rect 22373 17283 22431 17289
rect 22554 17280 22560 17292
rect 22612 17280 22618 17332
rect 23106 17320 23112 17332
rect 23067 17292 23112 17320
rect 23106 17280 23112 17292
rect 23164 17280 23170 17332
rect 23198 17280 23204 17332
rect 23256 17320 23262 17332
rect 24029 17323 24087 17329
rect 23256 17292 23428 17320
rect 23256 17280 23262 17292
rect 13814 17252 13820 17264
rect 7208 17224 12434 17252
rect 12544 17224 13820 17252
rect 7208 17184 7236 17224
rect 3804 17156 7236 17184
rect 7742 17144 7748 17196
rect 7800 17184 7806 17196
rect 8205 17187 8263 17193
rect 8205 17184 8217 17187
rect 7800 17156 8217 17184
rect 7800 17144 7806 17156
rect 8205 17153 8217 17156
rect 8251 17153 8263 17187
rect 8938 17184 8944 17196
rect 8899 17156 8944 17184
rect 8205 17147 8263 17153
rect 8938 17144 8944 17156
rect 8996 17144 9002 17196
rect 9214 17193 9220 17196
rect 9208 17184 9220 17193
rect 9175 17156 9220 17184
rect 9208 17147 9220 17156
rect 9214 17144 9220 17147
rect 9272 17144 9278 17196
rect 9490 17144 9496 17196
rect 9548 17184 9554 17196
rect 10781 17187 10839 17193
rect 10781 17184 10793 17187
rect 9548 17156 10793 17184
rect 9548 17144 9554 17156
rect 10781 17153 10793 17156
rect 10827 17153 10839 17187
rect 11698 17184 11704 17196
rect 11659 17156 11704 17184
rect 10781 17147 10839 17153
rect 11698 17144 11704 17156
rect 11756 17144 11762 17196
rect 12544 17193 12572 17224
rect 13814 17212 13820 17224
rect 13872 17212 13878 17264
rect 13998 17212 14004 17264
rect 14056 17252 14062 17264
rect 14056 17224 14596 17252
rect 14056 17212 14062 17224
rect 14568 17193 14596 17224
rect 15378 17212 15384 17264
rect 15436 17252 15442 17264
rect 15436 17224 16160 17252
rect 15436 17212 15442 17224
rect 12529 17187 12587 17193
rect 12529 17153 12541 17187
rect 12575 17153 12587 17187
rect 12529 17147 12587 17153
rect 12796 17187 12854 17193
rect 12796 17153 12808 17187
rect 12842 17184 12854 17187
rect 14369 17187 14427 17193
rect 14369 17184 14381 17187
rect 12842 17156 14381 17184
rect 12842 17153 12854 17156
rect 12796 17147 12854 17153
rect 14369 17153 14381 17156
rect 14415 17153 14427 17187
rect 14369 17147 14427 17153
rect 14553 17187 14611 17193
rect 14553 17153 14565 17187
rect 14599 17153 14611 17187
rect 14553 17147 14611 17153
rect 14734 17144 14740 17196
rect 14792 17184 14798 17196
rect 14829 17187 14887 17193
rect 14829 17184 14841 17187
rect 14792 17156 14841 17184
rect 14792 17144 14798 17156
rect 14829 17153 14841 17156
rect 14875 17153 14887 17187
rect 14829 17147 14887 17153
rect 15010 17144 15016 17196
rect 15068 17184 15074 17196
rect 15657 17187 15715 17193
rect 15657 17184 15669 17187
rect 15068 17156 15669 17184
rect 15068 17144 15074 17156
rect 15657 17153 15669 17156
rect 15703 17153 15715 17187
rect 15657 17147 15715 17153
rect 15838 17144 15844 17196
rect 15896 17184 15902 17196
rect 16132 17193 16160 17224
rect 16592 17224 16804 17252
rect 15933 17187 15991 17193
rect 15933 17184 15945 17187
rect 15896 17156 15945 17184
rect 15896 17144 15902 17156
rect 15933 17153 15945 17156
rect 15979 17153 15991 17187
rect 15933 17147 15991 17153
rect 16117 17187 16175 17193
rect 16117 17153 16129 17187
rect 16163 17153 16175 17187
rect 16117 17147 16175 17153
rect 8389 17119 8447 17125
rect 2148 17088 7788 17116
rect 1854 17008 1860 17060
rect 1912 17048 1918 17060
rect 3878 17048 3884 17060
rect 1912 17020 3884 17048
rect 1912 17008 1918 17020
rect 3878 17008 3884 17020
rect 3936 17008 3942 17060
rect 5166 17008 5172 17060
rect 5224 17048 5230 17060
rect 5261 17051 5319 17057
rect 5261 17048 5273 17051
rect 5224 17020 5273 17048
rect 5224 17008 5230 17020
rect 5261 17017 5273 17020
rect 5307 17017 5319 17051
rect 6733 17051 6791 17057
rect 5261 17011 5319 17017
rect 5368 17020 5580 17048
rect 1489 16983 1547 16989
rect 1489 16949 1501 16983
rect 1535 16980 1547 16983
rect 1762 16980 1768 16992
rect 1535 16952 1768 16980
rect 1535 16949 1547 16952
rect 1489 16943 1547 16949
rect 1762 16940 1768 16952
rect 1820 16940 1826 16992
rect 2133 16983 2191 16989
rect 2133 16949 2145 16983
rect 2179 16980 2191 16983
rect 5368 16980 5396 17020
rect 2179 16952 5396 16980
rect 5552 16980 5580 17020
rect 6733 17017 6745 17051
rect 6779 17048 6791 17051
rect 7466 17048 7472 17060
rect 6779 17020 7472 17048
rect 6779 17017 6791 17020
rect 6733 17011 6791 17017
rect 7466 17008 7472 17020
rect 7524 17008 7530 17060
rect 7760 17057 7788 17088
rect 8389 17085 8401 17119
rect 8435 17116 8447 17119
rect 8478 17116 8484 17128
rect 8435 17088 8484 17116
rect 8435 17085 8447 17088
rect 8389 17079 8447 17085
rect 8478 17076 8484 17088
rect 8536 17076 8542 17128
rect 10594 17076 10600 17128
rect 10652 17116 10658 17128
rect 11977 17119 12035 17125
rect 11977 17116 11989 17119
rect 10652 17088 11989 17116
rect 10652 17076 10658 17088
rect 11977 17085 11989 17088
rect 12023 17085 12035 17119
rect 11977 17079 12035 17085
rect 13538 17076 13544 17128
rect 13596 17116 13602 17128
rect 15473 17119 15531 17125
rect 13596 17088 14872 17116
rect 13596 17076 13602 17088
rect 7745 17051 7803 17057
rect 7745 17017 7757 17051
rect 7791 17017 7803 17051
rect 7745 17011 7803 17017
rect 8018 17008 8024 17060
rect 8076 17048 8082 17060
rect 8202 17048 8208 17060
rect 8076 17020 8208 17048
rect 8076 17008 8082 17020
rect 8202 17008 8208 17020
rect 8260 17008 8266 17060
rect 10226 17008 10232 17060
rect 10284 17048 10290 17060
rect 12250 17048 12256 17060
rect 10284 17020 12256 17048
rect 10284 17008 10290 17020
rect 12250 17008 12256 17020
rect 12308 17008 12314 17060
rect 14737 17051 14795 17057
rect 14737 17048 14749 17051
rect 13464 17020 14749 17048
rect 7006 16980 7012 16992
rect 5552 16952 7012 16980
rect 2179 16949 2191 16952
rect 2133 16943 2191 16949
rect 7006 16940 7012 16952
rect 7064 16940 7070 16992
rect 7101 16983 7159 16989
rect 7101 16949 7113 16983
rect 7147 16980 7159 16983
rect 7374 16980 7380 16992
rect 7147 16952 7380 16980
rect 7147 16949 7159 16952
rect 7101 16943 7159 16949
rect 7374 16940 7380 16952
rect 7432 16940 7438 16992
rect 7484 16980 7512 17008
rect 8386 16980 8392 16992
rect 7484 16952 8392 16980
rect 8386 16940 8392 16952
rect 8444 16940 8450 16992
rect 9674 16940 9680 16992
rect 9732 16980 9738 16992
rect 10321 16983 10379 16989
rect 10321 16980 10333 16983
rect 9732 16952 10333 16980
rect 9732 16940 9738 16952
rect 10321 16949 10333 16952
rect 10367 16980 10379 16983
rect 10870 16980 10876 16992
rect 10367 16952 10876 16980
rect 10367 16949 10379 16952
rect 10321 16943 10379 16949
rect 10870 16940 10876 16952
rect 10928 16940 10934 16992
rect 11882 16980 11888 16992
rect 11795 16952 11888 16980
rect 11882 16940 11888 16952
rect 11940 16980 11946 16992
rect 12158 16980 12164 16992
rect 11940 16952 12164 16980
rect 11940 16940 11946 16952
rect 12158 16940 12164 16952
rect 12216 16980 12222 16992
rect 13464 16980 13492 17020
rect 14737 17017 14749 17020
rect 14783 17017 14795 17051
rect 14844 17048 14872 17088
rect 15473 17085 15485 17119
rect 15519 17116 15531 17119
rect 16592 17116 16620 17224
rect 16666 17144 16672 17196
rect 16724 17144 16730 17196
rect 16776 17184 16804 17224
rect 17126 17212 17132 17264
rect 17184 17252 17190 17264
rect 17402 17252 17408 17264
rect 17184 17224 17408 17252
rect 17184 17212 17190 17224
rect 17402 17212 17408 17224
rect 17460 17212 17466 17264
rect 17862 17261 17868 17264
rect 17497 17255 17555 17261
rect 17497 17221 17509 17255
rect 17543 17252 17555 17255
rect 17856 17252 17868 17261
rect 17543 17224 17632 17252
rect 17823 17224 17868 17252
rect 17543 17221 17555 17224
rect 17497 17215 17555 17221
rect 16853 17187 16911 17193
rect 16853 17184 16865 17187
rect 16776 17156 16865 17184
rect 16853 17153 16865 17156
rect 16899 17153 16911 17187
rect 17034 17184 17040 17196
rect 16995 17156 17040 17184
rect 16853 17147 16911 17153
rect 17034 17144 17040 17156
rect 17092 17144 17098 17196
rect 17604 17193 17632 17224
rect 17856 17215 17868 17224
rect 17862 17212 17868 17215
rect 17920 17212 17926 17264
rect 17954 17212 17960 17264
rect 18012 17252 18018 17264
rect 19705 17255 19763 17261
rect 19705 17252 19717 17255
rect 18012 17224 19717 17252
rect 18012 17212 18018 17224
rect 19705 17221 19717 17224
rect 19751 17221 19763 17255
rect 19705 17215 19763 17221
rect 17596 17187 17654 17193
rect 17596 17153 17608 17187
rect 17642 17153 17654 17187
rect 17596 17147 17654 17153
rect 17687 17184 17816 17190
rect 17687 17162 18644 17184
rect 15519 17088 16620 17116
rect 16684 17116 16712 17144
rect 17129 17119 17187 17125
rect 17129 17116 17141 17119
rect 16684 17088 17141 17116
rect 15519 17085 15531 17088
rect 15473 17079 15531 17085
rect 17129 17085 17141 17088
rect 17175 17085 17187 17119
rect 17129 17079 17187 17085
rect 17221 17119 17279 17125
rect 17221 17085 17233 17119
rect 17267 17116 17279 17119
rect 17687 17116 17715 17162
rect 17788 17156 18644 17162
rect 17267 17088 17715 17116
rect 18616 17116 18644 17156
rect 18874 17144 18880 17196
rect 18932 17184 18938 17196
rect 19521 17187 19579 17193
rect 19521 17184 19533 17187
rect 18932 17156 19533 17184
rect 18932 17144 18938 17156
rect 19521 17153 19533 17156
rect 19567 17153 19579 17187
rect 19521 17147 19579 17153
rect 19720 17116 19748 17215
rect 19794 17212 19800 17264
rect 19852 17252 19858 17264
rect 19852 17224 20668 17252
rect 19852 17212 19858 17224
rect 19996 17196 20024 17224
rect 19978 17144 19984 17196
rect 20036 17144 20042 17196
rect 20346 17184 20352 17196
rect 20307 17156 20352 17184
rect 20346 17144 20352 17156
rect 20404 17144 20410 17196
rect 20640 17193 20668 17224
rect 21818 17212 21824 17264
rect 21876 17252 21882 17264
rect 23400 17252 23428 17292
rect 24029 17289 24041 17323
rect 24075 17320 24087 17323
rect 24302 17320 24308 17332
rect 24075 17292 24308 17320
rect 24075 17289 24087 17292
rect 24029 17283 24087 17289
rect 24302 17280 24308 17292
rect 24360 17280 24366 17332
rect 26973 17323 27031 17329
rect 26973 17289 26985 17323
rect 27019 17320 27031 17323
rect 27154 17320 27160 17332
rect 27019 17292 27160 17320
rect 27019 17289 27031 17292
rect 26973 17283 27031 17289
rect 27154 17280 27160 17292
rect 27212 17280 27218 17332
rect 29086 17280 29092 17332
rect 29144 17320 29150 17332
rect 29144 17292 29868 17320
rect 29144 17280 29150 17292
rect 24670 17252 24676 17264
rect 21876 17224 23336 17252
rect 23400 17224 24676 17252
rect 21876 17212 21882 17224
rect 20625 17187 20683 17193
rect 20625 17153 20637 17187
rect 20671 17153 20683 17187
rect 20625 17147 20683 17153
rect 20809 17187 20867 17193
rect 20809 17153 20821 17187
rect 20855 17184 20867 17187
rect 21726 17184 21732 17196
rect 20855 17156 21732 17184
rect 20855 17153 20867 17156
rect 20809 17147 20867 17153
rect 21726 17144 21732 17156
rect 21784 17144 21790 17196
rect 22005 17187 22063 17193
rect 22005 17153 22017 17187
rect 22051 17153 22063 17187
rect 22186 17184 22192 17196
rect 22147 17156 22192 17184
rect 22005 17147 22063 17153
rect 20714 17116 20720 17128
rect 18616 17088 19012 17116
rect 19720 17088 20720 17116
rect 17267 17085 17279 17088
rect 17221 17079 17279 17085
rect 15746 17048 15752 17060
rect 14844 17020 15752 17048
rect 14737 17011 14795 17017
rect 15746 17008 15752 17020
rect 15804 17008 15810 17060
rect 16669 17051 16727 17057
rect 16669 17048 16681 17051
rect 15856 17020 16681 17048
rect 13906 16980 13912 16992
rect 12216 16952 13492 16980
rect 13867 16952 13912 16980
rect 12216 16940 12222 16952
rect 13906 16940 13912 16952
rect 13964 16940 13970 16992
rect 15470 16940 15476 16992
rect 15528 16980 15534 16992
rect 15856 16980 15884 17020
rect 16669 17017 16681 17020
rect 16715 17017 16727 17051
rect 16669 17011 16727 17017
rect 16942 17008 16948 17060
rect 17000 17048 17006 17060
rect 17402 17048 17408 17060
rect 17000 17020 17408 17048
rect 17000 17008 17006 17020
rect 17402 17008 17408 17020
rect 17460 17048 17466 17060
rect 17497 17051 17555 17057
rect 17497 17048 17509 17051
rect 17460 17020 17509 17048
rect 17460 17008 17466 17020
rect 17497 17017 17509 17020
rect 17543 17017 17555 17051
rect 17497 17011 17555 17017
rect 15528 16952 15884 16980
rect 15528 16940 15534 16952
rect 16206 16940 16212 16992
rect 16264 16980 16270 16992
rect 18874 16980 18880 16992
rect 16264 16952 18880 16980
rect 16264 16940 16270 16952
rect 18874 16940 18880 16952
rect 18932 16940 18938 16992
rect 18984 16980 19012 17088
rect 20714 17076 20720 17088
rect 20772 17076 20778 17128
rect 20898 17076 20904 17128
rect 20956 17116 20962 17128
rect 22020 17116 22048 17147
rect 22186 17144 22192 17156
rect 22244 17144 22250 17196
rect 23308 17193 23336 17224
rect 24670 17212 24676 17224
rect 24728 17212 24734 17264
rect 27246 17212 27252 17264
rect 27304 17252 27310 17264
rect 27862 17255 27920 17261
rect 27862 17252 27874 17255
rect 27304 17224 27874 17252
rect 27304 17212 27310 17224
rect 27862 17221 27874 17224
rect 27908 17221 27920 17255
rect 27862 17215 27920 17221
rect 29840 17196 29868 17292
rect 30834 17252 30840 17264
rect 30300 17224 30840 17252
rect 23293 17187 23351 17193
rect 23293 17153 23305 17187
rect 23339 17153 23351 17187
rect 24210 17184 24216 17196
rect 24171 17156 24216 17184
rect 23293 17147 23351 17153
rect 24210 17144 24216 17156
rect 24268 17144 24274 17196
rect 24486 17184 24492 17196
rect 24447 17156 24492 17184
rect 24486 17144 24492 17156
rect 24544 17144 24550 17196
rect 24854 17144 24860 17196
rect 24912 17184 24918 17196
rect 25205 17187 25263 17193
rect 25205 17184 25217 17187
rect 24912 17156 25217 17184
rect 24912 17144 24918 17156
rect 25205 17153 25217 17156
rect 25251 17153 25263 17187
rect 25205 17147 25263 17153
rect 26602 17144 26608 17196
rect 26660 17184 26666 17196
rect 27157 17187 27215 17193
rect 27157 17184 27169 17187
rect 26660 17156 27169 17184
rect 26660 17144 26666 17156
rect 27157 17153 27169 17156
rect 27203 17153 27215 17187
rect 27614 17184 27620 17196
rect 27575 17156 27620 17184
rect 27157 17147 27215 17153
rect 27614 17144 27620 17156
rect 27672 17144 27678 17196
rect 29086 17144 29092 17196
rect 29144 17184 29150 17196
rect 29641 17187 29699 17193
rect 29641 17184 29653 17187
rect 29144 17156 29653 17184
rect 29144 17144 29150 17156
rect 29641 17153 29653 17156
rect 29687 17153 29699 17187
rect 29641 17147 29699 17153
rect 29822 17144 29828 17196
rect 29880 17184 29886 17196
rect 30300 17193 30328 17224
rect 30834 17212 30840 17224
rect 30892 17212 30898 17264
rect 32320 17252 33120 17266
rect 32232 17224 33120 17252
rect 30285 17187 30343 17193
rect 30285 17184 30297 17187
rect 29880 17156 30297 17184
rect 29880 17144 29886 17156
rect 30285 17153 30297 17156
rect 30331 17153 30343 17187
rect 30285 17147 30343 17153
rect 30561 17187 30619 17193
rect 30561 17153 30573 17187
rect 30607 17153 30619 17187
rect 30561 17147 30619 17153
rect 20956 17088 22048 17116
rect 23569 17119 23627 17125
rect 20956 17076 20962 17088
rect 23569 17085 23581 17119
rect 23615 17085 23627 17119
rect 24946 17116 24952 17128
rect 24907 17088 24952 17116
rect 23569 17079 23627 17085
rect 20162 17008 20168 17060
rect 20220 17048 20226 17060
rect 22922 17048 22928 17060
rect 20220 17020 22928 17048
rect 20220 17008 20226 17020
rect 22922 17008 22928 17020
rect 22980 17048 22986 17060
rect 23198 17048 23204 17060
rect 22980 17020 23204 17048
rect 22980 17008 22986 17020
rect 23198 17008 23204 17020
rect 23256 17008 23262 17060
rect 23584 17048 23612 17079
rect 24946 17076 24952 17088
rect 25004 17076 25010 17128
rect 30006 17076 30012 17128
rect 30064 17116 30070 17128
rect 30466 17116 30472 17128
rect 30064 17088 30472 17116
rect 30064 17076 30070 17088
rect 30466 17076 30472 17088
rect 30524 17116 30530 17128
rect 30576 17116 30604 17147
rect 30650 17144 30656 17196
rect 30708 17184 30714 17196
rect 30745 17187 30803 17193
rect 30745 17184 30757 17187
rect 30708 17156 30757 17184
rect 30708 17144 30714 17156
rect 30745 17153 30757 17156
rect 30791 17184 30803 17187
rect 31018 17184 31024 17196
rect 30791 17156 31024 17184
rect 30791 17153 30803 17156
rect 30745 17147 30803 17153
rect 31018 17144 31024 17156
rect 31076 17144 31082 17196
rect 30524 17088 30604 17116
rect 32232 17116 32260 17224
rect 32320 17210 33120 17224
rect 32232 17088 32352 17116
rect 30524 17076 30530 17088
rect 23584 17020 24992 17048
rect 22094 16980 22100 16992
rect 18984 16952 22100 16980
rect 22094 16940 22100 16952
rect 22152 16940 22158 16992
rect 23382 16940 23388 16992
rect 23440 16980 23446 16992
rect 23477 16983 23535 16989
rect 23477 16980 23489 16983
rect 23440 16952 23489 16980
rect 23440 16940 23446 16952
rect 23477 16949 23489 16952
rect 23523 16949 23535 16983
rect 23477 16943 23535 16949
rect 23750 16940 23756 16992
rect 23808 16980 23814 16992
rect 24397 16983 24455 16989
rect 24397 16980 24409 16983
rect 23808 16952 24409 16980
rect 23808 16940 23814 16952
rect 24397 16949 24409 16952
rect 24443 16949 24455 16983
rect 24397 16943 24455 16949
rect 24486 16940 24492 16992
rect 24544 16980 24550 16992
rect 24762 16980 24768 16992
rect 24544 16952 24768 16980
rect 24544 16940 24550 16952
rect 24762 16940 24768 16952
rect 24820 16940 24826 16992
rect 24964 16980 24992 17020
rect 25222 16980 25228 16992
rect 24964 16952 25228 16980
rect 25222 16940 25228 16952
rect 25280 16980 25286 16992
rect 26050 16980 26056 16992
rect 25280 16952 26056 16980
rect 25280 16940 25286 16952
rect 26050 16940 26056 16952
rect 26108 16980 26114 16992
rect 26329 16983 26387 16989
rect 26329 16980 26341 16983
rect 26108 16952 26341 16980
rect 26108 16940 26114 16952
rect 26329 16949 26341 16952
rect 26375 16949 26387 16983
rect 26329 16943 26387 16949
rect 28997 16983 29055 16989
rect 28997 16949 29009 16983
rect 29043 16980 29055 16983
rect 29178 16980 29184 16992
rect 29043 16952 29184 16980
rect 29043 16949 29055 16952
rect 28997 16943 29055 16949
rect 29178 16940 29184 16952
rect 29236 16940 29242 16992
rect 29454 16980 29460 16992
rect 29415 16952 29460 16980
rect 29454 16940 29460 16952
rect 29512 16940 29518 16992
rect 30101 16983 30159 16989
rect 30101 16949 30113 16983
rect 30147 16980 30159 16983
rect 30834 16980 30840 16992
rect 30147 16952 30840 16980
rect 30147 16949 30159 16952
rect 30101 16943 30159 16949
rect 30834 16940 30840 16952
rect 30892 16940 30898 16992
rect 1104 16890 32016 16912
rect 1104 16838 2136 16890
rect 2188 16838 12440 16890
rect 12492 16838 22744 16890
rect 22796 16838 32016 16890
rect 1104 16816 32016 16838
rect 6914 16736 6920 16788
rect 6972 16776 6978 16788
rect 7929 16779 7987 16785
rect 7929 16776 7941 16779
rect 6972 16748 7941 16776
rect 6972 16736 6978 16748
rect 7929 16745 7941 16748
rect 7975 16745 7987 16779
rect 7929 16739 7987 16745
rect 8297 16779 8355 16785
rect 8297 16745 8309 16779
rect 8343 16776 8355 16779
rect 8846 16776 8852 16788
rect 8343 16748 8852 16776
rect 8343 16745 8355 16748
rect 8297 16739 8355 16745
rect 8846 16736 8852 16748
rect 8904 16736 8910 16788
rect 9416 16748 11284 16776
rect 6089 16711 6147 16717
rect 6089 16677 6101 16711
rect 6135 16708 6147 16711
rect 6135 16680 8892 16708
rect 6135 16677 6147 16680
rect 6089 16671 6147 16677
rect 2590 16600 2596 16652
rect 2648 16600 2654 16652
rect 3786 16640 3792 16652
rect 3747 16612 3792 16640
rect 3786 16600 3792 16612
rect 3844 16600 3850 16652
rect 5258 16600 5264 16652
rect 5316 16600 5322 16652
rect 6917 16643 6975 16649
rect 6917 16609 6929 16643
rect 6963 16640 6975 16643
rect 7834 16640 7840 16652
rect 6963 16612 7840 16640
rect 6963 16609 6975 16612
rect 6917 16603 6975 16609
rect 7834 16600 7840 16612
rect 7892 16600 7898 16652
rect 8386 16640 8392 16652
rect 8347 16612 8392 16640
rect 8386 16600 8392 16612
rect 8444 16600 8450 16652
rect 2038 16532 2044 16584
rect 2096 16572 2102 16584
rect 2133 16575 2191 16581
rect 2133 16572 2145 16575
rect 2096 16544 2145 16572
rect 2096 16532 2102 16544
rect 2133 16541 2145 16544
rect 2179 16541 2191 16575
rect 2133 16535 2191 16541
rect 2225 16575 2283 16581
rect 2225 16541 2237 16575
rect 2271 16572 2283 16575
rect 2774 16572 2780 16584
rect 2271 16544 2780 16572
rect 2271 16541 2283 16544
rect 2225 16535 2283 16541
rect 2774 16532 2780 16544
rect 2832 16532 2838 16584
rect 3973 16575 4031 16581
rect 3973 16541 3985 16575
rect 4019 16572 4031 16575
rect 4246 16572 4252 16584
rect 4019 16544 4252 16572
rect 4019 16541 4031 16544
rect 3973 16535 4031 16541
rect 4246 16532 4252 16544
rect 4304 16532 4310 16584
rect 5077 16575 5135 16581
rect 5077 16541 5089 16575
rect 5123 16572 5135 16575
rect 5442 16572 5448 16584
rect 5123 16544 5448 16572
rect 5123 16541 5135 16544
rect 5077 16535 5135 16541
rect 5442 16532 5448 16544
rect 5500 16532 5506 16584
rect 6546 16532 6552 16584
rect 6604 16572 6610 16584
rect 7101 16575 7159 16581
rect 7101 16572 7113 16575
rect 6604 16544 7113 16572
rect 6604 16532 6610 16544
rect 7101 16541 7113 16544
rect 7147 16541 7159 16575
rect 7101 16535 7159 16541
rect 7190 16532 7196 16584
rect 7248 16572 7254 16584
rect 7374 16572 7380 16584
rect 7248 16544 7293 16572
rect 7335 16544 7380 16572
rect 7248 16532 7254 16544
rect 7374 16532 7380 16544
rect 7432 16532 7438 16584
rect 7469 16575 7527 16581
rect 7469 16541 7481 16575
rect 7515 16572 7527 16575
rect 7558 16572 7564 16584
rect 7515 16544 7564 16572
rect 7515 16541 7527 16544
rect 7469 16535 7527 16541
rect 7558 16532 7564 16544
rect 7616 16532 7622 16584
rect 8113 16575 8171 16581
rect 8113 16541 8125 16575
rect 8159 16572 8171 16575
rect 8570 16572 8576 16584
rect 8159 16544 8576 16572
rect 8159 16541 8171 16544
rect 8113 16535 8171 16541
rect 8570 16532 8576 16544
rect 8628 16532 8634 16584
rect 8864 16572 8892 16680
rect 8938 16600 8944 16652
rect 8996 16640 9002 16652
rect 9416 16649 9444 16748
rect 11256 16649 11284 16748
rect 11422 16736 11428 16788
rect 11480 16776 11486 16788
rect 11974 16776 11980 16788
rect 11480 16748 11980 16776
rect 11480 16736 11486 16748
rect 11974 16736 11980 16748
rect 12032 16736 12038 16788
rect 12158 16736 12164 16788
rect 12216 16776 12222 16788
rect 12618 16776 12624 16788
rect 12216 16748 12624 16776
rect 12216 16736 12222 16748
rect 12618 16736 12624 16748
rect 12676 16736 12682 16788
rect 22097 16779 22155 16785
rect 12811 16748 16068 16776
rect 12250 16668 12256 16720
rect 12308 16708 12314 16720
rect 12811 16708 12839 16748
rect 12308 16680 12839 16708
rect 16040 16708 16068 16748
rect 16776 16748 21128 16776
rect 16776 16708 16804 16748
rect 16040 16680 16804 16708
rect 12308 16668 12314 16680
rect 17310 16668 17316 16720
rect 17368 16708 17374 16720
rect 17497 16711 17555 16717
rect 17497 16708 17509 16711
rect 17368 16680 17509 16708
rect 17368 16668 17374 16680
rect 17497 16677 17509 16680
rect 17543 16677 17555 16711
rect 20990 16708 20996 16720
rect 17497 16671 17555 16677
rect 17696 16680 18092 16708
rect 9401 16643 9459 16649
rect 9401 16640 9413 16643
rect 8996 16612 9413 16640
rect 8996 16600 9002 16612
rect 9401 16609 9413 16612
rect 9447 16609 9459 16643
rect 9401 16603 9459 16609
rect 11241 16643 11299 16649
rect 11241 16609 11253 16643
rect 11287 16609 11299 16643
rect 11241 16603 11299 16609
rect 13814 16600 13820 16652
rect 13872 16640 13878 16652
rect 14093 16643 14151 16649
rect 14093 16640 14105 16643
rect 13872 16612 14105 16640
rect 13872 16600 13878 16612
rect 14093 16609 14105 16612
rect 14139 16609 14151 16643
rect 14093 16603 14151 16609
rect 15102 16600 15108 16652
rect 15160 16640 15166 16652
rect 15286 16640 15292 16652
rect 15160 16612 15292 16640
rect 15160 16600 15166 16612
rect 15286 16600 15292 16612
rect 15344 16600 15350 16652
rect 15378 16600 15384 16652
rect 15436 16640 15442 16652
rect 16758 16640 16764 16652
rect 15436 16612 16068 16640
rect 16719 16612 16764 16640
rect 15436 16600 15442 16612
rect 10502 16572 10508 16584
rect 8864 16544 10508 16572
rect 10502 16532 10508 16544
rect 10560 16532 10566 16584
rect 11054 16532 11060 16584
rect 11112 16572 11118 16584
rect 11508 16575 11566 16581
rect 11508 16572 11520 16575
rect 11112 16544 11520 16572
rect 11112 16532 11118 16544
rect 11508 16541 11520 16544
rect 11554 16541 11566 16575
rect 11508 16535 11566 16541
rect 11974 16532 11980 16584
rect 12032 16572 12038 16584
rect 14360 16575 14418 16581
rect 12032 16544 13400 16572
rect 12032 16532 12038 16544
rect 2590 16504 2596 16516
rect 2551 16476 2596 16504
rect 2590 16464 2596 16476
rect 2648 16464 2654 16516
rect 2961 16507 3019 16513
rect 2961 16473 2973 16507
rect 3007 16504 3019 16507
rect 4157 16507 4215 16513
rect 4157 16504 4169 16507
rect 3007 16476 4169 16504
rect 3007 16473 3019 16476
rect 2961 16467 3019 16473
rect 4157 16473 4169 16476
rect 4203 16473 4215 16507
rect 4157 16467 4215 16473
rect 5169 16507 5227 16513
rect 5169 16473 5181 16507
rect 5215 16473 5227 16507
rect 5534 16504 5540 16516
rect 5495 16476 5540 16504
rect 5169 16467 5227 16473
rect 1486 16396 1492 16448
rect 1544 16436 1550 16448
rect 1857 16439 1915 16445
rect 1857 16436 1869 16439
rect 1544 16408 1869 16436
rect 1544 16396 1550 16408
rect 1857 16405 1869 16408
rect 1903 16405 1915 16439
rect 1857 16399 1915 16405
rect 2038 16396 2044 16448
rect 2096 16436 2102 16448
rect 2406 16436 2412 16448
rect 2096 16408 2412 16436
rect 2096 16396 2102 16408
rect 2406 16396 2412 16408
rect 2464 16396 2470 16448
rect 3142 16436 3148 16448
rect 3103 16408 3148 16436
rect 3142 16396 3148 16408
rect 3200 16396 3206 16448
rect 4798 16436 4804 16448
rect 4759 16408 4804 16436
rect 4798 16396 4804 16408
rect 4856 16396 4862 16448
rect 5184 16436 5212 16467
rect 5534 16464 5540 16476
rect 5592 16464 5598 16516
rect 5905 16507 5963 16513
rect 5905 16473 5917 16507
rect 5951 16504 5963 16507
rect 8202 16504 8208 16516
rect 5951 16476 8208 16504
rect 5951 16473 5963 16476
rect 5905 16467 5963 16473
rect 8202 16464 8208 16476
rect 8260 16464 8266 16516
rect 9214 16464 9220 16516
rect 9272 16504 9278 16516
rect 9646 16507 9704 16513
rect 9646 16504 9658 16507
rect 9272 16476 9658 16504
rect 9272 16464 9278 16476
rect 9646 16473 9658 16476
rect 9692 16473 9704 16507
rect 9646 16467 9704 16473
rect 10962 16464 10968 16516
rect 11020 16504 11026 16516
rect 12802 16504 12808 16516
rect 11020 16476 12808 16504
rect 11020 16464 11026 16476
rect 12802 16464 12808 16476
rect 12860 16464 12866 16516
rect 13170 16464 13176 16516
rect 13228 16504 13234 16516
rect 13265 16507 13323 16513
rect 13265 16504 13277 16507
rect 13228 16476 13277 16504
rect 13228 16464 13234 16476
rect 13265 16473 13277 16476
rect 13311 16473 13323 16507
rect 13372 16504 13400 16544
rect 14360 16541 14372 16575
rect 14406 16572 14418 16575
rect 15470 16572 15476 16584
rect 14406 16544 15476 16572
rect 14406 16541 14418 16544
rect 14360 16535 14418 16541
rect 15470 16532 15476 16544
rect 15528 16532 15534 16584
rect 15102 16504 15108 16516
rect 13372 16476 15108 16504
rect 13265 16467 13323 16473
rect 15102 16464 15108 16476
rect 15160 16464 15166 16516
rect 16040 16504 16068 16612
rect 16758 16600 16764 16612
rect 16816 16600 16822 16652
rect 17402 16600 17408 16652
rect 17460 16640 17466 16652
rect 17696 16640 17724 16680
rect 17460 16612 17724 16640
rect 18064 16640 18092 16680
rect 19812 16680 20996 16708
rect 18874 16640 18880 16652
rect 18064 16612 18880 16640
rect 17460 16600 17466 16612
rect 18248 16584 18276 16612
rect 18874 16600 18880 16612
rect 18932 16600 18938 16652
rect 19150 16600 19156 16652
rect 19208 16640 19214 16652
rect 19812 16649 19840 16680
rect 20990 16668 20996 16680
rect 21048 16668 21054 16720
rect 21100 16708 21128 16748
rect 22097 16745 22109 16779
rect 22143 16776 22155 16779
rect 22370 16776 22376 16788
rect 22143 16748 22376 16776
rect 22143 16745 22155 16748
rect 22097 16739 22155 16745
rect 22370 16736 22376 16748
rect 22428 16736 22434 16788
rect 22922 16736 22928 16788
rect 22980 16776 22986 16788
rect 23382 16776 23388 16788
rect 22980 16748 23388 16776
rect 22980 16736 22986 16748
rect 23382 16736 23388 16748
rect 23440 16736 23446 16788
rect 24026 16736 24032 16788
rect 24084 16776 24090 16788
rect 24210 16776 24216 16788
rect 24084 16748 24216 16776
rect 24084 16736 24090 16748
rect 24210 16736 24216 16748
rect 24268 16736 24274 16788
rect 24394 16776 24400 16788
rect 24355 16748 24400 16776
rect 24394 16736 24400 16748
rect 24452 16736 24458 16788
rect 24670 16736 24676 16788
rect 24728 16776 24734 16788
rect 25961 16779 26019 16785
rect 25961 16776 25973 16779
rect 24728 16748 25973 16776
rect 24728 16736 24734 16748
rect 25961 16745 25973 16748
rect 26007 16745 26019 16779
rect 25961 16739 26019 16745
rect 26050 16736 26056 16788
rect 26108 16776 26114 16788
rect 26697 16779 26755 16785
rect 26697 16776 26709 16779
rect 26108 16748 26709 16776
rect 26108 16736 26114 16748
rect 26697 16745 26709 16748
rect 26743 16745 26755 16779
rect 26697 16739 26755 16745
rect 26804 16748 31754 16776
rect 26804 16708 26832 16748
rect 21100 16680 26832 16708
rect 29914 16668 29920 16720
rect 29972 16708 29978 16720
rect 30837 16711 30895 16717
rect 30837 16708 30849 16711
rect 29972 16680 30849 16708
rect 29972 16668 29978 16680
rect 30837 16677 30849 16680
rect 30883 16677 30895 16711
rect 31726 16708 31754 16748
rect 32324 16708 32352 17088
rect 31726 16680 32352 16708
rect 30837 16671 30895 16677
rect 19337 16643 19395 16649
rect 19337 16640 19349 16643
rect 19208 16612 19349 16640
rect 19208 16600 19214 16612
rect 19337 16609 19349 16612
rect 19383 16609 19395 16643
rect 19337 16603 19395 16609
rect 19797 16643 19855 16649
rect 19797 16609 19809 16643
rect 19843 16609 19855 16643
rect 19797 16603 19855 16609
rect 20809 16643 20867 16649
rect 20809 16609 20821 16643
rect 20855 16640 20867 16643
rect 20898 16640 20904 16652
rect 20855 16612 20904 16640
rect 20855 16609 20867 16612
rect 20809 16603 20867 16609
rect 20898 16600 20904 16612
rect 20956 16600 20962 16652
rect 21008 16640 21036 16668
rect 25038 16640 25044 16652
rect 21008 16612 21588 16640
rect 16117 16575 16175 16581
rect 16117 16541 16129 16575
rect 16163 16572 16175 16575
rect 16298 16572 16304 16584
rect 16163 16544 16304 16572
rect 16163 16541 16175 16544
rect 16117 16535 16175 16541
rect 16298 16532 16304 16544
rect 16356 16572 16362 16584
rect 16577 16575 16635 16581
rect 16577 16572 16589 16575
rect 16356 16544 16589 16572
rect 16356 16532 16362 16544
rect 16577 16541 16589 16544
rect 16623 16541 16635 16575
rect 16577 16535 16635 16541
rect 16669 16575 16727 16581
rect 16669 16541 16681 16575
rect 16715 16572 16727 16575
rect 17034 16572 17040 16584
rect 16715 16544 17040 16572
rect 16715 16541 16727 16544
rect 16669 16535 16727 16541
rect 17034 16532 17040 16544
rect 17092 16532 17098 16584
rect 17770 16572 17776 16584
rect 17731 16544 17776 16572
rect 17770 16532 17776 16544
rect 17828 16532 17834 16584
rect 18049 16575 18107 16581
rect 18049 16572 18061 16575
rect 17926 16544 18061 16572
rect 17926 16504 17954 16544
rect 18049 16541 18061 16544
rect 18095 16541 18107 16575
rect 18049 16535 18107 16541
rect 18230 16532 18236 16584
rect 18288 16532 18294 16584
rect 19518 16572 19524 16584
rect 19479 16544 19524 16572
rect 19518 16532 19524 16544
rect 19576 16532 19582 16584
rect 21560 16581 21588 16612
rect 22848 16612 25044 16640
rect 19705 16575 19763 16581
rect 19705 16541 19717 16575
rect 19751 16541 19763 16575
rect 20993 16575 21051 16581
rect 20993 16572 21005 16575
rect 19705 16535 19763 16541
rect 19904 16544 21005 16572
rect 15304 16476 15976 16504
rect 16040 16476 17954 16504
rect 19720 16504 19748 16535
rect 19794 16504 19800 16516
rect 19720 16476 19800 16504
rect 5718 16436 5724 16448
rect 5184 16408 5724 16436
rect 5718 16396 5724 16408
rect 5776 16396 5782 16448
rect 6730 16396 6736 16448
rect 6788 16436 6794 16448
rect 9490 16436 9496 16448
rect 6788 16408 9496 16436
rect 6788 16396 6794 16408
rect 9490 16396 9496 16408
rect 9548 16396 9554 16448
rect 9766 16396 9772 16448
rect 9824 16436 9830 16448
rect 10594 16436 10600 16448
rect 9824 16408 10600 16436
rect 9824 16396 9830 16408
rect 10594 16396 10600 16408
rect 10652 16436 10658 16448
rect 10778 16436 10784 16448
rect 10652 16408 10784 16436
rect 10652 16396 10658 16408
rect 10778 16396 10784 16408
rect 10836 16396 10842 16448
rect 11422 16396 11428 16448
rect 11480 16436 11486 16448
rect 12158 16436 12164 16448
rect 11480 16408 12164 16436
rect 11480 16396 11486 16408
rect 12158 16396 12164 16408
rect 12216 16396 12222 16448
rect 12250 16396 12256 16448
rect 12308 16436 12314 16448
rect 13357 16439 13415 16445
rect 13357 16436 13369 16439
rect 12308 16408 13369 16436
rect 12308 16396 12314 16408
rect 13357 16405 13369 16408
rect 13403 16405 13415 16439
rect 13357 16399 13415 16405
rect 14826 16396 14832 16448
rect 14884 16436 14890 16448
rect 15304 16436 15332 16476
rect 14884 16408 15332 16436
rect 14884 16396 14890 16408
rect 15378 16396 15384 16448
rect 15436 16436 15442 16448
rect 15473 16439 15531 16445
rect 15473 16436 15485 16439
rect 15436 16408 15485 16436
rect 15436 16396 15442 16408
rect 15473 16405 15485 16408
rect 15519 16405 15531 16439
rect 15473 16399 15531 16405
rect 15562 16396 15568 16448
rect 15620 16436 15626 16448
rect 15838 16436 15844 16448
rect 15620 16408 15844 16436
rect 15620 16396 15626 16408
rect 15838 16396 15844 16408
rect 15896 16396 15902 16448
rect 15948 16436 15976 16476
rect 19794 16464 19800 16476
rect 19852 16464 19858 16516
rect 16117 16439 16175 16445
rect 16117 16436 16129 16439
rect 15948 16408 16129 16436
rect 16117 16405 16129 16408
rect 16163 16405 16175 16439
rect 16117 16399 16175 16405
rect 16209 16439 16267 16445
rect 16209 16405 16221 16439
rect 16255 16436 16267 16439
rect 17957 16439 18015 16445
rect 17957 16436 17969 16439
rect 16255 16408 17969 16436
rect 16255 16405 16267 16408
rect 16209 16399 16267 16405
rect 17957 16405 17969 16408
rect 18003 16405 18015 16439
rect 17957 16399 18015 16405
rect 18598 16396 18604 16448
rect 18656 16436 18662 16448
rect 19904 16436 19932 16544
rect 20993 16541 21005 16544
rect 21039 16541 21051 16575
rect 20993 16535 21051 16541
rect 21269 16575 21327 16581
rect 21269 16541 21281 16575
rect 21315 16572 21327 16575
rect 21545 16575 21603 16581
rect 21315 16544 21496 16572
rect 21315 16541 21327 16544
rect 21269 16535 21327 16541
rect 21008 16504 21036 16535
rect 21468 16504 21496 16544
rect 21545 16541 21557 16575
rect 21591 16541 21603 16575
rect 21545 16535 21603 16541
rect 22278 16532 22284 16584
rect 22336 16532 22342 16584
rect 22370 16532 22376 16584
rect 22428 16572 22434 16584
rect 22848 16581 22876 16612
rect 25038 16600 25044 16612
rect 25096 16640 25102 16652
rect 25096 16612 25176 16640
rect 25096 16600 25102 16612
rect 22557 16575 22615 16581
rect 22557 16572 22569 16575
rect 22428 16544 22569 16572
rect 22428 16532 22434 16544
rect 22557 16541 22569 16544
rect 22603 16541 22615 16575
rect 22557 16535 22615 16541
rect 22833 16575 22891 16581
rect 22833 16541 22845 16575
rect 22879 16541 22891 16575
rect 22833 16535 22891 16541
rect 23017 16575 23075 16581
rect 23017 16541 23029 16575
rect 23063 16572 23075 16575
rect 23106 16572 23112 16584
rect 23063 16544 23112 16572
rect 23063 16541 23075 16544
rect 23017 16535 23075 16541
rect 22296 16504 22324 16532
rect 22848 16504 22876 16535
rect 23106 16532 23112 16544
rect 23164 16532 23170 16584
rect 23569 16575 23627 16581
rect 23569 16541 23581 16575
rect 23615 16572 23627 16575
rect 24302 16572 24308 16584
rect 23615 16544 24308 16572
rect 23615 16541 23627 16544
rect 23569 16535 23627 16541
rect 24302 16532 24308 16544
rect 24360 16572 24366 16584
rect 24486 16572 24492 16584
rect 24360 16544 24492 16572
rect 24360 16532 24366 16544
rect 24486 16532 24492 16544
rect 24544 16532 24550 16584
rect 24578 16532 24584 16584
rect 24636 16572 24642 16584
rect 25148 16581 25176 16612
rect 26142 16600 26148 16652
rect 26200 16640 26206 16652
rect 26200 16612 29592 16640
rect 26200 16600 26206 16612
rect 24857 16575 24915 16581
rect 24857 16572 24869 16575
rect 24636 16544 24869 16572
rect 24636 16532 24642 16544
rect 24857 16541 24869 16544
rect 24903 16541 24915 16575
rect 24857 16535 24915 16541
rect 25133 16575 25191 16581
rect 25133 16541 25145 16575
rect 25179 16541 25191 16575
rect 25133 16535 25191 16541
rect 25222 16532 25228 16584
rect 25280 16572 25286 16584
rect 25317 16575 25375 16581
rect 25317 16572 25329 16575
rect 25280 16544 25329 16572
rect 25280 16532 25286 16544
rect 25317 16541 25329 16544
rect 25363 16541 25375 16575
rect 25317 16535 25375 16541
rect 25774 16532 25780 16584
rect 25832 16572 25838 16584
rect 26605 16575 26663 16581
rect 26605 16572 26617 16575
rect 25832 16544 26617 16572
rect 25832 16532 25838 16544
rect 26605 16541 26617 16544
rect 26651 16572 26663 16575
rect 26694 16572 26700 16584
rect 26651 16544 26700 16572
rect 26651 16541 26663 16544
rect 26605 16535 26663 16541
rect 26694 16532 26700 16544
rect 26752 16532 26758 16584
rect 26786 16532 26792 16584
rect 26844 16572 26850 16584
rect 26881 16575 26939 16581
rect 26881 16572 26893 16575
rect 26844 16544 26893 16572
rect 26844 16532 26850 16544
rect 26881 16541 26893 16544
rect 26927 16541 26939 16575
rect 26881 16535 26939 16541
rect 27246 16532 27252 16584
rect 27304 16572 27310 16584
rect 27709 16575 27767 16581
rect 27709 16572 27721 16575
rect 27304 16544 27721 16572
rect 27304 16532 27310 16544
rect 27709 16541 27721 16544
rect 27755 16541 27767 16575
rect 27709 16535 27767 16541
rect 28261 16575 28319 16581
rect 28261 16541 28273 16575
rect 28307 16572 28319 16575
rect 28350 16572 28356 16584
rect 28307 16544 28356 16572
rect 28307 16541 28319 16544
rect 28261 16535 28319 16541
rect 28350 16532 28356 16544
rect 28408 16532 28414 16584
rect 29564 16581 29592 16612
rect 29549 16575 29607 16581
rect 29549 16541 29561 16575
rect 29595 16541 29607 16575
rect 29549 16535 29607 16541
rect 21008 16476 21312 16504
rect 21468 16476 22324 16504
rect 22572 16476 22876 16504
rect 18656 16408 19932 16436
rect 18656 16396 18662 16408
rect 20070 16396 20076 16448
rect 20128 16436 20134 16448
rect 21177 16439 21235 16445
rect 21177 16436 21189 16439
rect 20128 16408 21189 16436
rect 20128 16396 20134 16408
rect 21177 16405 21189 16408
rect 21223 16405 21235 16439
rect 21284 16436 21312 16476
rect 22572 16448 22600 16476
rect 23474 16464 23480 16516
rect 23532 16504 23538 16516
rect 25869 16507 25927 16513
rect 25869 16504 25881 16507
rect 23532 16476 25881 16504
rect 23532 16464 23538 16476
rect 25869 16473 25881 16476
rect 25915 16473 25927 16507
rect 25869 16467 25927 16473
rect 28445 16507 28503 16513
rect 28445 16473 28457 16507
rect 28491 16504 28503 16507
rect 28534 16504 28540 16516
rect 28491 16476 28540 16504
rect 28491 16473 28503 16476
rect 28445 16467 28503 16473
rect 28534 16464 28540 16476
rect 28592 16504 28598 16516
rect 31386 16504 31392 16516
rect 28592 16476 31392 16504
rect 28592 16464 28598 16476
rect 31386 16464 31392 16476
rect 31444 16464 31450 16516
rect 21637 16439 21695 16445
rect 21637 16436 21649 16439
rect 21284 16408 21649 16436
rect 21177 16399 21235 16405
rect 21637 16405 21649 16408
rect 21683 16405 21695 16439
rect 21637 16399 21695 16405
rect 22278 16396 22284 16448
rect 22336 16436 22342 16448
rect 22373 16439 22431 16445
rect 22373 16436 22385 16439
rect 22336 16408 22385 16436
rect 22336 16396 22342 16408
rect 22373 16405 22385 16408
rect 22419 16405 22431 16439
rect 22373 16399 22431 16405
rect 22554 16396 22560 16448
rect 22612 16396 22618 16448
rect 23753 16439 23811 16445
rect 23753 16405 23765 16439
rect 23799 16436 23811 16439
rect 23937 16439 23995 16445
rect 23937 16436 23949 16439
rect 23799 16408 23949 16436
rect 23799 16405 23811 16408
rect 23753 16399 23811 16405
rect 23937 16405 23949 16408
rect 23983 16405 23995 16439
rect 23937 16399 23995 16405
rect 24026 16396 24032 16448
rect 24084 16436 24090 16448
rect 24673 16439 24731 16445
rect 24673 16436 24685 16439
rect 24084 16408 24685 16436
rect 24084 16396 24090 16408
rect 24673 16405 24685 16408
rect 24719 16405 24731 16439
rect 24673 16399 24731 16405
rect 26050 16396 26056 16448
rect 26108 16436 26114 16448
rect 27157 16439 27215 16445
rect 27157 16436 27169 16439
rect 26108 16408 27169 16436
rect 26108 16396 26114 16408
rect 27157 16405 27169 16408
rect 27203 16405 27215 16439
rect 27157 16399 27215 16405
rect 1104 16346 32016 16368
rect 1104 16294 7288 16346
rect 7340 16294 17592 16346
rect 17644 16294 27896 16346
rect 27948 16294 32016 16346
rect 1104 16272 32016 16294
rect 5077 16235 5135 16241
rect 5077 16201 5089 16235
rect 5123 16232 5135 16235
rect 5534 16232 5540 16244
rect 5123 16204 5540 16232
rect 5123 16201 5135 16204
rect 5077 16195 5135 16201
rect 5534 16192 5540 16204
rect 5592 16192 5598 16244
rect 5905 16235 5963 16241
rect 5905 16201 5917 16235
rect 5951 16232 5963 16235
rect 6362 16232 6368 16244
rect 5951 16204 6368 16232
rect 5951 16201 5963 16204
rect 5905 16195 5963 16201
rect 6362 16192 6368 16204
rect 6420 16232 6426 16244
rect 7285 16235 7343 16241
rect 7285 16232 7297 16235
rect 6420 16204 7297 16232
rect 6420 16192 6426 16204
rect 7285 16201 7297 16204
rect 7331 16201 7343 16235
rect 7285 16195 7343 16201
rect 7374 16192 7380 16244
rect 7432 16232 7438 16244
rect 7469 16235 7527 16241
rect 7469 16232 7481 16235
rect 7432 16204 7481 16232
rect 7432 16192 7438 16204
rect 7469 16201 7481 16204
rect 7515 16201 7527 16235
rect 7469 16195 7527 16201
rect 8202 16192 8208 16244
rect 8260 16232 8266 16244
rect 8297 16235 8355 16241
rect 8297 16232 8309 16235
rect 8260 16204 8309 16232
rect 8260 16192 8266 16204
rect 8297 16201 8309 16204
rect 8343 16201 8355 16235
rect 9214 16232 9220 16244
rect 9175 16204 9220 16232
rect 8297 16195 8355 16201
rect 9214 16192 9220 16204
rect 9272 16192 9278 16244
rect 11790 16232 11796 16244
rect 11751 16204 11796 16232
rect 11790 16192 11796 16204
rect 11848 16192 11854 16244
rect 12342 16192 12348 16244
rect 12400 16232 12406 16244
rect 14366 16232 14372 16244
rect 12400 16204 14372 16232
rect 12400 16192 12406 16204
rect 14366 16192 14372 16204
rect 14424 16232 14430 16244
rect 18046 16232 18052 16244
rect 14424 16204 18052 16232
rect 14424 16192 14430 16204
rect 18046 16192 18052 16204
rect 18104 16192 18110 16244
rect 18417 16235 18475 16241
rect 18417 16232 18429 16235
rect 18156 16204 18429 16232
rect 2124 16167 2182 16173
rect 2124 16133 2136 16167
rect 2170 16164 2182 16167
rect 2222 16164 2228 16176
rect 2170 16136 2228 16164
rect 2170 16133 2182 16136
rect 2124 16127 2182 16133
rect 2222 16124 2228 16136
rect 2280 16124 2286 16176
rect 3142 16124 3148 16176
rect 3200 16164 3206 16176
rect 14826 16164 14832 16176
rect 3200 16136 14832 16164
rect 3200 16124 3206 16136
rect 14826 16124 14832 16136
rect 14884 16124 14890 16176
rect 15286 16124 15292 16176
rect 15344 16164 15350 16176
rect 15838 16164 15844 16176
rect 15344 16136 15844 16164
rect 15344 16124 15350 16136
rect 15838 16124 15844 16136
rect 15896 16124 15902 16176
rect 16117 16167 16175 16173
rect 16117 16133 16129 16167
rect 16163 16164 16175 16167
rect 16669 16167 16727 16173
rect 16163 16136 16611 16164
rect 16163 16133 16175 16136
rect 16117 16127 16175 16133
rect 3878 16056 3884 16108
rect 3936 16096 3942 16108
rect 4065 16099 4123 16105
rect 4065 16096 4077 16099
rect 3936 16068 4077 16096
rect 3936 16056 3942 16068
rect 4065 16065 4077 16068
rect 4111 16065 4123 16099
rect 4065 16059 4123 16065
rect 4430 16056 4436 16108
rect 4488 16096 4494 16108
rect 5445 16099 5503 16105
rect 5445 16096 5457 16099
rect 4488 16068 5457 16096
rect 4488 16056 4494 16068
rect 5445 16065 5457 16068
rect 5491 16065 5503 16099
rect 5445 16059 5503 16065
rect 5537 16099 5595 16105
rect 5537 16065 5549 16099
rect 5583 16096 5595 16099
rect 5905 16099 5963 16105
rect 5905 16096 5917 16099
rect 5583 16068 5917 16096
rect 5583 16065 5595 16068
rect 5537 16059 5595 16065
rect 5905 16065 5917 16068
rect 5951 16065 5963 16099
rect 5905 16059 5963 16065
rect 5994 16056 6000 16108
rect 6052 16096 6058 16108
rect 7558 16096 7564 16108
rect 6052 16068 7564 16096
rect 6052 16056 6058 16068
rect 7558 16056 7564 16068
rect 7616 16056 7622 16108
rect 7834 16056 7840 16108
rect 7892 16096 7898 16108
rect 8113 16099 8171 16105
rect 8113 16096 8125 16099
rect 7892 16068 8125 16096
rect 7892 16056 7898 16068
rect 8113 16065 8125 16068
rect 8159 16065 8171 16099
rect 8113 16059 8171 16065
rect 9401 16099 9459 16105
rect 9401 16065 9413 16099
rect 9447 16096 9459 16099
rect 10137 16099 10195 16105
rect 10137 16096 10149 16099
rect 9447 16068 10149 16096
rect 9447 16065 9459 16068
rect 9401 16059 9459 16065
rect 10137 16065 10149 16068
rect 10183 16065 10195 16099
rect 10318 16096 10324 16108
rect 10279 16068 10324 16096
rect 10137 16059 10195 16065
rect 10318 16056 10324 16068
rect 10376 16056 10382 16108
rect 10597 16099 10655 16105
rect 10597 16065 10609 16099
rect 10643 16065 10655 16099
rect 10778 16096 10784 16108
rect 10739 16068 10784 16096
rect 10597 16059 10655 16065
rect 1394 15988 1400 16040
rect 1452 16028 1458 16040
rect 1854 16028 1860 16040
rect 1452 16000 1860 16028
rect 1452 15988 1458 16000
rect 1854 15988 1860 16000
rect 1912 15988 1918 16040
rect 3789 16031 3847 16037
rect 3789 15997 3801 16031
rect 3835 15997 3847 16031
rect 3789 15991 3847 15997
rect 5629 16031 5687 16037
rect 5629 15997 5641 16031
rect 5675 15997 5687 16031
rect 5629 15991 5687 15997
rect 6917 16031 6975 16037
rect 6917 15997 6929 16031
rect 6963 15997 6975 16031
rect 6917 15991 6975 15997
rect 3237 15963 3295 15969
rect 3237 15929 3249 15963
rect 3283 15960 3295 15963
rect 3804 15960 3832 15991
rect 4338 15960 4344 15972
rect 3283 15932 4344 15960
rect 3283 15929 3295 15932
rect 3237 15923 3295 15929
rect 4338 15920 4344 15932
rect 4396 15920 4402 15972
rect 5074 15920 5080 15972
rect 5132 15960 5138 15972
rect 5644 15960 5672 15991
rect 5132 15932 5672 15960
rect 6932 15960 6960 15991
rect 7466 15988 7472 16040
rect 7524 16028 7530 16040
rect 7929 16031 7987 16037
rect 7929 16028 7941 16031
rect 7524 16000 7941 16028
rect 7524 15988 7530 16000
rect 7929 15997 7941 16000
rect 7975 15997 7987 16031
rect 9674 16028 9680 16040
rect 9635 16000 9680 16028
rect 7929 15991 7987 15997
rect 9674 15988 9680 16000
rect 9732 15988 9738 16040
rect 10612 16028 10640 16059
rect 10778 16056 10784 16068
rect 10836 16056 10842 16108
rect 11514 16056 11520 16108
rect 11572 16096 11578 16108
rect 11977 16099 12035 16105
rect 11977 16096 11989 16099
rect 11572 16068 11989 16096
rect 11572 16056 11578 16068
rect 11977 16065 11989 16068
rect 12023 16065 12035 16099
rect 11977 16059 12035 16065
rect 12253 16099 12311 16105
rect 12253 16065 12265 16099
rect 12299 16065 12311 16099
rect 12253 16059 12311 16065
rect 12437 16099 12495 16105
rect 12437 16065 12449 16099
rect 12483 16096 12495 16099
rect 12618 16096 12624 16108
rect 12483 16068 12624 16096
rect 12483 16065 12495 16068
rect 12437 16059 12495 16065
rect 12066 16028 12072 16040
rect 10612 16000 12072 16028
rect 12066 15988 12072 16000
rect 12124 16028 12130 16040
rect 12268 16028 12296 16059
rect 12618 16056 12624 16068
rect 12676 16056 12682 16108
rect 13541 16099 13599 16105
rect 13541 16096 13553 16099
rect 12728 16068 13553 16096
rect 12728 16028 12756 16068
rect 13541 16065 13553 16068
rect 13587 16065 13599 16099
rect 13541 16059 13599 16065
rect 13630 16056 13636 16108
rect 13688 16096 13694 16108
rect 13688 16068 14964 16096
rect 13688 16056 13694 16068
rect 12124 16000 12756 16028
rect 13265 16031 13323 16037
rect 12124 15988 12130 16000
rect 13265 15997 13277 16031
rect 13311 16028 13323 16031
rect 14366 16028 14372 16040
rect 13311 16000 14372 16028
rect 13311 15997 13323 16000
rect 13265 15991 13323 15997
rect 14366 15988 14372 16000
rect 14424 15988 14430 16040
rect 14936 16028 14964 16068
rect 15010 16056 15016 16108
rect 15068 16096 15074 16108
rect 15114 16099 15172 16105
rect 15114 16096 15126 16099
rect 15068 16068 15126 16096
rect 15068 16056 15074 16068
rect 15114 16065 15126 16068
rect 15160 16065 15172 16099
rect 15114 16059 15172 16065
rect 15381 16099 15439 16105
rect 15381 16065 15393 16099
rect 15427 16096 15439 16099
rect 15470 16096 15476 16108
rect 15427 16068 15476 16096
rect 15427 16065 15439 16068
rect 15381 16059 15439 16065
rect 15470 16056 15476 16068
rect 15528 16056 15534 16108
rect 15565 16099 15623 16105
rect 15565 16065 15577 16099
rect 15611 16096 15623 16099
rect 15654 16096 15660 16108
rect 15611 16068 15660 16096
rect 15611 16065 15623 16068
rect 15565 16059 15623 16065
rect 15654 16056 15660 16068
rect 15712 16096 15718 16108
rect 16583 16096 16611 16136
rect 16669 16133 16681 16167
rect 16715 16164 16727 16167
rect 17282 16167 17340 16173
rect 17282 16164 17294 16167
rect 16715 16136 17294 16164
rect 16715 16133 16727 16136
rect 16669 16127 16727 16133
rect 17282 16133 17294 16136
rect 17328 16133 17340 16167
rect 17282 16127 17340 16133
rect 18156 16096 18184 16204
rect 18417 16201 18429 16204
rect 18463 16201 18475 16235
rect 20254 16232 20260 16244
rect 20215 16204 20260 16232
rect 18417 16195 18475 16201
rect 20254 16192 20260 16204
rect 20312 16192 20318 16244
rect 21266 16192 21272 16244
rect 21324 16232 21330 16244
rect 23474 16232 23480 16244
rect 21324 16204 23480 16232
rect 21324 16192 21330 16204
rect 23474 16192 23480 16204
rect 23532 16192 23538 16244
rect 23658 16232 23664 16244
rect 23619 16204 23664 16232
rect 23658 16192 23664 16204
rect 23716 16192 23722 16244
rect 24394 16192 24400 16244
rect 24452 16232 24458 16244
rect 24949 16235 25007 16241
rect 24949 16232 24961 16235
rect 24452 16204 24961 16232
rect 24452 16192 24458 16204
rect 24949 16201 24961 16204
rect 24995 16201 25007 16235
rect 24949 16195 25007 16201
rect 25777 16235 25835 16241
rect 25777 16201 25789 16235
rect 25823 16232 25835 16235
rect 28258 16232 28264 16244
rect 25823 16204 28264 16232
rect 25823 16201 25835 16204
rect 25777 16195 25835 16201
rect 28258 16192 28264 16204
rect 28316 16192 28322 16244
rect 31205 16235 31263 16241
rect 29288 16204 31156 16232
rect 19150 16173 19156 16176
rect 19144 16164 19156 16173
rect 19111 16136 19156 16164
rect 19144 16127 19156 16136
rect 19150 16124 19156 16127
rect 19208 16124 19214 16176
rect 21085 16167 21143 16173
rect 21085 16164 21097 16167
rect 19260 16136 21097 16164
rect 18874 16096 18880 16108
rect 15712 16068 16528 16096
rect 16583 16068 18184 16096
rect 18835 16068 18880 16096
rect 15712 16056 15718 16068
rect 16117 16031 16175 16037
rect 16117 16028 16129 16031
rect 14936 16000 16129 16028
rect 16117 15997 16129 16000
rect 16163 15997 16175 16031
rect 16500 16028 16528 16068
rect 18874 16056 18880 16068
rect 18932 16056 18938 16108
rect 19260 16096 19288 16136
rect 21085 16133 21097 16136
rect 21131 16133 21143 16167
rect 21085 16127 21143 16133
rect 21450 16124 21456 16176
rect 21508 16164 21514 16176
rect 21508 16136 22315 16164
rect 21508 16124 21514 16136
rect 18984 16068 19288 16096
rect 17034 16028 17040 16040
rect 16500 16000 16804 16028
rect 16995 16000 17040 16028
rect 16117 15991 16175 15997
rect 7190 15960 7196 15972
rect 6932 15932 7196 15960
rect 5132 15920 5138 15932
rect 7190 15920 7196 15932
rect 7248 15920 7254 15972
rect 9585 15963 9643 15969
rect 9585 15929 9597 15963
rect 9631 15960 9643 15963
rect 10042 15960 10048 15972
rect 9631 15932 10048 15960
rect 9631 15929 9643 15932
rect 9585 15923 9643 15929
rect 10042 15920 10048 15932
rect 10100 15960 10106 15972
rect 12158 15960 12164 15972
rect 10100 15932 12164 15960
rect 10100 15920 10106 15932
rect 12158 15920 12164 15932
rect 12216 15920 12222 15972
rect 16669 15963 16727 15969
rect 16669 15960 16681 15963
rect 12728 15932 16681 15960
rect 937 15895 995 15901
rect 937 15861 949 15895
rect 983 15892 995 15895
rect 1854 15892 1860 15904
rect 983 15864 1860 15892
rect 983 15861 995 15864
rect 937 15855 995 15861
rect 1854 15852 1860 15864
rect 1912 15892 1918 15904
rect 6638 15892 6644 15904
rect 1912 15864 6644 15892
rect 1912 15852 1918 15864
rect 6638 15852 6644 15864
rect 6696 15852 6702 15904
rect 7285 15895 7343 15901
rect 7285 15861 7297 15895
rect 7331 15892 7343 15895
rect 7374 15892 7380 15904
rect 7331 15864 7380 15892
rect 7331 15861 7343 15864
rect 7285 15855 7343 15861
rect 7374 15852 7380 15864
rect 7432 15852 7438 15904
rect 9490 15852 9496 15904
rect 9548 15892 9554 15904
rect 12728 15892 12756 15932
rect 16669 15929 16681 15932
rect 16715 15929 16727 15963
rect 16776 15960 16804 16000
rect 17034 15988 17040 16000
rect 17092 15988 17098 16040
rect 18046 15988 18052 16040
rect 18104 16028 18110 16040
rect 18984 16028 19012 16068
rect 20254 16056 20260 16108
rect 20312 16096 20318 16108
rect 20717 16099 20775 16105
rect 20717 16096 20729 16099
rect 20312 16068 20729 16096
rect 20312 16056 20318 16068
rect 20717 16065 20729 16068
rect 20763 16065 20775 16099
rect 20717 16059 20775 16065
rect 21821 16099 21879 16105
rect 21821 16065 21833 16099
rect 21867 16096 21879 16099
rect 21910 16096 21916 16108
rect 21867 16068 21916 16096
rect 21867 16065 21879 16068
rect 21821 16059 21879 16065
rect 21910 16056 21916 16068
rect 21968 16056 21974 16108
rect 22094 16105 22100 16108
rect 22088 16059 22100 16105
rect 22152 16096 22158 16108
rect 22287 16096 22315 16136
rect 23198 16124 23204 16176
rect 23256 16164 23262 16176
rect 25222 16164 25228 16176
rect 23256 16136 25228 16164
rect 23256 16124 23262 16136
rect 25222 16124 25228 16136
rect 25280 16124 25286 16176
rect 26329 16167 26387 16173
rect 26329 16133 26341 16167
rect 26375 16164 26387 16167
rect 29288 16164 29316 16204
rect 26375 16136 29316 16164
rect 29365 16167 29423 16173
rect 26375 16133 26387 16136
rect 26329 16127 26387 16133
rect 29365 16133 29377 16167
rect 29411 16164 29423 16167
rect 30374 16164 30380 16176
rect 29411 16136 30380 16164
rect 29411 16133 29423 16136
rect 29365 16127 29423 16133
rect 30374 16124 30380 16136
rect 30432 16124 30438 16176
rect 31128 16164 31156 16204
rect 31205 16201 31217 16235
rect 31251 16232 31263 16235
rect 31294 16232 31300 16244
rect 31251 16204 31300 16232
rect 31251 16201 31263 16204
rect 31205 16195 31263 16201
rect 31294 16192 31300 16204
rect 31352 16192 31358 16244
rect 31478 16164 31484 16176
rect 31128 16136 31484 16164
rect 31478 16124 31484 16136
rect 31536 16124 31542 16176
rect 23566 16096 23572 16108
rect 22152 16068 22188 16096
rect 22287 16068 23572 16096
rect 22094 16056 22100 16059
rect 22152 16056 22158 16068
rect 23566 16056 23572 16068
rect 23624 16056 23630 16108
rect 23845 16099 23903 16105
rect 23845 16065 23857 16099
rect 23891 16096 23903 16099
rect 23934 16096 23940 16108
rect 23891 16068 23940 16096
rect 23891 16065 23903 16068
rect 23845 16059 23903 16065
rect 23934 16056 23940 16068
rect 23992 16056 23998 16108
rect 24394 16096 24400 16108
rect 24228 16068 24400 16096
rect 18104 16000 19012 16028
rect 18104 15988 18110 16000
rect 23382 15988 23388 16040
rect 23440 16028 23446 16040
rect 24228 16028 24256 16068
rect 24394 16056 24400 16068
rect 24452 16056 24458 16108
rect 24489 16099 24547 16105
rect 24489 16065 24501 16099
rect 24535 16096 24547 16099
rect 25958 16096 25964 16108
rect 24535 16068 25964 16096
rect 24535 16065 24547 16068
rect 24489 16059 24547 16065
rect 25958 16056 25964 16068
rect 26016 16056 26022 16108
rect 26050 16056 26056 16108
rect 26108 16096 26114 16108
rect 26108 16068 26153 16096
rect 26108 16056 26114 16068
rect 26970 16056 26976 16108
rect 27028 16096 27034 16108
rect 27065 16099 27123 16105
rect 27065 16096 27077 16099
rect 27028 16068 27077 16096
rect 27028 16056 27034 16068
rect 27065 16065 27077 16068
rect 27111 16065 27123 16099
rect 28261 16099 28319 16105
rect 27065 16059 27123 16065
rect 27264 16068 28212 16096
rect 27264 16040 27292 16068
rect 23440 16000 24256 16028
rect 24305 16031 24363 16037
rect 23440 15988 23446 16000
rect 24305 15997 24317 16031
rect 24351 16028 24363 16031
rect 24670 16028 24676 16040
rect 24351 16000 24676 16028
rect 24351 15997 24363 16000
rect 24305 15991 24363 15997
rect 24670 15988 24676 16000
rect 24728 15988 24734 16040
rect 24857 16031 24915 16037
rect 24857 15997 24869 16031
rect 24903 16028 24915 16031
rect 24949 16031 25007 16037
rect 24949 16028 24961 16031
rect 24903 16000 24961 16028
rect 24903 15997 24915 16000
rect 24857 15991 24915 15997
rect 24949 15997 24961 16000
rect 24995 15997 25007 16031
rect 24949 15991 25007 15997
rect 25777 16031 25835 16037
rect 25777 15997 25789 16031
rect 25823 16028 25835 16031
rect 25869 16031 25927 16037
rect 25869 16028 25881 16031
rect 25823 16000 25881 16028
rect 25823 15997 25835 16000
rect 25777 15991 25835 15997
rect 25869 15997 25881 16000
rect 25915 15997 25927 16031
rect 25869 15991 25927 15997
rect 26421 16031 26479 16037
rect 26421 15997 26433 16031
rect 26467 16028 26479 16031
rect 27246 16028 27252 16040
rect 26467 16000 27252 16028
rect 26467 15997 26479 16000
rect 26421 15991 26479 15997
rect 16942 15960 16948 15972
rect 16776 15932 16948 15960
rect 16669 15923 16727 15929
rect 16942 15920 16948 15932
rect 17000 15920 17006 15972
rect 24394 15960 24400 15972
rect 23584 15932 24400 15960
rect 9548 15864 12756 15892
rect 9548 15852 9554 15864
rect 14826 15852 14832 15904
rect 14884 15892 14890 15904
rect 14921 15895 14979 15901
rect 14921 15892 14933 15895
rect 14884 15864 14933 15892
rect 14884 15852 14890 15864
rect 14921 15861 14933 15864
rect 14967 15861 14979 15895
rect 14921 15855 14979 15861
rect 16298 15852 16304 15904
rect 16356 15892 16362 15904
rect 18506 15892 18512 15904
rect 16356 15864 18512 15892
rect 16356 15852 16362 15864
rect 18506 15852 18512 15864
rect 18564 15852 18570 15904
rect 20990 15852 20996 15904
rect 21048 15892 21054 15904
rect 21085 15895 21143 15901
rect 21085 15892 21097 15895
rect 21048 15864 21097 15892
rect 21048 15852 21054 15864
rect 21085 15861 21097 15864
rect 21131 15861 21143 15895
rect 21266 15892 21272 15904
rect 21227 15864 21272 15892
rect 21085 15855 21143 15861
rect 21266 15852 21272 15864
rect 21324 15852 21330 15904
rect 23106 15852 23112 15904
rect 23164 15892 23170 15904
rect 23201 15895 23259 15901
rect 23201 15892 23213 15895
rect 23164 15864 23213 15892
rect 23164 15852 23170 15864
rect 23201 15861 23213 15864
rect 23247 15892 23259 15895
rect 23584 15892 23612 15932
rect 24394 15920 24400 15932
rect 24452 15920 24458 15972
rect 24578 15920 24584 15972
rect 24636 15960 24642 15972
rect 24765 15963 24823 15969
rect 24765 15960 24777 15963
rect 24636 15932 24777 15960
rect 24636 15920 24642 15932
rect 24765 15929 24777 15932
rect 24811 15929 24823 15963
rect 24964 15960 24992 15991
rect 26436 15960 26464 15991
rect 27246 15988 27252 16000
rect 27304 15988 27310 16040
rect 27341 16031 27399 16037
rect 27341 15997 27353 16031
rect 27387 16028 27399 16031
rect 27522 16028 27528 16040
rect 27387 16000 27528 16028
rect 27387 15997 27399 16000
rect 27341 15991 27399 15997
rect 27522 15988 27528 16000
rect 27580 15988 27586 16040
rect 28077 16031 28135 16037
rect 28077 16028 28089 16031
rect 27632 16000 28089 16028
rect 24964 15932 26464 15960
rect 24765 15923 24823 15929
rect 23247 15864 23612 15892
rect 23247 15861 23259 15864
rect 23201 15855 23259 15861
rect 23658 15852 23664 15904
rect 23716 15892 23722 15904
rect 26234 15892 26240 15904
rect 23716 15864 26240 15892
rect 23716 15852 23722 15864
rect 26234 15852 26240 15864
rect 26292 15852 26298 15904
rect 27430 15892 27436 15904
rect 27391 15864 27436 15892
rect 27430 15852 27436 15864
rect 27488 15852 27494 15904
rect 27540 15892 27568 15988
rect 27632 15969 27660 16000
rect 28077 15997 28089 16000
rect 28123 15997 28135 16031
rect 28184 16028 28212 16068
rect 28261 16065 28273 16099
rect 28307 16096 28319 16099
rect 28994 16096 29000 16108
rect 28307 16068 29000 16096
rect 28307 16065 28319 16068
rect 28261 16059 28319 16065
rect 28994 16056 29000 16068
rect 29052 16056 29058 16108
rect 29181 16099 29239 16105
rect 29181 16065 29193 16099
rect 29227 16096 29239 16099
rect 29270 16096 29276 16108
rect 29227 16068 29276 16096
rect 29227 16065 29239 16068
rect 29181 16059 29239 16065
rect 29270 16056 29276 16068
rect 29328 16056 29334 16108
rect 29825 16099 29883 16105
rect 29825 16065 29837 16099
rect 29871 16096 29883 16099
rect 29914 16096 29920 16108
rect 29871 16068 29920 16096
rect 29871 16065 29883 16068
rect 29825 16059 29883 16065
rect 29914 16056 29920 16068
rect 29972 16056 29978 16108
rect 30092 16099 30150 16105
rect 30092 16065 30104 16099
rect 30138 16096 30150 16099
rect 30650 16096 30656 16108
rect 30138 16068 30656 16096
rect 30138 16065 30150 16068
rect 30092 16059 30150 16065
rect 30650 16056 30656 16068
rect 30708 16056 30714 16108
rect 28629 16031 28687 16037
rect 28629 16028 28641 16031
rect 28184 16000 28641 16028
rect 28077 15991 28135 15997
rect 28629 15997 28641 16000
rect 28675 15997 28687 16031
rect 28629 15991 28687 15997
rect 27617 15963 27675 15969
rect 27617 15929 27629 15963
rect 27663 15929 27675 15963
rect 27617 15923 27675 15929
rect 28442 15920 28448 15972
rect 28500 15960 28506 15972
rect 28537 15963 28595 15969
rect 28537 15960 28549 15963
rect 28500 15932 28549 15960
rect 28500 15920 28506 15932
rect 28537 15929 28549 15932
rect 28583 15929 28595 15963
rect 28537 15923 28595 15929
rect 28902 15892 28908 15904
rect 27540 15864 28908 15892
rect 28902 15852 28908 15864
rect 28960 15852 28966 15904
rect 1104 15802 32016 15824
rect 1104 15750 2136 15802
rect 2188 15750 12440 15802
rect 12492 15750 22744 15802
rect 22796 15750 32016 15802
rect 1104 15728 32016 15750
rect 1397 15691 1455 15697
rect 1397 15657 1409 15691
rect 1443 15688 1455 15691
rect 1486 15688 1492 15700
rect 1443 15660 1492 15688
rect 1443 15657 1455 15660
rect 1397 15651 1455 15657
rect 1486 15648 1492 15660
rect 1544 15648 1550 15700
rect 2590 15648 2596 15700
rect 2648 15688 2654 15700
rect 3789 15691 3847 15697
rect 3789 15688 3801 15691
rect 2648 15660 3801 15688
rect 2648 15648 2654 15660
rect 3789 15657 3801 15660
rect 3835 15657 3847 15691
rect 3789 15651 3847 15657
rect 4798 15648 4804 15700
rect 4856 15688 4862 15700
rect 4985 15691 5043 15697
rect 4985 15688 4997 15691
rect 4856 15660 4997 15688
rect 4856 15648 4862 15660
rect 4985 15657 4997 15660
rect 5031 15657 5043 15691
rect 7466 15688 7472 15700
rect 4985 15651 5043 15657
rect 5552 15660 7472 15688
rect 2866 15620 2872 15632
rect 2827 15592 2872 15620
rect 2866 15580 2872 15592
rect 2924 15580 2930 15632
rect 5074 15580 5080 15632
rect 5132 15620 5138 15632
rect 5552 15620 5580 15660
rect 7466 15648 7472 15660
rect 7524 15648 7530 15700
rect 7576 15660 13768 15688
rect 5132 15592 5580 15620
rect 5132 15580 5138 15592
rect 2041 15555 2099 15561
rect 2041 15521 2053 15555
rect 2087 15552 2099 15555
rect 3786 15552 3792 15564
rect 2087 15524 3792 15552
rect 2087 15521 2099 15524
rect 2041 15515 2099 15521
rect 3786 15512 3792 15524
rect 3844 15512 3850 15564
rect 4338 15552 4344 15564
rect 4299 15524 4344 15552
rect 4338 15512 4344 15524
rect 4396 15512 4402 15564
rect 5442 15552 5448 15564
rect 5403 15524 5448 15552
rect 5442 15512 5448 15524
rect 5500 15512 5506 15564
rect 5552 15561 5580 15592
rect 6273 15623 6331 15629
rect 6273 15589 6285 15623
rect 6319 15589 6331 15623
rect 6273 15583 6331 15589
rect 5537 15555 5595 15561
rect 5537 15521 5549 15555
rect 5583 15521 5595 15555
rect 6288 15552 6316 15583
rect 6638 15580 6644 15632
rect 6696 15620 6702 15632
rect 7101 15623 7159 15629
rect 6696 15592 7052 15620
rect 6696 15580 6702 15592
rect 6546 15552 6552 15564
rect 6288 15524 6552 15552
rect 5537 15515 5595 15521
rect 6546 15512 6552 15524
rect 6604 15512 6610 15564
rect 6822 15552 6828 15564
rect 6783 15524 6828 15552
rect 6822 15512 6828 15524
rect 6880 15512 6886 15564
rect 1765 15487 1823 15493
rect 1765 15453 1777 15487
rect 1811 15484 1823 15487
rect 1854 15484 1860 15496
rect 1811 15456 1860 15484
rect 1811 15453 1823 15456
rect 1765 15447 1823 15453
rect 1854 15444 1860 15456
rect 1912 15444 1918 15496
rect 2406 15444 2412 15496
rect 2464 15484 2470 15496
rect 2464 15456 6868 15484
rect 2464 15444 2470 15456
rect 0 15416 800 15430
rect 1486 15416 1492 15428
rect 0 15388 1492 15416
rect 0 15374 800 15388
rect 1486 15376 1492 15388
rect 1544 15376 1550 15428
rect 2314 15376 2320 15428
rect 2372 15416 2378 15428
rect 2593 15419 2651 15425
rect 2593 15416 2605 15419
rect 2372 15388 2605 15416
rect 2372 15376 2378 15388
rect 2593 15385 2605 15388
rect 2639 15385 2651 15419
rect 4157 15419 4215 15425
rect 4157 15416 4169 15419
rect 2593 15379 2651 15385
rect 2746 15388 4169 15416
rect 1857 15351 1915 15357
rect 1857 15317 1869 15351
rect 1903 15348 1915 15351
rect 2406 15348 2412 15360
rect 1903 15320 2412 15348
rect 1903 15317 1915 15320
rect 1857 15311 1915 15317
rect 2406 15308 2412 15320
rect 2464 15308 2470 15360
rect 2498 15308 2504 15360
rect 2556 15348 2562 15360
rect 2746 15348 2774 15388
rect 4157 15385 4169 15388
rect 4203 15385 4215 15419
rect 4157 15379 4215 15385
rect 4249 15419 4307 15425
rect 4249 15385 4261 15419
rect 4295 15416 4307 15419
rect 5353 15419 5411 15425
rect 4295 15388 4476 15416
rect 4295 15385 4307 15388
rect 4249 15379 4307 15385
rect 3050 15348 3056 15360
rect 2556 15320 2774 15348
rect 3011 15320 3056 15348
rect 2556 15308 2562 15320
rect 3050 15308 3056 15320
rect 3108 15308 3114 15360
rect 4448 15348 4476 15388
rect 5353 15385 5365 15419
rect 5399 15416 5411 15419
rect 5534 15416 5540 15428
rect 5399 15388 5540 15416
rect 5399 15385 5411 15388
rect 5353 15379 5411 15385
rect 5534 15376 5540 15388
rect 5592 15416 5598 15428
rect 6641 15419 6699 15425
rect 6641 15416 6653 15419
rect 5592 15388 6653 15416
rect 5592 15376 5598 15388
rect 6641 15385 6653 15388
rect 6687 15385 6699 15419
rect 6641 15379 6699 15385
rect 6270 15348 6276 15360
rect 4448 15320 6276 15348
rect 6270 15308 6276 15320
rect 6328 15348 6334 15360
rect 6730 15348 6736 15360
rect 6328 15320 6736 15348
rect 6328 15308 6334 15320
rect 6730 15308 6736 15320
rect 6788 15308 6794 15360
rect 6840 15348 6868 15456
rect 7024 15416 7052 15592
rect 7101 15589 7113 15623
rect 7147 15620 7159 15623
rect 7576 15620 7604 15660
rect 7147 15592 7604 15620
rect 7147 15589 7159 15592
rect 7101 15583 7159 15589
rect 7742 15580 7748 15632
rect 7800 15620 7806 15632
rect 8297 15623 8355 15629
rect 8297 15620 8309 15623
rect 7800 15592 8309 15620
rect 7800 15580 7806 15592
rect 8297 15589 8309 15592
rect 8343 15589 8355 15623
rect 8297 15583 8355 15589
rect 10502 15580 10508 15632
rect 10560 15620 10566 15632
rect 13633 15623 13691 15629
rect 13633 15620 13645 15623
rect 10560 15592 13645 15620
rect 10560 15580 10566 15592
rect 13633 15589 13645 15592
rect 13679 15589 13691 15623
rect 13740 15620 13768 15660
rect 13814 15648 13820 15700
rect 13872 15688 13878 15700
rect 15749 15691 15807 15697
rect 15749 15688 15761 15691
rect 13872 15660 15761 15688
rect 13872 15648 13878 15660
rect 15749 15657 15761 15660
rect 15795 15657 15807 15691
rect 15749 15651 15807 15657
rect 16482 15648 16488 15700
rect 16540 15688 16546 15700
rect 17954 15688 17960 15700
rect 16540 15660 17960 15688
rect 16540 15648 16546 15660
rect 17954 15648 17960 15660
rect 18012 15648 18018 15700
rect 18233 15691 18291 15697
rect 18233 15657 18245 15691
rect 18279 15688 18291 15691
rect 18322 15688 18328 15700
rect 18279 15660 18328 15688
rect 18279 15657 18291 15660
rect 18233 15651 18291 15657
rect 18322 15648 18328 15660
rect 18380 15648 18386 15700
rect 19518 15688 19524 15700
rect 19479 15660 19524 15688
rect 19518 15648 19524 15660
rect 19576 15648 19582 15700
rect 19886 15648 19892 15700
rect 19944 15688 19950 15700
rect 23658 15688 23664 15700
rect 19944 15660 23664 15688
rect 19944 15648 19950 15660
rect 23658 15648 23664 15660
rect 23716 15648 23722 15700
rect 23934 15648 23940 15700
rect 23992 15688 23998 15700
rect 24489 15691 24547 15697
rect 24489 15688 24501 15691
rect 23992 15660 24501 15688
rect 23992 15648 23998 15660
rect 24489 15657 24501 15660
rect 24535 15657 24547 15691
rect 24489 15651 24547 15657
rect 24949 15691 25007 15697
rect 24949 15657 24961 15691
rect 24995 15657 25007 15691
rect 24949 15651 25007 15657
rect 13740 15592 24256 15620
rect 13633 15583 13691 15589
rect 7285 15555 7343 15561
rect 7285 15521 7297 15555
rect 7331 15552 7343 15555
rect 8570 15552 8576 15564
rect 7331 15524 8576 15552
rect 7331 15521 7343 15524
rect 7285 15515 7343 15521
rect 8570 15512 8576 15524
rect 8628 15512 8634 15564
rect 8938 15552 8944 15564
rect 8899 15524 8944 15552
rect 8938 15512 8944 15524
rect 8996 15512 9002 15564
rect 13998 15552 14004 15564
rect 11164 15524 14004 15552
rect 7190 15444 7196 15496
rect 7248 15484 7254 15496
rect 11164 15493 11192 15524
rect 13998 15512 14004 15524
rect 14056 15512 14062 15564
rect 14108 15524 16611 15552
rect 8205 15487 8263 15493
rect 8205 15484 8217 15487
rect 7248 15456 8217 15484
rect 7248 15444 7254 15456
rect 8205 15453 8217 15456
rect 8251 15453 8263 15487
rect 8205 15447 8263 15453
rect 11149 15487 11207 15493
rect 11149 15453 11161 15487
rect 11195 15453 11207 15487
rect 11149 15447 11207 15453
rect 11333 15487 11391 15493
rect 11333 15453 11345 15487
rect 11379 15453 11391 15487
rect 11333 15447 11391 15453
rect 7285 15419 7343 15425
rect 7285 15416 7297 15419
rect 7024 15388 7297 15416
rect 7285 15385 7297 15388
rect 7331 15385 7343 15419
rect 7285 15379 7343 15385
rect 7561 15419 7619 15425
rect 7561 15385 7573 15419
rect 7607 15416 7619 15419
rect 8478 15416 8484 15428
rect 7607 15388 8484 15416
rect 7607 15385 7619 15388
rect 7561 15379 7619 15385
rect 8478 15376 8484 15388
rect 8536 15376 8542 15428
rect 9208 15419 9266 15425
rect 9208 15385 9220 15419
rect 9254 15416 9266 15419
rect 9306 15416 9312 15428
rect 9254 15388 9312 15416
rect 9254 15385 9266 15388
rect 9208 15379 9266 15385
rect 9306 15376 9312 15388
rect 9364 15376 9370 15428
rect 11348 15416 11376 15447
rect 11422 15444 11428 15496
rect 11480 15484 11486 15496
rect 11885 15487 11943 15493
rect 11480 15456 11525 15484
rect 11480 15444 11486 15456
rect 11885 15453 11897 15487
rect 11931 15453 11943 15487
rect 11885 15447 11943 15453
rect 11790 15416 11796 15428
rect 11348 15388 11796 15416
rect 11790 15376 11796 15388
rect 11848 15376 11854 15428
rect 11900 15416 11928 15447
rect 11974 15444 11980 15496
rect 12032 15484 12038 15496
rect 12161 15487 12219 15493
rect 12161 15484 12173 15487
rect 12032 15456 12173 15484
rect 12032 15444 12038 15456
rect 12161 15453 12173 15456
rect 12207 15484 12219 15487
rect 12342 15484 12348 15496
rect 12207 15456 12348 15484
rect 12207 15453 12219 15456
rect 12161 15447 12219 15453
rect 12342 15444 12348 15456
rect 12400 15444 12406 15496
rect 13357 15487 13415 15493
rect 13357 15453 13369 15487
rect 13403 15484 13415 15487
rect 13633 15487 13691 15493
rect 13633 15484 13645 15487
rect 13403 15456 13645 15484
rect 13403 15453 13415 15456
rect 13357 15447 13415 15453
rect 13633 15453 13645 15456
rect 13679 15453 13691 15487
rect 13633 15447 13691 15453
rect 13725 15487 13783 15493
rect 13725 15453 13737 15487
rect 13771 15484 13783 15487
rect 14108 15484 14136 15524
rect 13771 15456 14136 15484
rect 13771 15453 13783 15456
rect 13725 15447 13783 15453
rect 14182 15444 14188 15496
rect 14240 15484 14246 15496
rect 14458 15484 14464 15496
rect 14240 15456 14464 15484
rect 14240 15444 14246 15456
rect 14458 15444 14464 15456
rect 14516 15444 14522 15496
rect 15930 15444 15936 15496
rect 15988 15484 15994 15496
rect 16482 15484 16488 15496
rect 15988 15456 16488 15484
rect 15988 15444 15994 15456
rect 16482 15444 16488 15456
rect 16540 15444 16546 15496
rect 13170 15416 13176 15428
rect 11900 15388 13176 15416
rect 13170 15376 13176 15388
rect 13228 15416 13234 15428
rect 13541 15419 13599 15425
rect 13541 15416 13553 15419
rect 13228 15388 13553 15416
rect 13228 15376 13234 15388
rect 13541 15385 13553 15388
rect 13587 15416 13599 15419
rect 16583 15416 16611 15524
rect 17034 15512 17040 15564
rect 17092 15552 17098 15564
rect 17221 15555 17279 15561
rect 17221 15552 17233 15555
rect 17092 15524 17233 15552
rect 17092 15512 17098 15524
rect 17221 15521 17233 15524
rect 17267 15521 17279 15555
rect 17862 15552 17868 15564
rect 17823 15524 17868 15552
rect 17221 15515 17279 15521
rect 17862 15512 17868 15524
rect 17920 15512 17926 15564
rect 17954 15512 17960 15564
rect 18012 15552 18018 15564
rect 18690 15552 18696 15564
rect 18012 15524 18696 15552
rect 18012 15512 18018 15524
rect 18690 15512 18696 15524
rect 18748 15512 18754 15564
rect 20346 15552 20352 15564
rect 19720 15524 20352 15552
rect 19720 15496 19748 15524
rect 20346 15512 20352 15524
rect 20404 15512 20410 15564
rect 22922 15512 22928 15564
rect 22980 15552 22986 15564
rect 23106 15552 23112 15564
rect 22980 15524 23112 15552
rect 22980 15512 22986 15524
rect 23106 15512 23112 15524
rect 23164 15512 23170 15564
rect 23385 15555 23443 15561
rect 23385 15521 23397 15555
rect 23431 15552 23443 15555
rect 24228 15552 24256 15592
rect 24762 15580 24768 15632
rect 24820 15620 24826 15632
rect 24964 15620 24992 15651
rect 25590 15648 25596 15700
rect 25648 15688 25654 15700
rect 28994 15688 29000 15700
rect 25648 15660 28028 15688
rect 28955 15660 29000 15688
rect 25648 15648 25654 15660
rect 28000 15629 28028 15660
rect 28994 15648 29000 15660
rect 29052 15648 29058 15700
rect 30558 15648 30564 15700
rect 30616 15688 30622 15700
rect 30653 15691 30711 15697
rect 30653 15688 30665 15691
rect 30616 15660 30665 15688
rect 30616 15648 30622 15660
rect 30653 15657 30665 15660
rect 30699 15657 30711 15691
rect 30653 15651 30711 15657
rect 27985 15623 28043 15629
rect 24820 15592 24992 15620
rect 26620 15592 27752 15620
rect 24820 15580 24826 15592
rect 23431 15524 24164 15552
rect 24228 15524 25728 15552
rect 23431 15521 23443 15524
rect 23385 15515 23443 15521
rect 17129 15487 17187 15493
rect 17129 15453 17141 15487
rect 17175 15484 17187 15487
rect 17678 15484 17684 15496
rect 17175 15456 17684 15484
rect 17175 15453 17187 15456
rect 17129 15447 17187 15453
rect 17678 15444 17684 15456
rect 17736 15444 17742 15496
rect 18049 15487 18107 15493
rect 18049 15453 18061 15487
rect 18095 15484 18107 15487
rect 18782 15484 18788 15496
rect 18095 15456 18788 15484
rect 18095 15453 18107 15456
rect 18049 15447 18107 15453
rect 18782 15444 18788 15456
rect 18840 15444 18846 15496
rect 19702 15484 19708 15496
rect 19615 15456 19708 15484
rect 19702 15444 19708 15456
rect 19760 15444 19766 15496
rect 19978 15484 19984 15496
rect 19939 15456 19984 15484
rect 19978 15444 19984 15456
rect 20036 15444 20042 15496
rect 20165 15487 20223 15493
rect 20165 15453 20177 15487
rect 20211 15484 20223 15487
rect 20254 15484 20260 15496
rect 20211 15456 20260 15484
rect 20211 15453 20223 15456
rect 20165 15447 20223 15453
rect 20254 15444 20260 15456
rect 20312 15444 20318 15496
rect 20806 15484 20812 15496
rect 20767 15456 20812 15484
rect 20806 15444 20812 15456
rect 20864 15444 20870 15496
rect 23569 15487 23627 15493
rect 23569 15453 23581 15487
rect 23615 15453 23627 15487
rect 23750 15484 23756 15496
rect 23711 15456 23756 15484
rect 23569 15447 23627 15453
rect 17037 15419 17095 15425
rect 17037 15416 17049 15419
rect 13587 15388 14228 15416
rect 16583 15388 17049 15416
rect 13587 15385 13599 15388
rect 13541 15379 13599 15385
rect 14200 15360 14228 15388
rect 17037 15385 17049 15388
rect 17083 15416 17095 15419
rect 19242 15416 19248 15428
rect 17083 15388 19248 15416
rect 17083 15385 17095 15388
rect 17037 15379 17095 15385
rect 19242 15376 19248 15388
rect 19300 15376 19306 15428
rect 23382 15416 23388 15428
rect 21928 15388 23388 15416
rect 7101 15351 7159 15357
rect 7101 15348 7113 15351
rect 6840 15320 7113 15348
rect 7101 15317 7113 15320
rect 7147 15317 7159 15351
rect 7650 15348 7656 15360
rect 7611 15320 7656 15348
rect 7101 15311 7159 15317
rect 7650 15308 7656 15320
rect 7708 15308 7714 15360
rect 10321 15351 10379 15357
rect 10321 15317 10333 15351
rect 10367 15348 10379 15351
rect 10502 15348 10508 15360
rect 10367 15320 10508 15348
rect 10367 15317 10379 15320
rect 10321 15311 10379 15317
rect 10502 15308 10508 15320
rect 10560 15308 10566 15360
rect 10965 15351 11023 15357
rect 10965 15317 10977 15351
rect 11011 15348 11023 15351
rect 12158 15348 12164 15360
rect 11011 15320 12164 15348
rect 11011 15317 11023 15320
rect 10965 15311 11023 15317
rect 12158 15308 12164 15320
rect 12216 15308 12222 15360
rect 13633 15351 13691 15357
rect 13633 15317 13645 15351
rect 13679 15348 13691 15351
rect 14093 15351 14151 15357
rect 14093 15348 14105 15351
rect 13679 15320 14105 15348
rect 13679 15317 13691 15320
rect 13633 15311 13691 15317
rect 14093 15317 14105 15320
rect 14139 15317 14151 15351
rect 14093 15311 14151 15317
rect 14182 15308 14188 15360
rect 14240 15308 14246 15360
rect 14277 15351 14335 15357
rect 14277 15317 14289 15351
rect 14323 15348 14335 15351
rect 16206 15348 16212 15360
rect 14323 15320 16212 15348
rect 14323 15317 14335 15320
rect 14277 15311 14335 15317
rect 16206 15308 16212 15320
rect 16264 15308 16270 15360
rect 16669 15351 16727 15357
rect 16669 15317 16681 15351
rect 16715 15348 16727 15351
rect 16850 15348 16856 15360
rect 16715 15320 16856 15348
rect 16715 15317 16727 15320
rect 16669 15311 16727 15317
rect 16850 15308 16856 15320
rect 16908 15308 16914 15360
rect 19518 15308 19524 15360
rect 19576 15348 19582 15360
rect 21928 15348 21956 15388
rect 23382 15376 23388 15388
rect 23440 15376 23446 15428
rect 23584 15416 23612 15447
rect 23750 15444 23756 15456
rect 23808 15444 23814 15496
rect 23860 15493 24072 15494
rect 23845 15487 24087 15493
rect 23845 15453 23857 15487
rect 23891 15466 24041 15487
rect 23891 15453 23903 15466
rect 23845 15447 23903 15453
rect 24029 15453 24041 15466
rect 24075 15453 24087 15487
rect 24029 15447 24087 15453
rect 23658 15416 23664 15428
rect 23584 15388 23664 15416
rect 23658 15376 23664 15388
rect 23716 15376 23722 15428
rect 24136 15416 24164 15524
rect 24302 15444 24308 15496
rect 24360 15484 24366 15496
rect 24397 15487 24455 15493
rect 24397 15484 24409 15487
rect 24360 15456 24409 15484
rect 24360 15444 24366 15456
rect 24397 15453 24409 15456
rect 24443 15453 24455 15487
rect 24762 15484 24768 15496
rect 24723 15456 24768 15484
rect 24397 15447 24455 15453
rect 24762 15444 24768 15456
rect 24820 15444 24826 15496
rect 25590 15484 25596 15496
rect 25551 15456 25596 15484
rect 25590 15444 25596 15456
rect 25648 15444 25654 15496
rect 25700 15484 25728 15524
rect 26620 15484 26648 15592
rect 27525 15555 27583 15561
rect 27525 15521 27537 15555
rect 27571 15552 27583 15555
rect 27614 15552 27620 15564
rect 27571 15524 27620 15552
rect 27571 15521 27583 15524
rect 27525 15515 27583 15521
rect 27614 15512 27620 15524
rect 27672 15512 27678 15564
rect 27724 15552 27752 15592
rect 27985 15589 27997 15623
rect 28031 15589 28043 15623
rect 27985 15583 28043 15589
rect 30374 15580 30380 15632
rect 30432 15620 30438 15632
rect 31021 15623 31079 15629
rect 31021 15620 31033 15623
rect 30432 15592 31033 15620
rect 30432 15580 30438 15592
rect 31021 15589 31033 15592
rect 31067 15589 31079 15623
rect 31021 15583 31079 15589
rect 27724 15524 31754 15552
rect 27706 15484 27712 15496
rect 25700 15456 26648 15484
rect 27667 15456 27712 15484
rect 27706 15444 27712 15456
rect 27764 15444 27770 15496
rect 28077 15487 28135 15493
rect 28077 15453 28089 15487
rect 28123 15453 28135 15487
rect 28629 15487 28687 15493
rect 28629 15484 28641 15487
rect 28077 15447 28135 15453
rect 28184 15456 28641 15484
rect 24854 15416 24860 15428
rect 24136 15388 24860 15416
rect 24854 15376 24860 15388
rect 24912 15376 24918 15428
rect 25860 15419 25918 15425
rect 25860 15385 25872 15419
rect 25906 15416 25918 15419
rect 26878 15416 26884 15428
rect 25906 15388 26884 15416
rect 25906 15385 25918 15388
rect 25860 15379 25918 15385
rect 26878 15376 26884 15388
rect 26936 15376 26942 15428
rect 27246 15376 27252 15428
rect 27304 15416 27310 15428
rect 28092 15416 28120 15447
rect 27304 15388 28120 15416
rect 27304 15376 27310 15388
rect 19576 15320 21956 15348
rect 19576 15308 19582 15320
rect 22002 15308 22008 15360
rect 22060 15348 22066 15360
rect 22097 15351 22155 15357
rect 22097 15348 22109 15351
rect 22060 15320 22109 15348
rect 22060 15308 22066 15320
rect 22097 15317 22109 15320
rect 22143 15348 22155 15351
rect 22830 15348 22836 15360
rect 22143 15320 22836 15348
rect 22143 15317 22155 15320
rect 22097 15311 22155 15317
rect 22830 15308 22836 15320
rect 22888 15308 22894 15360
rect 24029 15351 24087 15357
rect 24029 15317 24041 15351
rect 24075 15348 24087 15351
rect 25774 15348 25780 15360
rect 24075 15320 25780 15348
rect 24075 15317 24087 15320
rect 24029 15311 24087 15317
rect 25774 15308 25780 15320
rect 25832 15308 25838 15360
rect 26970 15348 26976 15360
rect 26931 15320 26976 15348
rect 26970 15308 26976 15320
rect 27028 15348 27034 15360
rect 28184 15348 28212 15456
rect 28629 15453 28641 15456
rect 28675 15453 28687 15487
rect 28629 15447 28687 15453
rect 28721 15487 28779 15493
rect 28721 15453 28733 15487
rect 28767 15453 28779 15487
rect 28721 15447 28779 15453
rect 28813 15487 28871 15493
rect 28813 15453 28825 15487
rect 28859 15484 28871 15487
rect 28902 15484 28908 15496
rect 28859 15456 28908 15484
rect 28859 15453 28871 15456
rect 28813 15447 28871 15453
rect 28258 15376 28264 15428
rect 28316 15416 28322 15428
rect 28736 15416 28764 15447
rect 28902 15444 28908 15456
rect 28960 15444 28966 15496
rect 29733 15487 29791 15493
rect 29733 15453 29745 15487
rect 29779 15484 29791 15487
rect 29822 15484 29828 15496
rect 29779 15456 29828 15484
rect 29779 15453 29791 15456
rect 29733 15447 29791 15453
rect 29822 15444 29828 15456
rect 29880 15444 29886 15496
rect 30006 15484 30012 15496
rect 29967 15456 30012 15484
rect 30006 15444 30012 15456
rect 30064 15444 30070 15496
rect 30190 15484 30196 15496
rect 30151 15456 30196 15484
rect 30190 15444 30196 15456
rect 30248 15444 30254 15496
rect 30834 15484 30840 15496
rect 30795 15456 30840 15484
rect 30834 15444 30840 15456
rect 30892 15444 30898 15496
rect 31110 15444 31116 15496
rect 31168 15484 31174 15496
rect 31168 15456 31213 15484
rect 31168 15444 31174 15456
rect 29549 15419 29607 15425
rect 29549 15416 29561 15419
rect 28316 15388 28764 15416
rect 28828 15388 29561 15416
rect 28316 15376 28322 15388
rect 27028 15320 28212 15348
rect 27028 15308 27034 15320
rect 28718 15308 28724 15360
rect 28776 15348 28782 15360
rect 28828 15348 28856 15388
rect 29549 15385 29561 15388
rect 29595 15385 29607 15419
rect 31726 15416 31754 15524
rect 32320 15416 33120 15430
rect 31726 15388 33120 15416
rect 29549 15379 29607 15385
rect 32320 15374 33120 15388
rect 28776 15320 28856 15348
rect 28776 15308 28782 15320
rect 1104 15258 32016 15280
rect 1104 15206 7288 15258
rect 7340 15206 17592 15258
rect 17644 15206 27896 15258
rect 27948 15206 32016 15258
rect 1104 15184 32016 15206
rect 1670 15104 1676 15156
rect 1728 15144 1734 15156
rect 2222 15144 2228 15156
rect 1728 15116 2228 15144
rect 1728 15104 1734 15116
rect 2222 15104 2228 15116
rect 2280 15144 2286 15156
rect 2593 15147 2651 15153
rect 2593 15144 2605 15147
rect 2280 15116 2605 15144
rect 2280 15104 2286 15116
rect 2593 15113 2605 15116
rect 2639 15113 2651 15147
rect 2593 15107 2651 15113
rect 2866 15104 2872 15156
rect 2924 15144 2930 15156
rect 3878 15144 3884 15156
rect 2924 15116 3884 15144
rect 2924 15104 2930 15116
rect 3878 15104 3884 15116
rect 3936 15104 3942 15156
rect 3970 15104 3976 15156
rect 4028 15104 4034 15156
rect 4341 15147 4399 15153
rect 4341 15113 4353 15147
rect 4387 15144 4399 15147
rect 4890 15144 4896 15156
rect 4387 15116 4896 15144
rect 4387 15113 4399 15116
rect 4341 15107 4399 15113
rect 4890 15104 4896 15116
rect 4948 15144 4954 15156
rect 5442 15144 5448 15156
rect 4948 15116 5448 15144
rect 4948 15104 4954 15116
rect 5442 15104 5448 15116
rect 5500 15104 5506 15156
rect 5813 15147 5871 15153
rect 5813 15113 5825 15147
rect 5859 15113 5871 15147
rect 5813 15107 5871 15113
rect 1486 15076 1492 15088
rect 1447 15048 1492 15076
rect 1486 15036 1492 15048
rect 1544 15036 1550 15088
rect 2314 15036 2320 15088
rect 2372 15076 2378 15088
rect 3988 15076 4016 15104
rect 5828 15076 5856 15107
rect 6086 15104 6092 15156
rect 6144 15144 6150 15156
rect 14090 15144 14096 15156
rect 6144 15116 14096 15144
rect 6144 15104 6150 15116
rect 14090 15104 14096 15116
rect 14148 15104 14154 15156
rect 14918 15104 14924 15156
rect 14976 15144 14982 15156
rect 15381 15147 15439 15153
rect 14976 15116 15148 15144
rect 14976 15104 14982 15116
rect 6822 15076 6828 15088
rect 2372 15048 2636 15076
rect 2372 15036 2378 15048
rect 1026 14968 1032 15020
rect 1084 15008 1090 15020
rect 1670 15008 1676 15020
rect 1084 14980 1676 15008
rect 1084 14968 1090 14980
rect 1670 14968 1676 14980
rect 1728 14968 1734 15020
rect 2498 15008 2504 15020
rect 2459 14980 2504 15008
rect 2498 14968 2504 14980
rect 2556 14968 2562 15020
rect 1946 14900 1952 14952
rect 2004 14940 2010 14952
rect 2608 14940 2636 15048
rect 3804 15048 5212 15076
rect 5828 15048 6828 15076
rect 3513 15011 3571 15017
rect 3513 14977 3525 15011
rect 3559 15008 3571 15011
rect 3602 15008 3608 15020
rect 3559 14980 3608 15008
rect 3559 14977 3571 14980
rect 3513 14971 3571 14977
rect 3602 14968 3608 14980
rect 3660 14968 3666 15020
rect 3804 15017 3832 15048
rect 3789 15011 3847 15017
rect 3789 14977 3801 15011
rect 3835 14977 3847 15011
rect 3970 15008 3976 15020
rect 3931 14980 3976 15008
rect 3789 14971 3847 14977
rect 3970 14968 3976 14980
rect 4028 14968 4034 15020
rect 4700 15011 4758 15017
rect 4700 14977 4712 15011
rect 4746 15008 4758 15011
rect 5074 15008 5080 15020
rect 4746 14980 5080 15008
rect 4746 14977 4758 14980
rect 4700 14971 4758 14977
rect 5074 14968 5080 14980
rect 5132 14968 5138 15020
rect 5184 15008 5212 15048
rect 6822 15036 6828 15048
rect 6880 15036 6886 15088
rect 8938 15076 8944 15088
rect 7852 15048 8944 15076
rect 7650 15008 7656 15020
rect 5184 14980 7656 15008
rect 7650 14968 7656 14980
rect 7708 14968 7714 15020
rect 7852 15017 7880 15048
rect 8938 15036 8944 15048
rect 8996 15036 9002 15088
rect 11330 15076 11336 15088
rect 10244 15048 11336 15076
rect 7837 15011 7895 15017
rect 7837 14977 7849 15011
rect 7883 14977 7895 15011
rect 8093 15011 8151 15017
rect 8093 15008 8105 15011
rect 7837 14971 7895 14977
rect 7944 14980 8105 15008
rect 2777 14943 2835 14949
rect 2777 14940 2789 14943
rect 2004 14912 2544 14940
rect 2608 14912 2789 14940
rect 2004 14900 2010 14912
rect 1673 14875 1731 14881
rect 1673 14841 1685 14875
rect 1719 14872 1731 14875
rect 2516 14872 2544 14912
rect 2777 14909 2789 14912
rect 2823 14940 2835 14943
rect 3988 14940 4016 14968
rect 4430 14940 4436 14952
rect 2823 14912 4016 14940
rect 4391 14912 4436 14940
rect 2823 14909 2835 14912
rect 2777 14903 2835 14909
rect 4430 14900 4436 14912
rect 4488 14900 4494 14952
rect 7006 14900 7012 14952
rect 7064 14940 7070 14952
rect 7944 14940 7972 14980
rect 8093 14977 8105 14980
rect 8139 14977 8151 15011
rect 8093 14971 8151 14977
rect 8386 14968 8392 15020
rect 8444 15008 8450 15020
rect 10042 15008 10048 15020
rect 8444 14980 8892 15008
rect 10003 14980 10048 15008
rect 8444 14968 8450 14980
rect 7064 14912 7972 14940
rect 7064 14900 7070 14912
rect 3329 14875 3387 14881
rect 3329 14872 3341 14875
rect 1719 14844 2452 14872
rect 2516 14844 3341 14872
rect 1719 14841 1731 14844
rect 1673 14835 1731 14841
rect 1854 14764 1860 14816
rect 1912 14804 1918 14816
rect 2133 14807 2191 14813
rect 2133 14804 2145 14807
rect 1912 14776 2145 14804
rect 1912 14764 1918 14776
rect 2133 14773 2145 14776
rect 2179 14773 2191 14807
rect 2424 14804 2452 14844
rect 3329 14841 3341 14844
rect 3375 14841 3387 14875
rect 4341 14875 4399 14881
rect 4341 14872 4353 14875
rect 3329 14835 3387 14841
rect 3436 14844 4353 14872
rect 3436 14804 3464 14844
rect 4341 14841 4353 14844
rect 4387 14841 4399 14875
rect 7742 14872 7748 14884
rect 4341 14835 4399 14841
rect 6840 14844 7748 14872
rect 2424 14776 3464 14804
rect 2133 14767 2191 14773
rect 3510 14764 3516 14816
rect 3568 14804 3574 14816
rect 6840 14804 6868 14844
rect 7742 14832 7748 14844
rect 7800 14832 7806 14884
rect 8864 14872 8892 14980
rect 10042 14968 10048 14980
rect 10100 14968 10106 15020
rect 9214 14900 9220 14952
rect 9272 14940 9278 14952
rect 10244 14940 10272 15048
rect 11330 15036 11336 15048
rect 11388 15036 11394 15088
rect 12158 15085 12164 15088
rect 12152 15076 12164 15085
rect 12119 15048 12164 15076
rect 12152 15039 12164 15048
rect 12158 15036 12164 15039
rect 12216 15036 12222 15088
rect 15120 15076 15148 15116
rect 15381 15113 15393 15147
rect 15427 15144 15439 15147
rect 15654 15144 15660 15156
rect 15427 15116 15660 15144
rect 15427 15113 15439 15116
rect 15381 15107 15439 15113
rect 15654 15104 15660 15116
rect 15712 15104 15718 15156
rect 16025 15147 16083 15153
rect 16025 15113 16037 15147
rect 16071 15144 16083 15147
rect 16206 15144 16212 15156
rect 16071 15116 16212 15144
rect 16071 15113 16083 15116
rect 16025 15107 16083 15113
rect 16206 15104 16212 15116
rect 16264 15104 16270 15156
rect 16485 15147 16543 15153
rect 16485 15113 16497 15147
rect 16531 15144 16543 15147
rect 16942 15144 16948 15156
rect 16531 15116 16948 15144
rect 16531 15113 16543 15116
rect 16485 15107 16543 15113
rect 16942 15104 16948 15116
rect 17000 15104 17006 15156
rect 17037 15147 17095 15153
rect 17037 15113 17049 15147
rect 17083 15144 17095 15147
rect 17770 15144 17776 15156
rect 17083 15116 17776 15144
rect 17083 15113 17095 15116
rect 17037 15107 17095 15113
rect 17770 15104 17776 15116
rect 17828 15104 17834 15156
rect 17865 15147 17923 15153
rect 17865 15113 17877 15147
rect 17911 15144 17923 15147
rect 18138 15144 18144 15156
rect 17911 15116 18144 15144
rect 17911 15113 17923 15116
rect 17865 15107 17923 15113
rect 18138 15104 18144 15116
rect 18196 15104 18202 15156
rect 20990 15144 20996 15156
rect 19996 15116 20996 15144
rect 15473 15079 15531 15085
rect 15473 15076 15485 15079
rect 12268 15048 15047 15076
rect 15120 15048 15485 15076
rect 10321 15011 10379 15017
rect 10321 14977 10333 15011
rect 10367 14977 10379 15011
rect 10502 15008 10508 15020
rect 10463 14980 10508 15008
rect 10321 14971 10379 14977
rect 9272 14912 10272 14940
rect 10336 14940 10364 14971
rect 10502 14968 10508 14980
rect 10560 14968 10566 15020
rect 11238 14968 11244 15020
rect 11296 15008 11302 15020
rect 12268 15008 12296 15048
rect 11296 14980 12296 15008
rect 11296 14968 11302 14980
rect 13814 14968 13820 15020
rect 13872 15008 13878 15020
rect 14001 15011 14059 15017
rect 14001 15008 14013 15011
rect 13872 14980 14013 15008
rect 13872 14968 13878 14980
rect 14001 14977 14013 14980
rect 14047 14977 14059 15011
rect 14001 14971 14059 14977
rect 14268 15011 14326 15017
rect 14268 14977 14280 15011
rect 14314 15008 14326 15011
rect 14642 15008 14648 15020
rect 14314 14980 14648 15008
rect 14314 14977 14326 14980
rect 14268 14971 14326 14977
rect 14642 14968 14648 14980
rect 14700 14968 14706 15020
rect 11054 14940 11060 14952
rect 10336 14912 11060 14940
rect 9272 14900 9278 14912
rect 11054 14900 11060 14912
rect 11112 14900 11118 14952
rect 11882 14940 11888 14952
rect 11843 14912 11888 14940
rect 11882 14900 11888 14912
rect 11940 14900 11946 14952
rect 15019 14940 15047 15048
rect 15473 15045 15485 15048
rect 15519 15045 15531 15079
rect 15473 15039 15531 15045
rect 15838 15036 15844 15088
rect 15896 15076 15902 15088
rect 19996 15085 20024 15116
rect 20990 15104 20996 15116
rect 21048 15104 21054 15156
rect 22094 15104 22100 15156
rect 22152 15144 22158 15156
rect 22152 15116 22197 15144
rect 22152 15104 22158 15116
rect 23658 15104 23664 15156
rect 23716 15144 23722 15156
rect 24026 15144 24032 15156
rect 23716 15116 24032 15144
rect 23716 15104 23722 15116
rect 24026 15104 24032 15116
rect 24084 15104 24090 15156
rect 27430 15144 27436 15156
rect 24228 15116 27436 15144
rect 19797 15079 19855 15085
rect 19797 15076 19809 15079
rect 15896 15048 19809 15076
rect 15896 15036 15902 15048
rect 19797 15045 19809 15048
rect 19843 15045 19855 15079
rect 19797 15039 19855 15045
rect 19981 15079 20039 15085
rect 19981 15045 19993 15079
rect 20027 15045 20039 15079
rect 19981 15039 20039 15045
rect 20254 15036 20260 15088
rect 20312 15076 20318 15088
rect 20312 15048 21036 15076
rect 20312 15036 20318 15048
rect 15102 14968 15108 15020
rect 15160 15008 15166 15020
rect 15933 15011 15991 15017
rect 15933 15008 15945 15011
rect 15160 14980 15945 15008
rect 15160 14968 15166 14980
rect 15933 14977 15945 14980
rect 15979 14977 15991 15011
rect 15933 14971 15991 14977
rect 16114 14968 16120 15020
rect 16172 15008 16178 15020
rect 16485 15011 16543 15017
rect 16485 15008 16497 15011
rect 16172 14980 16497 15008
rect 16172 14968 16178 14980
rect 16485 14977 16497 14980
rect 16531 14977 16543 15011
rect 16758 15008 16764 15020
rect 16719 14980 16764 15008
rect 16485 14971 16543 14977
rect 16758 14968 16764 14980
rect 16816 14968 16822 15020
rect 16853 15011 16911 15017
rect 16853 14977 16865 15011
rect 16899 15008 16911 15011
rect 16942 15008 16948 15020
rect 16899 14980 16948 15008
rect 16899 14977 16911 14980
rect 16853 14971 16911 14977
rect 16942 14968 16948 14980
rect 17000 14968 17006 15020
rect 17865 15011 17923 15017
rect 17865 15008 17877 15011
rect 17420 14980 17877 15008
rect 17420 14940 17448 14980
rect 17865 14977 17877 14980
rect 17911 14977 17923 15011
rect 17865 14971 17923 14977
rect 17957 15011 18015 15017
rect 17957 14977 17969 15011
rect 18003 15008 18015 15011
rect 18506 15008 18512 15020
rect 18003 14980 18512 15008
rect 18003 14977 18015 14980
rect 17957 14971 18015 14977
rect 18506 14968 18512 14980
rect 18564 14968 18570 15020
rect 18874 15008 18880 15020
rect 18835 14980 18880 15008
rect 18874 14968 18880 14980
rect 18932 14968 18938 15020
rect 20898 15008 20904 15020
rect 20859 14980 20904 15008
rect 20898 14968 20904 14980
rect 20956 14968 20962 15020
rect 21008 15017 21036 15048
rect 22186 15036 22192 15088
rect 22244 15076 22250 15088
rect 22244 15048 22508 15076
rect 22244 15036 22250 15048
rect 20993 15011 21051 15017
rect 20993 14977 21005 15011
rect 21039 14977 21051 15011
rect 20993 14971 21051 14977
rect 21085 15011 21143 15017
rect 21085 14977 21097 15011
rect 21131 15008 21143 15011
rect 21266 15008 21272 15020
rect 21131 14980 21272 15008
rect 21131 14977 21143 14980
rect 21085 14971 21143 14977
rect 21266 14968 21272 14980
rect 21324 14968 21330 15020
rect 22278 15008 22284 15020
rect 22239 14980 22284 15008
rect 22278 14968 22284 14980
rect 22336 14968 22342 15020
rect 22480 15017 22508 15048
rect 23124 15048 23888 15076
rect 23124 15017 23152 15048
rect 23382 15017 23388 15020
rect 22465 15011 22523 15017
rect 22465 14977 22477 15011
rect 22511 14977 22523 15011
rect 22465 14971 22523 14977
rect 23109 15011 23167 15017
rect 23109 14977 23121 15011
rect 23155 14977 23167 15011
rect 23109 14971 23167 14977
rect 23376 14971 23388 15017
rect 23440 15008 23446 15020
rect 23860 15008 23888 15048
rect 23934 15036 23940 15088
rect 23992 15076 23998 15088
rect 24228 15076 24256 15116
rect 27430 15104 27436 15116
rect 27488 15104 27494 15156
rect 27617 15147 27675 15153
rect 27617 15113 27629 15147
rect 27663 15144 27675 15147
rect 27706 15144 27712 15156
rect 27663 15116 27712 15144
rect 27663 15113 27675 15116
rect 27617 15107 27675 15113
rect 27706 15104 27712 15116
rect 27764 15104 27770 15156
rect 29362 15104 29368 15156
rect 29420 15144 29426 15156
rect 29733 15147 29791 15153
rect 29733 15144 29745 15147
rect 29420 15116 29745 15144
rect 29420 15104 29426 15116
rect 29733 15113 29745 15116
rect 29779 15144 29791 15147
rect 30190 15144 30196 15156
rect 29779 15116 30196 15144
rect 29779 15113 29791 15116
rect 29733 15107 29791 15113
rect 30190 15104 30196 15116
rect 30248 15104 30254 15156
rect 30650 15144 30656 15156
rect 30611 15116 30656 15144
rect 30650 15104 30656 15116
rect 30708 15104 30714 15156
rect 24946 15076 24952 15088
rect 23992 15048 24256 15076
rect 24780 15048 24952 15076
rect 23992 15036 23998 15048
rect 24780 15020 24808 15048
rect 24946 15036 24952 15048
rect 25004 15076 25010 15088
rect 25590 15076 25596 15088
rect 25004 15048 25596 15076
rect 25004 15036 25010 15048
rect 25590 15036 25596 15048
rect 25648 15036 25654 15088
rect 26326 15036 26332 15088
rect 26384 15076 26390 15088
rect 28258 15076 28264 15088
rect 26384 15048 28264 15076
rect 26384 15036 26390 15048
rect 28258 15036 28264 15048
rect 28316 15036 28322 15088
rect 28994 15076 29000 15088
rect 28368 15048 29000 15076
rect 24762 15008 24768 15020
rect 23440 14980 23476 15008
rect 23860 15006 24164 15008
rect 24228 15006 24768 15008
rect 23860 14980 24768 15006
rect 23382 14968 23388 14971
rect 23440 14968 23446 14980
rect 24136 14978 24256 14980
rect 24762 14968 24768 14980
rect 24820 14968 24826 15020
rect 24857 15011 24915 15017
rect 24857 14977 24869 15011
rect 24903 15008 24915 15011
rect 25041 15011 25099 15017
rect 25041 15008 25053 15011
rect 24903 14980 25053 15008
rect 24903 14977 24915 14980
rect 24857 14971 24915 14977
rect 25041 14977 25053 14980
rect 25087 14977 25099 15011
rect 25222 15008 25228 15020
rect 25183 14980 25228 15008
rect 25041 14971 25099 14977
rect 25222 14968 25228 14980
rect 25280 14968 25286 15020
rect 25961 15011 26019 15017
rect 25961 14977 25973 15011
rect 26007 14977 26019 15011
rect 25961 14971 26019 14977
rect 15019 14912 17448 14940
rect 18138 14900 18144 14952
rect 18196 14940 18202 14952
rect 18892 14940 18920 14968
rect 18196 14912 18920 14940
rect 20165 14943 20223 14949
rect 18196 14900 18202 14912
rect 20165 14909 20177 14943
rect 20211 14940 20223 14943
rect 20809 14943 20867 14949
rect 20809 14940 20821 14943
rect 20211 14912 20821 14940
rect 20211 14909 20223 14912
rect 20165 14903 20223 14909
rect 20809 14909 20821 14912
rect 20855 14909 20867 14943
rect 22186 14940 22192 14952
rect 20809 14903 20867 14909
rect 21376 14912 22192 14940
rect 13538 14872 13544 14884
rect 8864 14844 9996 14872
rect 3568 14776 6868 14804
rect 6917 14807 6975 14813
rect 3568 14764 3574 14776
rect 6917 14773 6929 14807
rect 6963 14804 6975 14807
rect 7190 14804 7196 14816
rect 6963 14776 7196 14804
rect 6963 14773 6975 14776
rect 6917 14767 6975 14773
rect 7190 14764 7196 14776
rect 7248 14804 7254 14816
rect 7374 14804 7380 14816
rect 7248 14776 7380 14804
rect 7248 14764 7254 14776
rect 7374 14764 7380 14776
rect 7432 14764 7438 14816
rect 7466 14764 7472 14816
rect 7524 14804 7530 14816
rect 9217 14807 9275 14813
rect 9217 14804 9229 14807
rect 7524 14776 9229 14804
rect 7524 14764 7530 14776
rect 9217 14773 9229 14776
rect 9263 14804 9275 14807
rect 9398 14804 9404 14816
rect 9263 14776 9404 14804
rect 9263 14773 9275 14776
rect 9217 14767 9275 14773
rect 9398 14764 9404 14776
rect 9456 14764 9462 14816
rect 9490 14764 9496 14816
rect 9548 14804 9554 14816
rect 9861 14807 9919 14813
rect 9861 14804 9873 14807
rect 9548 14776 9873 14804
rect 9548 14764 9554 14776
rect 9861 14773 9873 14776
rect 9907 14773 9919 14807
rect 9968 14804 9996 14844
rect 12811 14844 13544 14872
rect 12811 14804 12839 14844
rect 13538 14832 13544 14844
rect 13596 14832 13602 14884
rect 17862 14872 17868 14884
rect 14936 14844 17868 14872
rect 14936 14816 14964 14844
rect 17862 14832 17868 14844
rect 17920 14832 17926 14884
rect 18322 14872 18328 14884
rect 18283 14844 18328 14872
rect 18322 14832 18328 14844
rect 18380 14832 18386 14884
rect 20625 14875 20683 14881
rect 20625 14841 20637 14875
rect 20671 14872 20683 14875
rect 21376 14872 21404 14912
rect 22186 14900 22192 14912
rect 22244 14900 22250 14952
rect 22557 14943 22615 14949
rect 22557 14909 22569 14943
rect 22603 14940 22615 14943
rect 22922 14940 22928 14952
rect 22603 14912 22928 14940
rect 22603 14909 22615 14912
rect 22557 14903 22615 14909
rect 22922 14900 22928 14912
rect 22980 14900 22986 14952
rect 24486 14900 24492 14952
rect 24544 14940 24550 14952
rect 25976 14940 26004 14971
rect 26142 14968 26148 15020
rect 26200 15008 26206 15020
rect 26237 15011 26295 15017
rect 26237 15008 26249 15011
rect 26200 14980 26249 15008
rect 26200 14968 26206 14980
rect 26237 14977 26249 14980
rect 26283 14977 26295 15011
rect 26237 14971 26295 14977
rect 26421 15011 26479 15017
rect 26421 14977 26433 15011
rect 26467 15008 26479 15011
rect 26970 15008 26976 15020
rect 26467 14980 26976 15008
rect 26467 14977 26479 14980
rect 26421 14971 26479 14977
rect 26970 14968 26976 14980
rect 27028 14968 27034 15020
rect 27065 15011 27123 15017
rect 27065 14977 27077 15011
rect 27111 15008 27123 15011
rect 27246 15008 27252 15020
rect 27111 14980 27252 15008
rect 27111 14977 27123 14980
rect 27065 14971 27123 14977
rect 27246 14968 27252 14980
rect 27304 14968 27310 15020
rect 28368 15017 28396 15048
rect 28994 15036 29000 15048
rect 29052 15076 29058 15088
rect 29914 15076 29920 15088
rect 29052 15048 29920 15076
rect 29052 15036 29058 15048
rect 29914 15036 29920 15048
rect 29972 15036 29978 15088
rect 28626 15017 28632 15020
rect 28353 15011 28411 15017
rect 28353 14977 28365 15011
rect 28399 14977 28411 15011
rect 28353 14971 28411 14977
rect 28620 14971 28632 15017
rect 28684 15008 28690 15020
rect 28684 14980 28720 15008
rect 28626 14968 28632 14971
rect 28684 14968 28690 14980
rect 30742 14968 30748 15020
rect 30800 15008 30806 15020
rect 30837 15011 30895 15017
rect 30837 15008 30849 15011
rect 30800 14980 30849 15008
rect 30800 14968 30806 14980
rect 30837 14977 30849 14980
rect 30883 14977 30895 15011
rect 30837 14971 30895 14977
rect 31018 14968 31024 15020
rect 31076 15008 31082 15020
rect 31113 15011 31171 15017
rect 31113 15008 31125 15011
rect 31076 14980 31125 15008
rect 31076 14968 31082 14980
rect 31113 14977 31125 14980
rect 31159 14977 31171 15011
rect 31113 14971 31171 14977
rect 24544 14912 26004 14940
rect 24544 14900 24550 14912
rect 25240 14884 25268 14912
rect 26786 14900 26792 14952
rect 26844 14940 26850 14952
rect 27338 14940 27344 14952
rect 26844 14912 27344 14940
rect 26844 14900 26850 14912
rect 27338 14900 27344 14912
rect 27396 14900 27402 14952
rect 24857 14875 24915 14881
rect 24857 14872 24869 14875
rect 20671 14844 21404 14872
rect 24412 14844 24869 14872
rect 20671 14841 20683 14844
rect 20625 14835 20683 14841
rect 9968 14776 12839 14804
rect 13265 14807 13323 14813
rect 9861 14767 9919 14773
rect 13265 14773 13277 14807
rect 13311 14804 13323 14807
rect 14734 14804 14740 14816
rect 13311 14776 14740 14804
rect 13311 14773 13323 14776
rect 13265 14767 13323 14773
rect 14734 14764 14740 14776
rect 14792 14764 14798 14816
rect 14918 14764 14924 14816
rect 14976 14764 14982 14816
rect 15473 14807 15531 14813
rect 15473 14773 15485 14807
rect 15519 14804 15531 14807
rect 15654 14804 15660 14816
rect 15519 14776 15660 14804
rect 15519 14773 15531 14776
rect 15473 14767 15531 14773
rect 15654 14764 15660 14776
rect 15712 14764 15718 14816
rect 15746 14764 15752 14816
rect 15804 14804 15810 14816
rect 16022 14804 16028 14816
rect 15804 14776 16028 14804
rect 15804 14764 15810 14776
rect 16022 14764 16028 14776
rect 16080 14764 16086 14816
rect 16206 14764 16212 14816
rect 16264 14804 16270 14816
rect 17402 14804 17408 14816
rect 16264 14776 17408 14804
rect 16264 14764 16270 14776
rect 17402 14764 17408 14776
rect 17460 14764 17466 14816
rect 17678 14764 17684 14816
rect 17736 14804 17742 14816
rect 18417 14807 18475 14813
rect 18417 14804 18429 14807
rect 17736 14776 18429 14804
rect 17736 14764 17742 14776
rect 18417 14773 18429 14776
rect 18463 14773 18475 14807
rect 18417 14767 18475 14773
rect 19061 14807 19119 14813
rect 19061 14773 19073 14807
rect 19107 14804 19119 14807
rect 19886 14804 19892 14816
rect 19107 14776 19892 14804
rect 19107 14773 19119 14776
rect 19061 14767 19119 14773
rect 19886 14764 19892 14776
rect 19944 14764 19950 14816
rect 20714 14764 20720 14816
rect 20772 14804 20778 14816
rect 24412 14804 24440 14844
rect 24857 14841 24869 14844
rect 24903 14841 24915 14875
rect 24857 14835 24915 14841
rect 25222 14832 25228 14884
rect 25280 14832 25286 14884
rect 30374 14832 30380 14884
rect 30432 14872 30438 14884
rect 31021 14875 31079 14881
rect 31021 14872 31033 14875
rect 30432 14844 31033 14872
rect 30432 14832 30438 14844
rect 31021 14841 31033 14844
rect 31067 14841 31079 14875
rect 31021 14835 31079 14841
rect 20772 14776 24440 14804
rect 24489 14807 24547 14813
rect 20772 14764 20778 14776
rect 24489 14773 24501 14807
rect 24535 14804 24547 14807
rect 25038 14804 25044 14816
rect 24535 14776 25044 14804
rect 24535 14773 24547 14776
rect 24489 14767 24547 14773
rect 25038 14764 25044 14776
rect 25096 14764 25102 14816
rect 25777 14807 25835 14813
rect 25777 14773 25789 14807
rect 25823 14804 25835 14807
rect 27062 14804 27068 14816
rect 25823 14776 27068 14804
rect 25823 14773 25835 14776
rect 25777 14767 25835 14773
rect 27062 14764 27068 14776
rect 27120 14764 27126 14816
rect 27154 14764 27160 14816
rect 27212 14804 27218 14816
rect 27212 14776 27257 14804
rect 27212 14764 27218 14776
rect 1104 14714 32016 14736
rect 1104 14662 2136 14714
rect 2188 14662 12440 14714
rect 12492 14662 22744 14714
rect 22796 14662 32016 14714
rect 1104 14640 32016 14662
rect 2682 14560 2688 14612
rect 2740 14600 2746 14612
rect 3510 14600 3516 14612
rect 2740 14572 3516 14600
rect 2740 14560 2746 14572
rect 3510 14560 3516 14572
rect 3568 14560 3574 14612
rect 5442 14560 5448 14612
rect 5500 14600 5506 14612
rect 6822 14600 6828 14612
rect 5500 14572 6828 14600
rect 5500 14560 5506 14572
rect 6822 14560 6828 14572
rect 6880 14560 6886 14612
rect 8202 14560 8208 14612
rect 8260 14600 8266 14612
rect 8297 14603 8355 14609
rect 8297 14600 8309 14603
rect 8260 14572 8309 14600
rect 8260 14560 8266 14572
rect 8297 14569 8309 14572
rect 8343 14569 8355 14603
rect 9766 14600 9772 14612
rect 8297 14563 8355 14569
rect 8864 14572 9772 14600
rect 2406 14492 2412 14544
rect 2464 14532 2470 14544
rect 4062 14532 4068 14544
rect 2464 14504 4068 14532
rect 2464 14492 2470 14504
rect 4062 14492 4068 14504
rect 4120 14492 4126 14544
rect 4433 14467 4491 14473
rect 4433 14433 4445 14467
rect 4479 14464 4491 14467
rect 4614 14464 4620 14476
rect 4479 14436 4620 14464
rect 4479 14433 4491 14436
rect 4433 14427 4491 14433
rect 4614 14424 4620 14436
rect 4672 14424 4678 14476
rect 6086 14464 6092 14476
rect 5000 14436 6092 14464
rect 1394 14396 1400 14408
rect 1355 14368 1400 14396
rect 1394 14356 1400 14368
rect 1452 14356 1458 14408
rect 4154 14356 4160 14408
rect 4212 14396 4218 14408
rect 5000 14405 5028 14436
rect 6086 14424 6092 14436
rect 6144 14424 6150 14476
rect 6270 14464 6276 14476
rect 6231 14436 6276 14464
rect 6270 14424 6276 14436
rect 6328 14424 6334 14476
rect 8754 14464 8760 14476
rect 8050 14436 8760 14464
rect 8754 14424 8760 14436
rect 8812 14424 8818 14476
rect 4249 14399 4307 14405
rect 4249 14396 4261 14399
rect 4212 14368 4261 14396
rect 4212 14356 4218 14368
rect 4249 14365 4261 14368
rect 4295 14365 4307 14399
rect 4249 14359 4307 14365
rect 4985 14399 5043 14405
rect 4985 14365 4997 14399
rect 5031 14365 5043 14399
rect 5166 14396 5172 14408
rect 5127 14368 5172 14396
rect 4985 14359 5043 14365
rect 5166 14356 5172 14368
rect 5224 14356 5230 14408
rect 5350 14356 5356 14408
rect 5408 14396 5414 14408
rect 5997 14399 6055 14405
rect 5997 14396 6009 14399
rect 5408 14368 6009 14396
rect 5408 14356 5414 14368
rect 5997 14365 6009 14368
rect 6043 14365 6055 14399
rect 5997 14359 6055 14365
rect 7377 14399 7435 14405
rect 7377 14365 7389 14399
rect 7423 14396 7435 14399
rect 8864 14396 8892 14572
rect 9766 14560 9772 14572
rect 9824 14600 9830 14612
rect 10502 14600 10508 14612
rect 9824 14572 10508 14600
rect 9824 14560 9830 14572
rect 10502 14560 10508 14572
rect 10560 14560 10566 14612
rect 13998 14560 14004 14612
rect 14056 14600 14062 14612
rect 14093 14603 14151 14609
rect 14093 14600 14105 14603
rect 14056 14572 14105 14600
rect 14056 14560 14062 14572
rect 14093 14569 14105 14572
rect 14139 14569 14151 14603
rect 14093 14563 14151 14569
rect 14182 14560 14188 14612
rect 14240 14600 14246 14612
rect 15194 14600 15200 14612
rect 14240 14572 15200 14600
rect 14240 14560 14246 14572
rect 15194 14560 15200 14572
rect 15252 14560 15258 14612
rect 15289 14603 15347 14609
rect 15289 14569 15301 14603
rect 15335 14600 15347 14603
rect 23382 14600 23388 14612
rect 15335 14572 18368 14600
rect 23343 14572 23388 14600
rect 15335 14569 15347 14572
rect 15289 14563 15347 14569
rect 9677 14535 9735 14541
rect 9677 14501 9689 14535
rect 9723 14532 9735 14535
rect 9950 14532 9956 14544
rect 9723 14504 9956 14532
rect 9723 14501 9735 14504
rect 9677 14495 9735 14501
rect 9950 14492 9956 14504
rect 10008 14492 10014 14544
rect 13538 14532 13544 14544
rect 13451 14504 13544 14532
rect 13538 14492 13544 14504
rect 13596 14532 13602 14544
rect 17681 14535 17739 14541
rect 17681 14532 17693 14535
rect 13596 14504 17693 14532
rect 13596 14492 13602 14504
rect 17681 14501 17693 14504
rect 17727 14501 17739 14535
rect 17681 14495 17739 14501
rect 8938 14424 8944 14476
rect 8996 14464 9002 14476
rect 10229 14467 10287 14473
rect 10229 14464 10241 14467
rect 8996 14436 10241 14464
rect 8996 14424 9002 14436
rect 10229 14433 10241 14436
rect 10275 14433 10287 14467
rect 10229 14427 10287 14433
rect 13170 14424 13176 14476
rect 13228 14464 13234 14476
rect 13228 14436 14320 14464
rect 13228 14424 13234 14436
rect 7423 14368 8892 14396
rect 9493 14399 9551 14405
rect 7423 14365 7435 14368
rect 7377 14359 7435 14365
rect 9493 14365 9505 14399
rect 9539 14396 9551 14399
rect 9582 14396 9588 14408
rect 9539 14368 9588 14396
rect 9539 14365 9551 14368
rect 9493 14359 9551 14365
rect 9582 14356 9588 14368
rect 9640 14356 9646 14408
rect 9769 14399 9827 14405
rect 9769 14365 9781 14399
rect 9815 14396 9827 14399
rect 9861 14399 9919 14405
rect 9861 14396 9873 14399
rect 9815 14368 9873 14396
rect 9815 14365 9827 14368
rect 9769 14359 9827 14365
rect 9861 14365 9873 14368
rect 9907 14396 9919 14399
rect 11698 14396 11704 14408
rect 9907 14368 11704 14396
rect 9907 14365 9919 14368
rect 9861 14359 9919 14365
rect 11698 14356 11704 14368
rect 11756 14356 11762 14408
rect 11882 14356 11888 14408
rect 11940 14396 11946 14408
rect 12158 14396 12164 14408
rect 11940 14368 12164 14396
rect 11940 14356 11946 14368
rect 12158 14356 12164 14368
rect 12216 14396 12222 14408
rect 13814 14396 13820 14408
rect 12216 14368 13820 14396
rect 12216 14356 12222 14368
rect 13814 14356 13820 14368
rect 13872 14356 13878 14408
rect 14292 14405 14320 14436
rect 15470 14424 15476 14476
rect 15528 14464 15534 14476
rect 15528 14436 15884 14464
rect 15528 14424 15534 14436
rect 14277 14399 14335 14405
rect 14277 14365 14289 14399
rect 14323 14365 14335 14399
rect 14277 14359 14335 14365
rect 14553 14399 14611 14405
rect 14553 14365 14565 14399
rect 14599 14365 14611 14399
rect 14734 14396 14740 14408
rect 14695 14368 14740 14396
rect 14553 14359 14611 14365
rect 1664 14331 1722 14337
rect 1664 14297 1676 14331
rect 1710 14328 1722 14331
rect 2682 14328 2688 14340
rect 1710 14300 2688 14328
rect 1710 14297 1722 14300
rect 1664 14291 1722 14297
rect 2682 14288 2688 14300
rect 2740 14288 2746 14340
rect 5077 14331 5135 14337
rect 5077 14297 5089 14331
rect 5123 14328 5135 14331
rect 6914 14328 6920 14340
rect 5123 14300 6920 14328
rect 5123 14297 5135 14300
rect 5077 14291 5135 14297
rect 6914 14288 6920 14300
rect 6972 14288 6978 14340
rect 7285 14331 7343 14337
rect 7285 14297 7297 14331
rect 7331 14297 7343 14331
rect 7742 14328 7748 14340
rect 7703 14300 7748 14328
rect 7285 14291 7343 14297
rect 2774 14260 2780 14272
rect 2735 14232 2780 14260
rect 2774 14220 2780 14232
rect 2832 14220 2838 14272
rect 3510 14220 3516 14272
rect 3568 14260 3574 14272
rect 3789 14263 3847 14269
rect 3789 14260 3801 14263
rect 3568 14232 3801 14260
rect 3568 14220 3574 14232
rect 3789 14229 3801 14232
rect 3835 14229 3847 14263
rect 3789 14223 3847 14229
rect 4157 14263 4215 14269
rect 4157 14229 4169 14263
rect 4203 14260 4215 14263
rect 4338 14260 4344 14272
rect 4203 14232 4344 14260
rect 4203 14229 4215 14232
rect 4157 14223 4215 14229
rect 4338 14220 4344 14232
rect 4396 14260 4402 14272
rect 5442 14260 5448 14272
rect 4396 14232 5448 14260
rect 4396 14220 4402 14232
rect 5442 14220 5448 14232
rect 5500 14220 5506 14272
rect 5629 14263 5687 14269
rect 5629 14229 5641 14263
rect 5675 14260 5687 14263
rect 5718 14260 5724 14272
rect 5675 14232 5724 14260
rect 5675 14229 5687 14232
rect 5629 14223 5687 14229
rect 5718 14220 5724 14232
rect 5776 14220 5782 14272
rect 6089 14263 6147 14269
rect 6089 14229 6101 14263
rect 6135 14260 6147 14263
rect 6178 14260 6184 14272
rect 6135 14232 6184 14260
rect 6135 14229 6147 14232
rect 6089 14223 6147 14229
rect 6178 14220 6184 14232
rect 6236 14220 6242 14272
rect 6546 14220 6552 14272
rect 6604 14260 6610 14272
rect 7009 14263 7067 14269
rect 7009 14260 7021 14263
rect 6604 14232 7021 14260
rect 6604 14220 6610 14232
rect 7009 14229 7021 14232
rect 7055 14229 7067 14263
rect 7300 14260 7328 14291
rect 7742 14288 7748 14300
rect 7800 14288 7806 14340
rect 9309 14331 9367 14337
rect 9309 14297 9321 14331
rect 9355 14328 9367 14331
rect 10474 14331 10532 14337
rect 10474 14328 10486 14331
rect 9355 14300 10486 14328
rect 9355 14297 9367 14300
rect 9309 14291 9367 14297
rect 10474 14297 10486 14300
rect 10520 14297 10532 14331
rect 10474 14291 10532 14297
rect 11974 14288 11980 14340
rect 12032 14328 12038 14340
rect 12406 14331 12464 14337
rect 12406 14328 12418 14331
rect 12032 14300 12418 14328
rect 12032 14288 12038 14300
rect 12406 14297 12418 14300
rect 12452 14297 12464 14331
rect 12406 14291 12464 14297
rect 13446 14288 13452 14340
rect 13504 14328 13510 14340
rect 14568 14328 14596 14359
rect 14734 14356 14740 14368
rect 14792 14356 14798 14408
rect 15010 14356 15016 14408
rect 15068 14396 15074 14408
rect 15856 14405 15884 14436
rect 15930 14424 15936 14476
rect 15988 14464 15994 14476
rect 17310 14464 17316 14476
rect 15988 14436 17316 14464
rect 15988 14424 15994 14436
rect 17310 14424 17316 14436
rect 17368 14424 17374 14476
rect 18340 14464 18368 14572
rect 23382 14560 23388 14572
rect 23440 14560 23446 14612
rect 25958 14600 25964 14612
rect 25919 14572 25964 14600
rect 25958 14560 25964 14572
rect 26016 14560 26022 14612
rect 27430 14600 27436 14612
rect 27391 14572 27436 14600
rect 27430 14560 27436 14572
rect 27488 14560 27494 14612
rect 27614 14560 27620 14612
rect 27672 14600 27678 14612
rect 27709 14603 27767 14609
rect 27709 14600 27721 14603
rect 27672 14572 27721 14600
rect 27672 14560 27678 14572
rect 27709 14569 27721 14572
rect 27755 14569 27767 14603
rect 27709 14563 27767 14569
rect 28537 14603 28595 14609
rect 28537 14569 28549 14603
rect 28583 14600 28595 14603
rect 28626 14600 28632 14612
rect 28583 14572 28632 14600
rect 28583 14569 28595 14572
rect 28537 14563 28595 14569
rect 28626 14560 28632 14572
rect 28684 14560 28690 14612
rect 18690 14492 18696 14544
rect 18748 14532 18754 14544
rect 19521 14535 19579 14541
rect 19521 14532 19533 14535
rect 18748 14504 19533 14532
rect 18748 14492 18754 14504
rect 19521 14501 19533 14504
rect 19567 14532 19579 14535
rect 23290 14532 23296 14544
rect 19567 14504 23296 14532
rect 19567 14501 19579 14504
rect 19521 14495 19579 14501
rect 23290 14492 23296 14504
rect 23348 14492 23354 14544
rect 24397 14535 24455 14541
rect 24397 14532 24409 14535
rect 23584 14504 24409 14532
rect 18509 14467 18567 14473
rect 18509 14464 18521 14467
rect 18340 14436 18521 14464
rect 18509 14433 18521 14436
rect 18555 14433 18567 14467
rect 22830 14464 22836 14476
rect 18509 14427 18567 14433
rect 19260 14436 22836 14464
rect 15565 14399 15623 14405
rect 15565 14396 15577 14399
rect 15068 14368 15577 14396
rect 15068 14356 15074 14368
rect 15565 14365 15577 14368
rect 15611 14365 15623 14399
rect 15565 14359 15623 14365
rect 15841 14399 15899 14405
rect 15841 14365 15853 14399
rect 15887 14365 15899 14399
rect 15841 14359 15899 14365
rect 16025 14399 16083 14405
rect 16025 14365 16037 14399
rect 16071 14396 16083 14399
rect 16114 14396 16120 14408
rect 16071 14368 16120 14396
rect 16071 14365 16083 14368
rect 16025 14359 16083 14365
rect 16114 14356 16120 14368
rect 16172 14356 16178 14408
rect 16945 14399 17003 14405
rect 16945 14365 16957 14399
rect 16991 14365 17003 14399
rect 16945 14359 17003 14365
rect 13504 14300 14596 14328
rect 13504 14288 13510 14300
rect 15102 14288 15108 14340
rect 15160 14328 15166 14340
rect 16960 14328 16988 14359
rect 17034 14356 17040 14408
rect 17092 14396 17098 14408
rect 17221 14399 17279 14405
rect 17221 14396 17233 14399
rect 17092 14368 17233 14396
rect 17092 14356 17098 14368
rect 17221 14365 17233 14368
rect 17267 14365 17279 14399
rect 17221 14359 17279 14365
rect 17681 14399 17739 14405
rect 17681 14365 17693 14399
rect 17727 14396 17739 14399
rect 17926 14396 18092 14406
rect 18325 14399 18383 14405
rect 18325 14396 18337 14399
rect 17727 14378 18337 14396
rect 17727 14368 17954 14378
rect 18064 14368 18337 14378
rect 17727 14365 17739 14368
rect 17681 14359 17739 14365
rect 18325 14365 18337 14368
rect 18371 14365 18383 14399
rect 18325 14359 18383 14365
rect 18417 14399 18475 14405
rect 18417 14365 18429 14399
rect 18463 14396 18475 14399
rect 18463 14368 18644 14396
rect 18463 14365 18475 14368
rect 18417 14359 18475 14365
rect 15160 14300 16988 14328
rect 17236 14328 17264 14359
rect 18616 14328 18644 14368
rect 18690 14328 18696 14340
rect 17236 14300 18554 14328
rect 18616 14300 18696 14328
rect 15160 14288 15166 14300
rect 7926 14260 7932 14272
rect 7300 14232 7932 14260
rect 7009 14223 7067 14229
rect 7926 14220 7932 14232
rect 7984 14220 7990 14272
rect 8113 14263 8171 14269
rect 8113 14229 8125 14263
rect 8159 14260 8171 14263
rect 8202 14260 8208 14272
rect 8159 14232 8208 14260
rect 8159 14229 8171 14232
rect 8113 14223 8171 14229
rect 8202 14220 8208 14232
rect 8260 14220 8266 14272
rect 8294 14220 8300 14272
rect 8352 14260 8358 14272
rect 9398 14260 9404 14272
rect 8352 14232 9404 14260
rect 8352 14220 8358 14232
rect 9398 14220 9404 14232
rect 9456 14260 9462 14272
rect 9861 14263 9919 14269
rect 9861 14260 9873 14263
rect 9456 14232 9873 14260
rect 9456 14220 9462 14232
rect 9861 14229 9873 14232
rect 9907 14229 9919 14263
rect 11606 14260 11612 14272
rect 11567 14232 11612 14260
rect 9861 14223 9919 14229
rect 11606 14220 11612 14232
rect 11664 14220 11670 14272
rect 12986 14220 12992 14272
rect 13044 14260 13050 14272
rect 13722 14260 13728 14272
rect 13044 14232 13728 14260
rect 13044 14220 13050 14232
rect 13722 14220 13728 14232
rect 13780 14260 13786 14272
rect 15289 14263 15347 14269
rect 15289 14260 15301 14263
rect 13780 14232 15301 14260
rect 13780 14220 13786 14232
rect 15289 14229 15301 14232
rect 15335 14229 15347 14263
rect 15289 14223 15347 14229
rect 15381 14263 15439 14269
rect 15381 14229 15393 14263
rect 15427 14260 15439 14263
rect 15746 14260 15752 14272
rect 15427 14232 15752 14260
rect 15427 14229 15439 14232
rect 15381 14223 15439 14229
rect 15746 14220 15752 14232
rect 15804 14220 15810 14272
rect 17957 14263 18015 14269
rect 17957 14229 17969 14263
rect 18003 14260 18015 14263
rect 18230 14260 18236 14272
rect 18003 14232 18236 14260
rect 18003 14229 18015 14232
rect 17957 14223 18015 14229
rect 18230 14220 18236 14232
rect 18288 14220 18294 14272
rect 18526 14260 18554 14300
rect 18690 14288 18696 14300
rect 18748 14288 18754 14340
rect 19260 14260 19288 14436
rect 22830 14424 22836 14436
rect 22888 14424 22894 14476
rect 19337 14399 19395 14405
rect 19337 14365 19349 14399
rect 19383 14396 19395 14399
rect 19426 14396 19432 14408
rect 19383 14368 19432 14396
rect 19383 14365 19395 14368
rect 19337 14359 19395 14365
rect 19426 14356 19432 14368
rect 19484 14396 19490 14408
rect 20073 14399 20131 14405
rect 19484 14368 19932 14396
rect 19484 14356 19490 14368
rect 18526 14232 19288 14260
rect 19904 14260 19932 14368
rect 20073 14365 20085 14399
rect 20119 14396 20131 14399
rect 20622 14396 20628 14408
rect 20119 14368 20628 14396
rect 20119 14365 20131 14368
rect 20073 14359 20131 14365
rect 20622 14356 20628 14368
rect 20680 14356 20686 14408
rect 22370 14356 22376 14408
rect 22428 14396 22434 14408
rect 22465 14399 22523 14405
rect 22465 14396 22477 14399
rect 22428 14368 22477 14396
rect 22428 14356 22434 14368
rect 22465 14365 22477 14368
rect 22511 14365 22523 14399
rect 22465 14359 22523 14365
rect 22480 14328 22508 14359
rect 22554 14356 22560 14408
rect 22612 14396 22618 14408
rect 22741 14399 22799 14405
rect 22741 14396 22753 14399
rect 22612 14368 22753 14396
rect 22612 14356 22618 14368
rect 22741 14365 22753 14368
rect 22787 14365 22799 14399
rect 22922 14396 22928 14408
rect 22883 14368 22928 14396
rect 22741 14359 22799 14365
rect 22922 14356 22928 14368
rect 22980 14356 22986 14408
rect 23584 14405 23612 14504
rect 24397 14501 24409 14504
rect 24443 14501 24455 14535
rect 24946 14532 24952 14544
rect 24397 14495 24455 14501
rect 24872 14504 24952 14532
rect 23569 14399 23627 14405
rect 23569 14365 23581 14399
rect 23615 14365 23627 14399
rect 23569 14359 23627 14365
rect 23658 14356 23664 14408
rect 23716 14396 23722 14408
rect 23753 14399 23811 14405
rect 23753 14396 23765 14399
rect 23716 14368 23765 14396
rect 23716 14356 23722 14368
rect 23753 14365 23765 14368
rect 23799 14365 23811 14399
rect 23753 14359 23811 14365
rect 23845 14399 23903 14405
rect 23845 14365 23857 14399
rect 23891 14396 23903 14399
rect 24302 14396 24308 14408
rect 23891 14368 24308 14396
rect 23891 14365 23903 14368
rect 23845 14359 23903 14365
rect 24302 14356 24308 14368
rect 24360 14374 24366 14408
rect 24872 14405 24900 14504
rect 24946 14492 24952 14504
rect 25004 14492 25010 14544
rect 25038 14492 25044 14544
rect 25096 14532 25102 14544
rect 26234 14532 26240 14544
rect 25096 14504 25176 14532
rect 25096 14492 25102 14504
rect 24581 14399 24639 14405
rect 24360 14356 24440 14374
rect 24581 14365 24593 14399
rect 24627 14365 24639 14399
rect 24872 14399 24948 14405
rect 24872 14368 24902 14399
rect 24581 14359 24639 14365
rect 24890 14365 24902 14368
rect 24936 14365 24948 14399
rect 24890 14359 24948 14365
rect 25053 14399 25111 14405
rect 25053 14365 25065 14399
rect 25099 14396 25111 14399
rect 25148 14396 25176 14504
rect 25792 14504 26240 14532
rect 25792 14464 25820 14504
rect 26234 14492 26240 14504
rect 26292 14492 26298 14544
rect 26326 14492 26332 14544
rect 26384 14532 26390 14544
rect 29730 14532 29736 14544
rect 26384 14504 29736 14532
rect 26384 14492 26390 14504
rect 29730 14492 29736 14504
rect 29788 14492 29794 14544
rect 25700 14436 25820 14464
rect 25700 14405 25728 14436
rect 25958 14424 25964 14476
rect 26016 14464 26022 14476
rect 29825 14467 29883 14473
rect 29825 14464 29837 14467
rect 26016 14436 29837 14464
rect 26016 14424 26022 14436
rect 29825 14433 29837 14436
rect 29871 14433 29883 14467
rect 29825 14427 29883 14433
rect 25099 14368 25176 14396
rect 25593 14399 25651 14405
rect 25099 14365 25111 14368
rect 25053 14359 25111 14365
rect 25593 14365 25605 14399
rect 25639 14365 25651 14399
rect 25593 14359 25651 14365
rect 25685 14399 25743 14405
rect 25685 14365 25697 14399
rect 25731 14365 25743 14399
rect 25685 14359 25743 14365
rect 25777 14399 25835 14405
rect 25777 14365 25789 14399
rect 25823 14365 25835 14399
rect 25777 14359 25835 14365
rect 24320 14346 24440 14356
rect 23382 14328 23388 14340
rect 22480 14300 23388 14328
rect 23382 14288 23388 14300
rect 23440 14288 23446 14340
rect 21174 14260 21180 14272
rect 19904 14232 21180 14260
rect 21174 14220 21180 14232
rect 21232 14220 21238 14272
rect 21358 14260 21364 14272
rect 21319 14232 21364 14260
rect 21358 14220 21364 14232
rect 21416 14220 21422 14272
rect 21818 14220 21824 14272
rect 21876 14260 21882 14272
rect 22281 14263 22339 14269
rect 22281 14260 22293 14263
rect 21876 14232 22293 14260
rect 21876 14220 21882 14232
rect 22281 14229 22293 14232
rect 22327 14229 22339 14263
rect 22281 14223 22339 14229
rect 23290 14220 23296 14272
rect 23348 14260 23354 14272
rect 24026 14260 24032 14272
rect 23348 14232 24032 14260
rect 23348 14220 23354 14232
rect 24026 14220 24032 14232
rect 24084 14220 24090 14272
rect 24412 14260 24440 14346
rect 24486 14288 24492 14340
rect 24544 14328 24550 14340
rect 24596 14328 24624 14359
rect 25608 14328 25636 14359
rect 24544 14300 24624 14328
rect 24657 14300 25636 14328
rect 24544 14288 24550 14300
rect 24657 14260 24685 14300
rect 24412 14232 24685 14260
rect 24854 14220 24860 14272
rect 24912 14260 24918 14272
rect 25792 14260 25820 14359
rect 26234 14356 26240 14408
rect 26292 14396 26298 14408
rect 27154 14396 27160 14408
rect 26292 14368 27160 14396
rect 26292 14356 26298 14368
rect 27154 14356 27160 14368
rect 27212 14356 27218 14408
rect 27246 14356 27252 14408
rect 27304 14396 27310 14408
rect 27433 14399 27491 14405
rect 27433 14396 27445 14399
rect 27304 14368 27445 14396
rect 27304 14356 27310 14368
rect 27433 14365 27445 14368
rect 27479 14365 27491 14399
rect 28718 14396 28724 14408
rect 28679 14368 28724 14396
rect 27433 14359 27491 14365
rect 28718 14356 28724 14368
rect 28776 14356 28782 14408
rect 28905 14399 28963 14405
rect 28905 14365 28917 14399
rect 28951 14365 28963 14399
rect 28905 14359 28963 14365
rect 28997 14399 29055 14405
rect 28997 14365 29009 14399
rect 29043 14396 29055 14399
rect 29178 14396 29184 14408
rect 29043 14368 29184 14396
rect 29043 14365 29055 14368
rect 28997 14359 29055 14365
rect 26513 14331 26571 14337
rect 26513 14297 26525 14331
rect 26559 14297 26571 14331
rect 26513 14291 26571 14297
rect 26697 14331 26755 14337
rect 26697 14297 26709 14331
rect 26743 14328 26755 14331
rect 28920 14328 28948 14359
rect 29178 14356 29184 14368
rect 29236 14356 29242 14408
rect 29454 14356 29460 14408
rect 29512 14396 29518 14408
rect 30081 14399 30139 14405
rect 30081 14396 30093 14399
rect 29512 14368 30093 14396
rect 29512 14356 29518 14368
rect 30081 14365 30093 14368
rect 30127 14365 30139 14399
rect 30081 14359 30139 14365
rect 29914 14328 29920 14340
rect 26743 14300 29920 14328
rect 26743 14297 26755 14300
rect 26697 14291 26755 14297
rect 24912 14232 25820 14260
rect 26528 14260 26556 14291
rect 29914 14288 29920 14300
rect 29972 14288 29978 14340
rect 29270 14260 29276 14272
rect 26528 14232 29276 14260
rect 24912 14220 24918 14232
rect 29270 14220 29276 14232
rect 29328 14220 29334 14272
rect 29638 14220 29644 14272
rect 29696 14260 29702 14272
rect 31205 14263 31263 14269
rect 31205 14260 31217 14263
rect 29696 14232 31217 14260
rect 29696 14220 29702 14232
rect 31205 14229 31217 14232
rect 31251 14229 31263 14263
rect 31205 14223 31263 14229
rect 1104 14170 32016 14192
rect 1104 14118 7288 14170
rect 7340 14118 17592 14170
rect 17644 14118 27896 14170
rect 27948 14118 32016 14170
rect 1104 14096 32016 14118
rect 1854 14016 1860 14068
rect 1912 14056 1918 14068
rect 2777 14059 2835 14065
rect 2777 14056 2789 14059
rect 1912 14028 2789 14056
rect 1912 14016 1918 14028
rect 2777 14025 2789 14028
rect 2823 14025 2835 14059
rect 3881 14059 3939 14065
rect 3881 14056 3893 14059
rect 2777 14019 2835 14025
rect 2945 14028 3893 14056
rect 2133 13991 2191 13997
rect 2133 13957 2145 13991
rect 2179 13988 2191 13991
rect 2945 13988 2973 14028
rect 3881 14025 3893 14028
rect 3927 14025 3939 14059
rect 3881 14019 3939 14025
rect 4065 14059 4123 14065
rect 4065 14025 4077 14059
rect 4111 14056 4123 14059
rect 4111 14028 7420 14056
rect 4111 14025 4123 14028
rect 4065 14019 4123 14025
rect 3050 13988 3056 14000
rect 2179 13960 2973 13988
rect 3011 13960 3056 13988
rect 2179 13957 2191 13960
rect 2133 13951 2191 13957
rect 3050 13948 3056 13960
rect 3108 13948 3114 14000
rect 3142 13948 3148 14000
rect 3200 13988 3206 14000
rect 3510 13988 3516 14000
rect 3200 13960 3245 13988
rect 3471 13960 3516 13988
rect 3200 13948 3206 13960
rect 3510 13948 3516 13960
rect 3568 13948 3574 14000
rect 4246 13948 4252 14000
rect 4304 13988 4310 14000
rect 5534 13988 5540 14000
rect 4304 13960 5540 13988
rect 4304 13948 4310 13960
rect 5534 13948 5540 13960
rect 5592 13948 5598 14000
rect 6178 13948 6184 14000
rect 6236 13988 6242 14000
rect 7009 13991 7067 13997
rect 7009 13988 7021 13991
rect 6236 13960 7021 13988
rect 6236 13948 6242 13960
rect 7009 13957 7021 13960
rect 7055 13957 7067 13991
rect 7009 13951 7067 13957
rect 1302 13880 1308 13932
rect 1360 13920 1366 13932
rect 1949 13923 2007 13929
rect 1949 13920 1961 13923
rect 1360 13892 1961 13920
rect 1360 13880 1366 13892
rect 1949 13889 1961 13892
rect 1995 13889 2007 13923
rect 1949 13883 2007 13889
rect 3970 13880 3976 13932
rect 4028 13920 4034 13932
rect 4893 13923 4951 13929
rect 4893 13920 4905 13923
rect 4028 13892 4905 13920
rect 4028 13880 4034 13892
rect 4893 13889 4905 13892
rect 4939 13889 4951 13923
rect 4893 13883 4951 13889
rect 5258 13880 5264 13932
rect 5316 13920 5322 13932
rect 6917 13923 6975 13929
rect 6917 13920 6929 13923
rect 5316 13892 6929 13920
rect 5316 13880 5322 13892
rect 6917 13889 6929 13892
rect 6963 13889 6975 13923
rect 7392 13920 7420 14028
rect 7926 14016 7932 14068
rect 7984 14056 7990 14068
rect 8205 14059 8263 14065
rect 8205 14056 8217 14059
rect 7984 14028 8217 14056
rect 7984 14016 7990 14028
rect 8205 14025 8217 14028
rect 8251 14025 8263 14059
rect 8941 14059 8999 14065
rect 8941 14056 8953 14059
rect 8205 14019 8263 14025
rect 8588 14028 8953 14056
rect 7650 13948 7656 14000
rect 7708 13988 7714 14000
rect 8588 13988 8616 14028
rect 8941 14025 8953 14028
rect 8987 14025 8999 14059
rect 8941 14019 8999 14025
rect 9582 14016 9588 14068
rect 9640 14056 9646 14068
rect 10321 14059 10379 14065
rect 10321 14056 10333 14059
rect 9640 14028 10333 14056
rect 9640 14016 9646 14028
rect 10321 14025 10333 14028
rect 10367 14025 10379 14059
rect 10321 14019 10379 14025
rect 10502 14016 10508 14068
rect 10560 14056 10566 14068
rect 12618 14056 12624 14068
rect 10560 14028 12624 14056
rect 10560 14016 10566 14028
rect 12618 14016 12624 14028
rect 12676 14056 12682 14068
rect 14642 14056 14648 14068
rect 12676 14028 13124 14056
rect 14603 14028 14648 14056
rect 12676 14016 12682 14028
rect 12986 13988 12992 14000
rect 7708 13960 8616 13988
rect 8772 13960 12992 13988
rect 7708 13948 7714 13960
rect 8386 13920 8392 13932
rect 7392 13892 8392 13920
rect 6917 13883 6975 13889
rect 8386 13880 8392 13892
rect 8444 13880 8450 13932
rect 8665 13923 8723 13929
rect 8665 13889 8677 13923
rect 8711 13920 8723 13923
rect 8772 13920 8800 13960
rect 12986 13948 12992 13960
rect 13044 13948 13050 14000
rect 8711 13892 8800 13920
rect 8849 13923 8907 13929
rect 8711 13889 8723 13892
rect 8665 13883 8723 13889
rect 8849 13889 8861 13923
rect 8895 13920 8907 13923
rect 8941 13923 8999 13929
rect 8941 13920 8953 13923
rect 8895 13892 8953 13920
rect 8895 13889 8907 13892
rect 8849 13883 8907 13889
rect 8941 13889 8953 13892
rect 8987 13920 8999 13923
rect 9122 13920 9128 13932
rect 8987 13892 9128 13920
rect 8987 13889 8999 13892
rect 8941 13883 8999 13889
rect 9122 13880 9128 13892
rect 9180 13880 9186 13932
rect 9490 13920 9496 13932
rect 9451 13892 9496 13920
rect 9490 13880 9496 13892
rect 9548 13880 9554 13932
rect 9677 13923 9735 13929
rect 9677 13889 9689 13923
rect 9723 13920 9735 13923
rect 9950 13920 9956 13932
rect 9723 13892 9956 13920
rect 9723 13889 9735 13892
rect 9677 13883 9735 13889
rect 9950 13880 9956 13892
rect 10008 13880 10014 13932
rect 10042 13880 10048 13932
rect 10100 13920 10106 13932
rect 10226 13920 10232 13932
rect 10100 13892 10232 13920
rect 10100 13880 10106 13892
rect 10226 13880 10232 13892
rect 10284 13920 10290 13932
rect 10502 13920 10508 13932
rect 10284 13892 10508 13920
rect 10284 13880 10290 13892
rect 10502 13880 10508 13892
rect 10560 13880 10566 13932
rect 10781 13923 10839 13929
rect 10781 13889 10793 13923
rect 10827 13920 10839 13923
rect 10870 13920 10876 13932
rect 10827 13892 10876 13920
rect 10827 13889 10839 13892
rect 10781 13883 10839 13889
rect 10870 13880 10876 13892
rect 10928 13880 10934 13932
rect 10965 13923 11023 13929
rect 10965 13889 10977 13923
rect 11011 13920 11023 13923
rect 11606 13920 11612 13932
rect 11011 13892 11612 13920
rect 11011 13889 11023 13892
rect 10965 13883 11023 13889
rect 2780 13864 2832 13870
rect 1765 13855 1823 13861
rect 1765 13821 1777 13855
rect 1811 13852 1823 13855
rect 2314 13852 2320 13864
rect 1811 13824 2320 13852
rect 1811 13821 1823 13824
rect 1765 13815 1823 13821
rect 2314 13812 2320 13824
rect 2372 13812 2378 13864
rect 4614 13852 4620 13864
rect 4575 13824 4620 13852
rect 4614 13812 4620 13824
rect 4672 13812 4678 13864
rect 5442 13812 5448 13864
rect 5500 13852 5506 13864
rect 7193 13855 7251 13861
rect 5500 13824 7144 13852
rect 5500 13812 5506 13824
rect 2780 13806 2832 13812
rect 6546 13784 6552 13796
rect 6507 13756 6552 13784
rect 6546 13744 6552 13756
rect 6604 13744 6610 13796
rect 7116 13784 7144 13824
rect 7193 13821 7205 13855
rect 7239 13852 7251 13855
rect 7745 13855 7803 13861
rect 7745 13852 7757 13855
rect 7239 13824 7757 13852
rect 7239 13821 7251 13824
rect 7193 13815 7251 13821
rect 7745 13821 7757 13824
rect 7791 13852 7803 13855
rect 8294 13852 8300 13864
rect 7791 13824 8300 13852
rect 7791 13821 7803 13824
rect 7745 13815 7803 13821
rect 8294 13812 8300 13824
rect 8352 13812 8358 13864
rect 8754 13812 8760 13864
rect 8812 13852 8818 13864
rect 9769 13855 9827 13861
rect 9769 13852 9781 13855
rect 8812 13824 9781 13852
rect 8812 13812 8818 13824
rect 9769 13821 9781 13824
rect 9815 13852 9827 13855
rect 10980 13852 11008 13883
rect 11606 13880 11612 13892
rect 11664 13880 11670 13932
rect 11974 13920 11980 13932
rect 11935 13892 11980 13920
rect 11974 13880 11980 13892
rect 12032 13880 12038 13932
rect 13096 13929 13124 14028
rect 14642 14016 14648 14028
rect 14700 14016 14706 14068
rect 14734 14016 14740 14068
rect 14792 14056 14798 14068
rect 16206 14056 16212 14068
rect 14792 14028 16212 14056
rect 14792 14016 14798 14028
rect 16206 14016 16212 14028
rect 16264 14016 16270 14068
rect 16666 14056 16672 14068
rect 16627 14028 16672 14056
rect 16666 14016 16672 14028
rect 16724 14016 16730 14068
rect 19242 14056 19248 14068
rect 16776 14028 17172 14056
rect 14093 13991 14151 13997
rect 14093 13957 14105 13991
rect 14139 13988 14151 13991
rect 15289 13991 15347 13997
rect 15289 13988 15301 13991
rect 14139 13960 15301 13988
rect 14139 13957 14151 13960
rect 14093 13951 14151 13957
rect 15289 13957 15301 13960
rect 15335 13957 15347 13991
rect 16776 13988 16804 14028
rect 17037 13991 17095 13997
rect 17037 13988 17049 13991
rect 15289 13951 15347 13957
rect 15488 13960 16804 13988
rect 16868 13960 17049 13988
rect 12161 13923 12219 13929
rect 12161 13889 12173 13923
rect 12207 13920 12219 13923
rect 12897 13923 12955 13929
rect 12897 13920 12909 13923
rect 12207 13892 12909 13920
rect 12207 13889 12219 13892
rect 12161 13883 12219 13889
rect 12897 13889 12909 13892
rect 12943 13889 12955 13923
rect 12897 13883 12955 13889
rect 13081 13923 13139 13929
rect 13081 13889 13093 13923
rect 13127 13920 13139 13923
rect 13170 13920 13176 13932
rect 13127 13892 13176 13920
rect 13127 13889 13139 13892
rect 13081 13883 13139 13889
rect 13170 13880 13176 13892
rect 13228 13880 13234 13932
rect 13357 13923 13415 13929
rect 13357 13889 13369 13923
rect 13403 13920 13415 13923
rect 13446 13920 13452 13932
rect 13403 13892 13452 13920
rect 13403 13889 13415 13892
rect 13357 13883 13415 13889
rect 13446 13880 13452 13892
rect 13504 13880 13510 13932
rect 13538 13880 13544 13932
rect 13596 13920 13602 13932
rect 14001 13923 14059 13929
rect 13596 13892 13641 13920
rect 13596 13880 13602 13892
rect 14001 13889 14013 13923
rect 14047 13889 14059 13923
rect 14001 13883 14059 13889
rect 14185 13923 14243 13929
rect 14185 13889 14197 13923
rect 14231 13920 14243 13923
rect 14277 13923 14335 13929
rect 14277 13920 14289 13923
rect 14231 13892 14289 13920
rect 14231 13889 14243 13892
rect 14185 13883 14243 13889
rect 14277 13889 14289 13892
rect 14323 13920 14335 13923
rect 14642 13920 14648 13932
rect 14323 13892 14648 13920
rect 14323 13889 14335 13892
rect 14277 13883 14335 13889
rect 12342 13852 12348 13864
rect 9815 13824 11008 13852
rect 12303 13824 12348 13852
rect 9815 13821 9827 13824
rect 9769 13815 9827 13821
rect 12342 13812 12348 13824
rect 12400 13812 12406 13864
rect 12437 13855 12495 13861
rect 12437 13821 12449 13855
rect 12483 13852 12495 13855
rect 13906 13852 13912 13864
rect 12483 13824 13912 13852
rect 12483 13821 12495 13824
rect 12437 13815 12495 13821
rect 13906 13812 13912 13824
rect 13964 13812 13970 13864
rect 14016 13852 14044 13883
rect 14642 13880 14648 13892
rect 14700 13880 14706 13932
rect 14826 13920 14832 13932
rect 14787 13892 14832 13920
rect 14826 13880 14832 13892
rect 14884 13880 14890 13932
rect 15105 13923 15163 13929
rect 15105 13889 15117 13923
rect 15151 13920 15163 13923
rect 15378 13920 15384 13932
rect 15151 13892 15384 13920
rect 15151 13889 15163 13892
rect 15105 13883 15163 13889
rect 15378 13880 15384 13892
rect 15436 13880 15442 13932
rect 15488 13852 15516 13960
rect 15749 13923 15807 13929
rect 15749 13889 15761 13923
rect 15795 13920 15807 13923
rect 15838 13920 15844 13932
rect 15795 13892 15844 13920
rect 15795 13889 15807 13892
rect 15749 13883 15807 13889
rect 15838 13880 15844 13892
rect 15896 13880 15902 13932
rect 15930 13880 15936 13932
rect 15988 13920 15994 13932
rect 16482 13920 16488 13932
rect 15988 13892 16488 13920
rect 15988 13880 15994 13892
rect 16482 13880 16488 13892
rect 16540 13880 16546 13932
rect 16868 13920 16896 13960
rect 17037 13957 17049 13960
rect 17083 13957 17095 13991
rect 17144 13988 17172 14028
rect 17236 14028 19248 14056
rect 17236 13988 17264 14028
rect 19242 14016 19248 14028
rect 19300 14016 19306 14068
rect 19978 14016 19984 14068
rect 20036 14016 20042 14068
rect 20990 14016 20996 14068
rect 21048 14056 21054 14068
rect 21177 14059 21235 14065
rect 21177 14056 21189 14059
rect 21048 14028 21189 14056
rect 21048 14016 21054 14028
rect 21177 14025 21189 14028
rect 21223 14025 21235 14059
rect 21177 14019 21235 14025
rect 21726 14016 21732 14068
rect 21784 14056 21790 14068
rect 21784 14028 22094 14056
rect 21784 14016 21790 14028
rect 18138 13988 18144 14000
rect 17144 13960 17264 13988
rect 17972 13960 18144 13988
rect 17037 13951 17095 13957
rect 16776 13892 16896 13920
rect 16776 13864 16804 13892
rect 16942 13880 16948 13932
rect 17000 13920 17006 13932
rect 17972 13929 18000 13960
rect 18138 13948 18144 13960
rect 18196 13988 18202 14000
rect 19996 13988 20024 14016
rect 21358 13988 21364 14000
rect 18196 13960 21364 13988
rect 18196 13948 18202 13960
rect 19812 13929 19840 13960
rect 21358 13948 21364 13960
rect 21416 13948 21422 14000
rect 22066 13997 22094 14028
rect 22922 14016 22928 14068
rect 22980 14056 22986 14068
rect 23201 14059 23259 14065
rect 23201 14056 23213 14059
rect 22980 14028 23213 14056
rect 22980 14016 22986 14028
rect 23201 14025 23213 14028
rect 23247 14056 23259 14059
rect 24670 14056 24676 14068
rect 23247 14028 24676 14056
rect 23247 14025 23259 14028
rect 23201 14019 23259 14025
rect 24670 14016 24676 14028
rect 24728 14016 24734 14068
rect 24854 14016 24860 14068
rect 24912 14056 24918 14068
rect 25130 14056 25136 14068
rect 24912 14028 25136 14056
rect 24912 14016 24918 14028
rect 25130 14016 25136 14028
rect 25188 14016 25194 14068
rect 25958 14056 25964 14068
rect 25516 14028 25964 14056
rect 22066 13991 22124 13997
rect 22066 13957 22078 13991
rect 22112 13957 22124 13991
rect 22066 13951 22124 13957
rect 23937 13991 23995 13997
rect 23937 13957 23949 13991
rect 23983 13988 23995 13991
rect 25516 13988 25544 14028
rect 25958 14016 25964 14028
rect 26016 14016 26022 14068
rect 26237 14059 26295 14065
rect 26237 14025 26249 14059
rect 26283 14056 26295 14059
rect 28813 14059 28871 14065
rect 26283 14028 28672 14056
rect 26283 14025 26295 14028
rect 26237 14019 26295 14025
rect 26142 13988 26148 14000
rect 23983 13960 25544 13988
rect 25608 13960 26148 13988
rect 23983 13957 23995 13960
rect 23937 13951 23995 13957
rect 17957 13923 18015 13929
rect 17000 13892 17448 13920
rect 17000 13880 17006 13892
rect 14016 13824 15516 13852
rect 15562 13812 15568 13864
rect 15620 13852 15626 13864
rect 16025 13855 16083 13861
rect 16025 13852 16037 13855
rect 15620 13824 16037 13852
rect 15620 13812 15626 13824
rect 16025 13821 16037 13824
rect 16071 13852 16083 13855
rect 16206 13852 16212 13864
rect 16071 13824 16212 13852
rect 16071 13821 16083 13824
rect 16025 13815 16083 13821
rect 16206 13812 16212 13824
rect 16264 13812 16270 13864
rect 16758 13812 16764 13864
rect 16816 13812 16822 13864
rect 16850 13812 16856 13864
rect 16908 13852 16914 13864
rect 17129 13855 17187 13861
rect 17129 13852 17141 13855
rect 16908 13824 17141 13852
rect 16908 13812 16914 13824
rect 17129 13821 17141 13824
rect 17175 13821 17187 13855
rect 17129 13815 17187 13821
rect 17221 13855 17279 13861
rect 17221 13821 17233 13855
rect 17267 13821 17279 13855
rect 17420 13852 17448 13892
rect 17957 13889 17969 13923
rect 18003 13889 18015 13923
rect 18224 13923 18282 13929
rect 18224 13920 18236 13923
rect 17957 13883 18015 13889
rect 18064 13892 18236 13920
rect 18064 13852 18092 13892
rect 18224 13889 18236 13892
rect 18270 13889 18282 13923
rect 18224 13883 18282 13889
rect 19797 13923 19855 13929
rect 19797 13889 19809 13923
rect 19843 13889 19855 13923
rect 19797 13883 19855 13889
rect 19886 13880 19892 13932
rect 19944 13920 19950 13932
rect 20053 13923 20111 13929
rect 20053 13920 20065 13923
rect 19944 13892 20065 13920
rect 19944 13880 19950 13892
rect 20053 13889 20065 13892
rect 20099 13889 20111 13923
rect 20053 13883 20111 13889
rect 21174 13880 21180 13932
rect 21232 13920 21238 13932
rect 22922 13920 22928 13932
rect 21232 13892 22928 13920
rect 21232 13880 21238 13892
rect 22922 13880 22928 13892
rect 22980 13880 22986 13932
rect 24397 13923 24455 13929
rect 24397 13889 24409 13923
rect 24443 13920 24455 13923
rect 25133 13923 25191 13929
rect 25133 13920 25145 13923
rect 24443 13892 25145 13920
rect 24443 13889 24455 13892
rect 24397 13883 24455 13889
rect 25133 13889 25145 13892
rect 25179 13889 25191 13923
rect 25133 13883 25191 13889
rect 25222 13880 25228 13932
rect 25280 13920 25286 13932
rect 25317 13923 25375 13929
rect 25317 13920 25329 13923
rect 25280 13892 25329 13920
rect 25280 13880 25286 13892
rect 25317 13889 25329 13892
rect 25363 13889 25375 13923
rect 25317 13883 25375 13889
rect 25498 13880 25504 13932
rect 25556 13920 25562 13932
rect 25608 13929 25636 13960
rect 26142 13948 26148 13960
rect 26200 13948 26206 14000
rect 28644 13997 28672 14028
rect 28813 14025 28825 14059
rect 28859 14056 28871 14059
rect 29086 14056 29092 14068
rect 28859 14028 29092 14056
rect 28859 14025 28871 14028
rect 28813 14019 28871 14025
rect 29086 14016 29092 14028
rect 29144 14016 29150 14068
rect 29641 14059 29699 14065
rect 29641 14025 29653 14059
rect 29687 14056 29699 14059
rect 30926 14056 30932 14068
rect 29687 14028 30932 14056
rect 29687 14025 29699 14028
rect 29641 14019 29699 14025
rect 30926 14016 30932 14028
rect 30984 14016 30990 14068
rect 28718 13997 28724 14000
rect 28445 13991 28503 13997
rect 26436 13960 28396 13988
rect 25593 13923 25651 13929
rect 25593 13920 25605 13923
rect 25556 13892 25605 13920
rect 25556 13880 25562 13892
rect 25593 13889 25605 13892
rect 25639 13889 25651 13923
rect 25774 13920 25780 13932
rect 25735 13892 25780 13920
rect 25593 13883 25651 13889
rect 25774 13880 25780 13892
rect 25832 13880 25838 13932
rect 26436 13929 26464 13960
rect 26421 13923 26479 13929
rect 26421 13889 26433 13923
rect 26467 13889 26479 13923
rect 26421 13883 26479 13889
rect 27062 13880 27068 13932
rect 27120 13920 27126 13932
rect 27157 13923 27215 13929
rect 27157 13920 27169 13923
rect 27120 13892 27169 13920
rect 27120 13880 27126 13892
rect 27157 13889 27169 13892
rect 27203 13889 27215 13923
rect 27157 13883 27215 13889
rect 27433 13923 27491 13929
rect 27433 13889 27445 13923
rect 27479 13920 27491 13923
rect 27522 13920 27528 13932
rect 27479 13892 27528 13920
rect 27479 13889 27491 13892
rect 27433 13883 27491 13889
rect 27522 13880 27528 13892
rect 27580 13880 27586 13932
rect 17420 13824 18092 13852
rect 17221 13815 17279 13821
rect 7650 13784 7656 13796
rect 7116 13756 7656 13784
rect 7650 13744 7656 13756
rect 7708 13744 7714 13796
rect 8018 13784 8024 13796
rect 7979 13756 8024 13784
rect 8018 13744 8024 13756
rect 8076 13744 8082 13796
rect 9306 13784 9312 13796
rect 8266 13756 8800 13784
rect 9267 13756 9312 13784
rect 4338 13676 4344 13728
rect 4396 13716 4402 13728
rect 8266 13716 8294 13756
rect 8662 13716 8668 13728
rect 4396 13688 8294 13716
rect 8623 13688 8668 13716
rect 4396 13676 4402 13688
rect 8662 13676 8668 13688
rect 8720 13676 8726 13728
rect 8772 13716 8800 13756
rect 9306 13744 9312 13756
rect 9364 13744 9370 13796
rect 10980 13756 15700 13784
rect 10980 13716 11008 13756
rect 8772 13688 11008 13716
rect 11054 13676 11060 13728
rect 11112 13716 11118 13728
rect 11514 13716 11520 13728
rect 11112 13688 11520 13716
rect 11112 13676 11118 13688
rect 11514 13676 11520 13688
rect 11572 13676 11578 13728
rect 11698 13676 11704 13728
rect 11756 13716 11762 13728
rect 12986 13716 12992 13728
rect 11756 13688 12992 13716
rect 11756 13676 11762 13688
rect 12986 13676 12992 13688
rect 13044 13676 13050 13728
rect 13538 13676 13544 13728
rect 13596 13716 13602 13728
rect 14277 13719 14335 13725
rect 14277 13716 14289 13719
rect 13596 13688 14289 13716
rect 13596 13676 13602 13688
rect 14277 13685 14289 13688
rect 14323 13685 14335 13719
rect 15010 13716 15016 13728
rect 14971 13688 15016 13716
rect 14277 13679 14335 13685
rect 15010 13676 15016 13688
rect 15068 13676 15074 13728
rect 15289 13719 15347 13725
rect 15289 13685 15301 13719
rect 15335 13716 15347 13719
rect 15378 13716 15384 13728
rect 15335 13688 15384 13716
rect 15335 13685 15347 13688
rect 15289 13679 15347 13685
rect 15378 13676 15384 13688
rect 15436 13676 15442 13728
rect 15562 13716 15568 13728
rect 15523 13688 15568 13716
rect 15562 13676 15568 13688
rect 15620 13676 15626 13728
rect 15672 13716 15700 13756
rect 16114 13744 16120 13796
rect 16172 13784 16178 13796
rect 17236 13784 17264 13815
rect 21358 13812 21364 13864
rect 21416 13852 21422 13864
rect 21821 13855 21879 13861
rect 21821 13852 21833 13855
rect 21416 13824 21833 13852
rect 21416 13812 21422 13824
rect 21821 13821 21833 13824
rect 21867 13821 21879 13855
rect 21821 13815 21879 13821
rect 23750 13812 23756 13864
rect 23808 13852 23814 13864
rect 24581 13855 24639 13861
rect 24581 13852 24593 13855
rect 23808 13824 24593 13852
rect 23808 13812 23814 13824
rect 24581 13821 24593 13824
rect 24627 13821 24639 13855
rect 24581 13815 24639 13821
rect 24670 13812 24676 13864
rect 24728 13852 24734 13864
rect 27798 13852 27804 13864
rect 24728 13824 24773 13852
rect 26206 13824 26648 13852
rect 24728 13812 24734 13824
rect 16172 13756 17264 13784
rect 16172 13744 16178 13756
rect 17402 13744 17408 13796
rect 17460 13784 17466 13796
rect 17460 13756 18000 13784
rect 17460 13744 17466 13756
rect 17678 13716 17684 13728
rect 15672 13688 17684 13716
rect 17678 13676 17684 13688
rect 17736 13676 17742 13728
rect 17972 13716 18000 13756
rect 22830 13744 22836 13796
rect 22888 13784 22894 13796
rect 26206 13784 26234 13824
rect 22888 13756 26234 13784
rect 22888 13744 22894 13756
rect 18322 13716 18328 13728
rect 17972 13688 18328 13716
rect 18322 13676 18328 13688
rect 18380 13676 18386 13728
rect 18690 13676 18696 13728
rect 18748 13716 18754 13728
rect 19337 13719 19395 13725
rect 19337 13716 19349 13719
rect 18748 13688 19349 13716
rect 18748 13676 18754 13688
rect 19337 13685 19349 13688
rect 19383 13716 19395 13719
rect 20990 13716 20996 13728
rect 19383 13688 20996 13716
rect 19383 13685 19395 13688
rect 19337 13679 19395 13685
rect 20990 13676 20996 13688
rect 21048 13676 21054 13728
rect 22002 13676 22008 13728
rect 22060 13716 22066 13728
rect 23937 13719 23995 13725
rect 23937 13716 23949 13719
rect 22060 13688 23949 13716
rect 22060 13676 22066 13688
rect 23937 13685 23949 13688
rect 23983 13685 23995 13719
rect 24210 13716 24216 13728
rect 24171 13688 24216 13716
rect 23937 13679 23995 13685
rect 24210 13676 24216 13688
rect 24268 13676 24274 13728
rect 26620 13716 26648 13824
rect 27448 13824 27804 13852
rect 26878 13744 26884 13796
rect 26936 13784 26942 13796
rect 26973 13787 27031 13793
rect 26973 13784 26985 13787
rect 26936 13756 26985 13784
rect 26936 13744 26942 13756
rect 26973 13753 26985 13756
rect 27019 13753 27031 13787
rect 26973 13747 27031 13753
rect 27154 13744 27160 13796
rect 27212 13784 27218 13796
rect 27341 13787 27399 13793
rect 27341 13784 27353 13787
rect 27212 13756 27353 13784
rect 27212 13744 27218 13756
rect 27341 13753 27353 13756
rect 27387 13753 27399 13787
rect 27341 13747 27399 13753
rect 27448 13716 27476 13824
rect 27798 13812 27804 13824
rect 27856 13812 27862 13864
rect 28368 13852 28396 13960
rect 28445 13957 28457 13991
rect 28491 13957 28503 13991
rect 28644 13991 28724 13997
rect 28644 13960 28673 13991
rect 28445 13951 28503 13957
rect 28661 13957 28673 13960
rect 28707 13957 28724 13991
rect 28661 13951 28724 13957
rect 28460 13920 28488 13951
rect 28718 13948 28724 13951
rect 28776 13948 28782 14000
rect 29917 13991 29975 13997
rect 29917 13957 29929 13991
rect 29963 13988 29975 13991
rect 29963 13960 31340 13988
rect 29963 13957 29975 13960
rect 29917 13951 29975 13957
rect 29178 13920 29184 13932
rect 28460 13892 29184 13920
rect 29178 13880 29184 13892
rect 29236 13880 29242 13932
rect 29273 13923 29331 13929
rect 29273 13889 29285 13923
rect 29319 13920 29331 13923
rect 30926 13920 30932 13932
rect 29319 13892 30932 13920
rect 29319 13889 29331 13892
rect 29273 13883 29331 13889
rect 30926 13880 30932 13892
rect 30984 13880 30990 13932
rect 31110 13920 31116 13932
rect 31071 13892 31116 13920
rect 31110 13880 31116 13892
rect 31168 13880 31174 13932
rect 31312 13929 31340 13960
rect 31297 13923 31355 13929
rect 31297 13889 31309 13923
rect 31343 13889 31355 13923
rect 31297 13883 31355 13889
rect 29086 13852 29092 13864
rect 28368 13824 29092 13852
rect 29086 13812 29092 13824
rect 29144 13812 29150 13864
rect 29730 13812 29736 13864
rect 29788 13852 29794 13864
rect 30285 13855 30343 13861
rect 30285 13852 30297 13855
rect 29788 13824 30297 13852
rect 29788 13812 29794 13824
rect 30285 13821 30297 13824
rect 30331 13821 30343 13855
rect 30834 13852 30840 13864
rect 30795 13824 30840 13852
rect 30285 13815 30343 13821
rect 30834 13812 30840 13824
rect 30892 13812 30898 13864
rect 29825 13787 29883 13793
rect 29825 13753 29837 13787
rect 29871 13784 29883 13787
rect 29917 13787 29975 13793
rect 29917 13784 29929 13787
rect 29871 13756 29929 13784
rect 29871 13753 29883 13756
rect 29825 13747 29883 13753
rect 29917 13753 29929 13756
rect 29963 13753 29975 13787
rect 29917 13747 29975 13753
rect 28626 13716 28632 13728
rect 26620 13688 27476 13716
rect 28587 13688 28632 13716
rect 28626 13676 28632 13688
rect 28684 13676 28690 13728
rect 29638 13716 29644 13728
rect 29599 13688 29644 13716
rect 29638 13676 29644 13688
rect 29696 13676 29702 13728
rect 1104 13626 32016 13648
rect 0 13580 800 13594
rect 0 13552 888 13580
rect 1104 13574 2136 13626
rect 2188 13574 12440 13626
rect 12492 13574 22744 13626
rect 22796 13574 32016 13626
rect 32320 13580 33120 13594
rect 1104 13552 32016 13574
rect 32048 13552 33120 13580
rect 0 13538 800 13552
rect 860 13444 888 13552
rect 2682 13512 2688 13524
rect 2643 13484 2688 13512
rect 2682 13472 2688 13484
rect 2740 13472 2746 13524
rect 3050 13512 3056 13524
rect 3011 13484 3056 13512
rect 3050 13472 3056 13484
rect 3108 13472 3114 13524
rect 3142 13472 3148 13524
rect 3200 13472 3206 13524
rect 7098 13512 7104 13524
rect 7059 13484 7104 13512
rect 7098 13472 7104 13484
rect 7156 13512 7162 13524
rect 7466 13512 7472 13524
rect 7156 13484 7472 13512
rect 7156 13472 7162 13484
rect 7466 13472 7472 13484
rect 7524 13472 7530 13524
rect 7653 13515 7711 13521
rect 7653 13481 7665 13515
rect 7699 13512 7711 13515
rect 7742 13512 7748 13524
rect 7699 13484 7748 13512
rect 7699 13481 7711 13484
rect 7653 13475 7711 13481
rect 7742 13472 7748 13484
rect 7800 13472 7806 13524
rect 8662 13472 8668 13524
rect 8720 13512 8726 13524
rect 16577 13515 16635 13521
rect 8720 13484 16436 13512
rect 8720 13472 8726 13484
rect 860 13416 1440 13444
rect 1412 13385 1440 13416
rect 2314 13404 2320 13456
rect 2372 13444 2378 13456
rect 3160 13444 3188 13472
rect 3602 13444 3608 13456
rect 2372 13416 3608 13444
rect 2372 13404 2378 13416
rect 3602 13404 3608 13416
rect 3660 13404 3666 13456
rect 4341 13447 4399 13453
rect 4341 13413 4353 13447
rect 4387 13444 4399 13447
rect 4706 13444 4712 13456
rect 4387 13416 4712 13444
rect 4387 13413 4399 13416
rect 4341 13407 4399 13413
rect 4706 13404 4712 13416
rect 4764 13404 4770 13456
rect 7558 13404 7564 13456
rect 7616 13444 7622 13456
rect 8018 13444 8024 13456
rect 7616 13416 8024 13444
rect 7616 13404 7622 13416
rect 8018 13404 8024 13416
rect 8076 13404 8082 13456
rect 8386 13444 8392 13456
rect 8220 13416 8392 13444
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13345 1455 13379
rect 1397 13339 1455 13345
rect 1486 13336 1492 13388
rect 1544 13376 1550 13388
rect 3145 13379 3203 13385
rect 1544 13348 3096 13376
rect 1544 13336 1550 13348
rect 1673 13311 1731 13317
rect 1673 13277 1685 13311
rect 1719 13308 1731 13311
rect 2498 13308 2504 13320
rect 1719 13280 2504 13308
rect 1719 13277 1731 13280
rect 1673 13271 1731 13277
rect 2498 13268 2504 13280
rect 2556 13268 2562 13320
rect 2869 13311 2927 13317
rect 2869 13277 2881 13311
rect 2915 13277 2927 13311
rect 3068 13308 3096 13348
rect 3145 13345 3157 13379
rect 3191 13376 3203 13379
rect 3970 13376 3976 13388
rect 3191 13348 3976 13376
rect 3191 13345 3203 13348
rect 3145 13339 3203 13345
rect 3970 13336 3976 13348
rect 4028 13336 4034 13388
rect 5442 13336 5448 13388
rect 5500 13336 5506 13388
rect 6822 13336 6828 13388
rect 6880 13376 6886 13388
rect 8113 13379 8171 13385
rect 8113 13376 8125 13379
rect 6880 13348 8125 13376
rect 6880 13336 6886 13348
rect 8113 13345 8125 13348
rect 8159 13345 8171 13379
rect 8113 13339 8171 13345
rect 3786 13308 3792 13320
rect 3068 13280 3792 13308
rect 2869 13271 2927 13277
rect 2884 13172 2912 13271
rect 3786 13268 3792 13280
rect 3844 13308 3850 13320
rect 4982 13308 4988 13320
rect 3844 13280 4988 13308
rect 3844 13268 3850 13280
rect 4982 13268 4988 13280
rect 5040 13308 5046 13320
rect 5040 13280 5672 13308
rect 5040 13268 5046 13280
rect 3970 13240 3976 13252
rect 3931 13212 3976 13240
rect 3970 13200 3976 13212
rect 4028 13200 4034 13252
rect 5353 13243 5411 13249
rect 5353 13240 5365 13243
rect 4448 13212 5365 13240
rect 3510 13172 3516 13184
rect 2884 13144 3516 13172
rect 3510 13132 3516 13144
rect 3568 13132 3574 13184
rect 4448 13181 4476 13212
rect 5353 13209 5365 13212
rect 5399 13209 5411 13243
rect 5353 13203 5411 13209
rect 5445 13243 5503 13249
rect 5445 13209 5457 13243
rect 5491 13240 5503 13243
rect 5534 13240 5540 13252
rect 5491 13212 5540 13240
rect 5491 13209 5503 13212
rect 5445 13203 5503 13209
rect 5534 13200 5540 13212
rect 5592 13200 5598 13252
rect 5644 13240 5672 13280
rect 5718 13268 5724 13320
rect 5776 13308 5782 13320
rect 5813 13311 5871 13317
rect 5813 13308 5825 13311
rect 5776 13280 5825 13308
rect 5776 13268 5782 13280
rect 5813 13277 5825 13280
rect 5859 13277 5871 13311
rect 5813 13271 5871 13277
rect 6914 13268 6920 13320
rect 6972 13308 6978 13320
rect 7009 13311 7067 13317
rect 7009 13308 7021 13311
rect 6972 13280 7021 13308
rect 6972 13268 6978 13280
rect 7009 13277 7021 13280
rect 7055 13308 7067 13311
rect 8220 13308 8248 13416
rect 8386 13404 8392 13416
rect 8444 13404 8450 13456
rect 8478 13404 8484 13456
rect 8536 13444 8542 13456
rect 10410 13444 10416 13456
rect 8536 13416 10416 13444
rect 8536 13404 8542 13416
rect 10410 13404 10416 13416
rect 10468 13404 10474 13456
rect 11514 13404 11520 13456
rect 11572 13444 11578 13456
rect 14185 13447 14243 13453
rect 11572 13416 12848 13444
rect 11572 13404 11578 13416
rect 8297 13379 8355 13385
rect 8297 13345 8309 13379
rect 8343 13345 8355 13379
rect 9398 13376 9404 13388
rect 9359 13348 9404 13376
rect 8297 13339 8355 13345
rect 7055 13280 8248 13308
rect 8312 13308 8340 13339
rect 9398 13336 9404 13348
rect 9456 13336 9462 13388
rect 9125 13311 9183 13317
rect 9125 13308 9137 13311
rect 8312 13280 9137 13308
rect 7055 13277 7067 13280
rect 7009 13271 7067 13277
rect 9125 13277 9137 13280
rect 9171 13277 9183 13311
rect 9125 13271 9183 13277
rect 10505 13311 10563 13317
rect 10505 13277 10517 13311
rect 10551 13308 10563 13311
rect 12158 13308 12164 13320
rect 10551 13280 12164 13308
rect 10551 13277 10563 13280
rect 10505 13271 10563 13277
rect 8754 13240 8760 13252
rect 5644 13212 8760 13240
rect 8754 13200 8760 13212
rect 8812 13200 8818 13252
rect 4433 13175 4491 13181
rect 4433 13141 4445 13175
rect 4479 13141 4491 13175
rect 4433 13135 4491 13141
rect 4798 13132 4804 13184
rect 4856 13172 4862 13184
rect 5077 13175 5135 13181
rect 5077 13172 5089 13175
rect 4856 13144 5089 13172
rect 4856 13132 4862 13144
rect 5077 13141 5089 13144
rect 5123 13141 5135 13175
rect 6178 13172 6184 13184
rect 6139 13144 6184 13172
rect 5077 13135 5135 13141
rect 6178 13132 6184 13144
rect 6236 13132 6242 13184
rect 6365 13175 6423 13181
rect 6365 13141 6377 13175
rect 6411 13172 6423 13175
rect 7098 13172 7104 13184
rect 6411 13144 7104 13172
rect 6411 13141 6423 13144
rect 6365 13135 6423 13141
rect 7098 13132 7104 13144
rect 7156 13132 7162 13184
rect 7650 13132 7656 13184
rect 7708 13172 7714 13184
rect 8021 13175 8079 13181
rect 8021 13172 8033 13175
rect 7708 13144 8033 13172
rect 7708 13132 7714 13144
rect 8021 13141 8033 13144
rect 8067 13141 8079 13175
rect 9140 13172 9168 13271
rect 12158 13268 12164 13280
rect 12216 13268 12222 13320
rect 12529 13311 12587 13317
rect 12529 13277 12541 13311
rect 12575 13308 12587 13311
rect 12618 13308 12624 13320
rect 12575 13280 12624 13308
rect 12575 13277 12587 13280
rect 12529 13271 12587 13277
rect 12618 13268 12624 13280
rect 12676 13268 12682 13320
rect 12820 13317 12848 13416
rect 14185 13413 14197 13447
rect 14231 13444 14243 13447
rect 15102 13444 15108 13456
rect 14231 13416 15108 13444
rect 14231 13413 14243 13416
rect 14185 13407 14243 13413
rect 15102 13404 15108 13416
rect 15160 13404 15166 13456
rect 15381 13447 15439 13453
rect 15381 13413 15393 13447
rect 15427 13444 15439 13447
rect 15930 13444 15936 13456
rect 15427 13416 15936 13444
rect 15427 13413 15439 13416
rect 15381 13407 15439 13413
rect 15930 13404 15936 13416
rect 15988 13404 15994 13456
rect 16408 13444 16436 13484
rect 16577 13481 16589 13515
rect 16623 13512 16635 13515
rect 16758 13512 16764 13524
rect 16623 13484 16764 13512
rect 16623 13481 16635 13484
rect 16577 13475 16635 13481
rect 16758 13472 16764 13484
rect 16816 13472 16822 13524
rect 16850 13472 16856 13524
rect 16908 13512 16914 13524
rect 17126 13512 17132 13524
rect 16908 13484 17132 13512
rect 16908 13472 16914 13484
rect 17126 13472 17132 13484
rect 17184 13472 17190 13524
rect 17313 13515 17371 13521
rect 17313 13481 17325 13515
rect 17359 13512 17371 13515
rect 17770 13512 17776 13524
rect 17359 13484 17776 13512
rect 17359 13481 17371 13484
rect 17313 13475 17371 13481
rect 17770 13472 17776 13484
rect 17828 13512 17834 13524
rect 17828 13484 18276 13512
rect 17828 13472 17834 13484
rect 18138 13444 18144 13456
rect 16408 13416 18144 13444
rect 18138 13404 18144 13416
rect 18196 13404 18202 13456
rect 18248 13444 18276 13484
rect 18322 13472 18328 13524
rect 18380 13512 18386 13524
rect 18417 13515 18475 13521
rect 18417 13512 18429 13515
rect 18380 13484 18429 13512
rect 18380 13472 18386 13484
rect 18417 13481 18429 13484
rect 18463 13512 18475 13515
rect 19334 13512 19340 13524
rect 18463 13484 19340 13512
rect 18463 13481 18475 13484
rect 18417 13475 18475 13481
rect 19334 13472 19340 13484
rect 19392 13472 19398 13524
rect 19429 13515 19487 13521
rect 19429 13481 19441 13515
rect 19475 13512 19487 13515
rect 19475 13484 20944 13512
rect 19475 13481 19487 13484
rect 19429 13475 19487 13481
rect 19794 13444 19800 13456
rect 18248 13416 19800 13444
rect 19794 13404 19800 13416
rect 19852 13404 19858 13456
rect 20916 13444 20944 13484
rect 21726 13472 21732 13524
rect 21784 13512 21790 13524
rect 21821 13515 21879 13521
rect 21821 13512 21833 13515
rect 21784 13484 21833 13512
rect 21784 13472 21790 13484
rect 21821 13481 21833 13484
rect 21867 13481 21879 13515
rect 21821 13475 21879 13481
rect 22094 13472 22100 13524
rect 22152 13512 22158 13524
rect 22189 13515 22247 13521
rect 22189 13512 22201 13515
rect 22152 13484 22201 13512
rect 22152 13472 22158 13484
rect 22189 13481 22201 13484
rect 22235 13481 22247 13515
rect 22189 13475 22247 13481
rect 23566 13472 23572 13524
rect 23624 13512 23630 13524
rect 24302 13512 24308 13524
rect 23624 13484 24308 13512
rect 23624 13472 23630 13484
rect 24302 13472 24308 13484
rect 24360 13472 24366 13524
rect 25498 13512 25504 13524
rect 24780 13484 25504 13512
rect 24780 13444 24808 13484
rect 25498 13472 25504 13484
rect 25556 13472 25562 13524
rect 25774 13472 25780 13524
rect 25832 13512 25838 13524
rect 26145 13515 26203 13521
rect 26145 13512 26157 13515
rect 25832 13484 26157 13512
rect 25832 13472 25838 13484
rect 26145 13481 26157 13484
rect 26191 13481 26203 13515
rect 26145 13475 26203 13481
rect 26510 13472 26516 13524
rect 26568 13512 26574 13524
rect 26973 13515 27031 13521
rect 26973 13512 26985 13515
rect 26568 13484 26985 13512
rect 26568 13472 26574 13484
rect 26973 13481 26985 13484
rect 27019 13512 27031 13515
rect 27154 13512 27160 13524
rect 27019 13484 27160 13512
rect 27019 13481 27031 13484
rect 26973 13475 27031 13481
rect 27154 13472 27160 13484
rect 27212 13472 27218 13524
rect 27338 13472 27344 13524
rect 27396 13512 27402 13524
rect 27617 13515 27675 13521
rect 27617 13512 27629 13515
rect 27396 13484 27629 13512
rect 27396 13472 27402 13484
rect 27617 13481 27629 13484
rect 27663 13481 27675 13515
rect 27617 13475 27675 13481
rect 28537 13515 28595 13521
rect 28537 13481 28549 13515
rect 28583 13512 28595 13515
rect 28626 13512 28632 13524
rect 28583 13484 28632 13512
rect 28583 13481 28595 13484
rect 28537 13475 28595 13481
rect 28626 13472 28632 13484
rect 28684 13512 28690 13524
rect 28813 13515 28871 13521
rect 28813 13512 28825 13515
rect 28684 13484 28825 13512
rect 28684 13472 28690 13484
rect 28813 13481 28825 13484
rect 28859 13481 28871 13515
rect 28813 13475 28871 13481
rect 28997 13515 29055 13521
rect 28997 13481 29009 13515
rect 29043 13512 29055 13515
rect 29086 13512 29092 13524
rect 29043 13484 29092 13512
rect 29043 13481 29055 13484
rect 28997 13475 29055 13481
rect 29086 13472 29092 13484
rect 29144 13472 29150 13524
rect 29914 13512 29920 13524
rect 29875 13484 29920 13512
rect 29914 13472 29920 13484
rect 29972 13472 29978 13524
rect 30926 13512 30932 13524
rect 30887 13484 30932 13512
rect 30926 13472 30932 13484
rect 30984 13472 30990 13524
rect 31110 13512 31116 13524
rect 31071 13484 31116 13512
rect 31110 13472 31116 13484
rect 31168 13472 31174 13524
rect 20916 13416 24808 13444
rect 25958 13404 25964 13456
rect 26016 13444 26022 13456
rect 32048 13444 32076 13552
rect 32320 13538 33120 13552
rect 26016 13416 32076 13444
rect 26016 13404 26022 13416
rect 15746 13376 15752 13388
rect 14108 13348 15516 13376
rect 12805 13311 12863 13317
rect 12805 13277 12817 13311
rect 12851 13277 12863 13311
rect 12986 13308 12992 13320
rect 12947 13280 12992 13308
rect 12805 13271 12863 13277
rect 12986 13268 12992 13280
rect 13044 13268 13050 13320
rect 14108 13317 14136 13348
rect 14093 13311 14151 13317
rect 14093 13277 14105 13311
rect 14139 13277 14151 13311
rect 14093 13271 14151 13277
rect 14182 13268 14188 13320
rect 14240 13308 14246 13320
rect 14642 13318 14648 13320
rect 14277 13311 14335 13317
rect 14277 13308 14289 13311
rect 14240 13280 14289 13308
rect 14240 13268 14246 13280
rect 14277 13277 14289 13280
rect 14323 13308 14335 13311
rect 14568 13308 14648 13318
rect 14323 13290 14648 13308
rect 14323 13280 14596 13290
rect 14323 13277 14335 13280
rect 14277 13271 14335 13277
rect 14642 13268 14648 13290
rect 14700 13318 14706 13320
rect 14700 13290 15047 13318
rect 14700 13268 14706 13290
rect 10772 13243 10830 13249
rect 10772 13209 10784 13243
rect 10818 13240 10830 13243
rect 11330 13240 11336 13252
rect 10818 13212 11336 13240
rect 10818 13209 10830 13212
rect 10772 13203 10830 13209
rect 11330 13200 11336 13212
rect 11388 13200 11394 13252
rect 13906 13200 13912 13252
rect 13964 13240 13970 13252
rect 14829 13243 14887 13249
rect 14829 13240 14841 13243
rect 13964 13212 14841 13240
rect 13964 13200 13970 13212
rect 14829 13209 14841 13212
rect 14875 13240 14887 13243
rect 14918 13240 14924 13252
rect 14875 13212 14924 13240
rect 14875 13209 14887 13212
rect 14829 13203 14887 13209
rect 14918 13200 14924 13212
rect 14976 13200 14982 13252
rect 15019 13249 15047 13290
rect 15102 13268 15108 13320
rect 15160 13308 15166 13320
rect 15381 13311 15439 13317
rect 15381 13308 15393 13311
rect 15160 13280 15393 13308
rect 15160 13268 15166 13280
rect 15381 13277 15393 13280
rect 15427 13277 15439 13311
rect 15381 13271 15439 13277
rect 15013 13243 15071 13249
rect 15013 13209 15025 13243
rect 15059 13209 15071 13243
rect 15013 13203 15071 13209
rect 11885 13175 11943 13181
rect 11885 13172 11897 13175
rect 9140 13144 11897 13172
rect 8021 13135 8079 13141
rect 11885 13141 11897 13144
rect 11931 13141 11943 13175
rect 12342 13172 12348 13184
rect 12303 13144 12348 13172
rect 11885 13135 11943 13141
rect 12342 13132 12348 13144
rect 12400 13132 12406 13184
rect 12802 13132 12808 13184
rect 12860 13172 12866 13184
rect 15102 13172 15108 13184
rect 12860 13144 15108 13172
rect 12860 13132 12866 13144
rect 15102 13132 15108 13144
rect 15160 13132 15166 13184
rect 15488 13172 15516 13348
rect 15580 13348 15752 13376
rect 15580 13317 15608 13348
rect 15746 13336 15752 13348
rect 15804 13336 15810 13388
rect 16206 13376 16212 13388
rect 16167 13348 16212 13376
rect 16206 13336 16212 13348
rect 16264 13336 16270 13388
rect 19426 13376 19432 13388
rect 17788 13348 19432 13376
rect 15565 13311 15623 13317
rect 15565 13277 15577 13311
rect 15611 13277 15623 13311
rect 15565 13271 15623 13277
rect 16298 13268 16304 13320
rect 16356 13308 16362 13320
rect 16393 13311 16451 13317
rect 16393 13308 16405 13311
rect 16356 13280 16405 13308
rect 16356 13268 16362 13280
rect 16393 13277 16405 13280
rect 16439 13277 16451 13311
rect 16393 13271 16451 13277
rect 16482 13268 16488 13320
rect 16540 13308 16546 13320
rect 17788 13308 17816 13348
rect 19426 13336 19432 13348
rect 19484 13336 19490 13388
rect 19978 13376 19984 13388
rect 19939 13348 19984 13376
rect 19978 13336 19984 13348
rect 20036 13336 20042 13388
rect 20990 13336 20996 13388
rect 21048 13376 21054 13388
rect 22281 13379 22339 13385
rect 22281 13376 22293 13379
rect 21048 13348 22293 13376
rect 21048 13336 21054 13348
rect 22281 13345 22293 13348
rect 22327 13345 22339 13379
rect 22281 13339 22339 13345
rect 22370 13336 22376 13388
rect 22428 13376 22434 13388
rect 22554 13376 22560 13388
rect 22428 13348 22560 13376
rect 22428 13336 22434 13348
rect 22554 13336 22560 13348
rect 22612 13376 22618 13388
rect 24762 13376 24768 13388
rect 22612 13348 23704 13376
rect 24723 13348 24768 13376
rect 22612 13336 22618 13348
rect 18782 13308 18788 13320
rect 16540 13280 17816 13308
rect 17871 13280 18788 13308
rect 16540 13268 16546 13280
rect 15749 13243 15807 13249
rect 15749 13209 15761 13243
rect 15795 13240 15807 13243
rect 15838 13240 15844 13252
rect 15795 13212 15844 13240
rect 15795 13209 15807 13212
rect 15749 13203 15807 13209
rect 15838 13200 15844 13212
rect 15896 13200 15902 13252
rect 17221 13243 17279 13249
rect 15948 13212 16620 13240
rect 15948 13172 15976 13212
rect 15488 13144 15976 13172
rect 16592 13172 16620 13212
rect 17221 13209 17233 13243
rect 17267 13240 17279 13243
rect 17494 13240 17500 13252
rect 17267 13212 17500 13240
rect 17267 13209 17279 13212
rect 17221 13203 17279 13209
rect 17494 13200 17500 13212
rect 17552 13200 17558 13252
rect 17871 13240 17899 13280
rect 18782 13268 18788 13280
rect 18840 13268 18846 13320
rect 19150 13268 19156 13320
rect 19208 13308 19214 13320
rect 19337 13311 19395 13317
rect 19337 13308 19349 13311
rect 19208 13280 19349 13308
rect 19208 13268 19214 13280
rect 19337 13277 19349 13280
rect 19383 13308 19395 13311
rect 19383 13280 20484 13308
rect 19383 13277 19395 13280
rect 19337 13271 19395 13277
rect 17788 13212 17899 13240
rect 17788 13172 17816 13212
rect 17954 13200 17960 13252
rect 18012 13240 18018 13252
rect 18012 13212 18057 13240
rect 18012 13200 18018 13212
rect 18138 13200 18144 13252
rect 18196 13240 18202 13252
rect 20226 13243 20284 13249
rect 20226 13240 20238 13243
rect 18196 13212 20238 13240
rect 18196 13200 18202 13212
rect 20226 13209 20238 13212
rect 20272 13209 20284 13243
rect 20456 13240 20484 13280
rect 21818 13268 21824 13320
rect 21876 13308 21882 13320
rect 22005 13311 22063 13317
rect 22005 13308 22017 13311
rect 21876 13280 22017 13308
rect 21876 13268 21882 13280
rect 22005 13277 22017 13280
rect 22051 13277 22063 13311
rect 23382 13308 23388 13320
rect 23343 13280 23388 13308
rect 22005 13271 22063 13277
rect 23382 13268 23388 13280
rect 23440 13268 23446 13320
rect 23676 13317 23704 13348
rect 24762 13336 24768 13348
rect 24820 13336 24826 13388
rect 27062 13376 27068 13388
rect 27023 13348 27068 13376
rect 27062 13336 27068 13348
rect 27120 13336 27126 13388
rect 27448 13348 27660 13376
rect 23661 13311 23719 13317
rect 23661 13277 23673 13311
rect 23707 13277 23719 13311
rect 23661 13271 23719 13277
rect 23845 13311 23903 13317
rect 23845 13277 23857 13311
rect 23891 13308 23903 13311
rect 23934 13308 23940 13320
rect 23891 13280 23940 13308
rect 23891 13277 23903 13280
rect 23845 13271 23903 13277
rect 23934 13268 23940 13280
rect 23992 13268 23998 13320
rect 24210 13268 24216 13320
rect 24268 13308 24274 13320
rect 25021 13311 25079 13317
rect 25021 13308 25033 13311
rect 24268 13280 25033 13308
rect 24268 13268 24274 13280
rect 25021 13277 25033 13280
rect 25067 13277 25079 13311
rect 26786 13308 26792 13320
rect 26747 13280 26792 13308
rect 25021 13271 25079 13277
rect 26786 13268 26792 13280
rect 26844 13268 26850 13320
rect 22554 13240 22560 13252
rect 20456 13212 22560 13240
rect 20226 13203 20284 13209
rect 22554 13200 22560 13212
rect 22612 13200 22618 13252
rect 22922 13200 22928 13252
rect 22980 13240 22986 13252
rect 23952 13240 23980 13268
rect 24670 13240 24676 13252
rect 22980 13212 23704 13240
rect 23952 13212 24676 13240
rect 22980 13200 22986 13212
rect 16592 13144 17816 13172
rect 18233 13175 18291 13181
rect 18233 13141 18245 13175
rect 18279 13172 18291 13175
rect 18417 13175 18475 13181
rect 18417 13172 18429 13175
rect 18279 13144 18429 13172
rect 18279 13141 18291 13144
rect 18233 13135 18291 13141
rect 18417 13141 18429 13144
rect 18463 13141 18475 13175
rect 18417 13135 18475 13141
rect 19242 13132 19248 13184
rect 19300 13172 19306 13184
rect 21361 13175 21419 13181
rect 21361 13172 21373 13175
rect 19300 13144 21373 13172
rect 19300 13132 19306 13144
rect 21361 13141 21373 13144
rect 21407 13172 21419 13175
rect 21910 13172 21916 13184
rect 21407 13144 21916 13172
rect 21407 13141 21419 13144
rect 21361 13135 21419 13141
rect 21910 13132 21916 13144
rect 21968 13132 21974 13184
rect 23201 13175 23259 13181
rect 23201 13141 23213 13175
rect 23247 13172 23259 13175
rect 23566 13172 23572 13184
rect 23247 13144 23572 13172
rect 23247 13141 23259 13144
rect 23201 13135 23259 13141
rect 23566 13132 23572 13144
rect 23624 13132 23630 13184
rect 23676 13172 23704 13212
rect 24670 13200 24676 13212
rect 24728 13200 24734 13252
rect 25682 13200 25688 13252
rect 25740 13240 25746 13252
rect 27448 13240 27476 13348
rect 27525 13311 27583 13317
rect 27525 13277 27537 13311
rect 27571 13277 27583 13311
rect 27632 13308 27660 13348
rect 27706 13336 27712 13388
rect 27764 13376 27770 13388
rect 27801 13379 27859 13385
rect 27801 13376 27813 13379
rect 27764 13348 27813 13376
rect 27764 13336 27770 13348
rect 27801 13345 27813 13348
rect 27847 13345 27859 13379
rect 27801 13339 27859 13345
rect 28718 13336 28724 13388
rect 28776 13376 28782 13388
rect 28776 13348 30696 13376
rect 28776 13336 28782 13348
rect 28537 13311 28595 13317
rect 28537 13308 28549 13311
rect 27632 13280 28549 13308
rect 27525 13271 27583 13277
rect 28537 13277 28549 13280
rect 28583 13277 28595 13311
rect 28537 13271 28595 13277
rect 25740 13212 27476 13240
rect 25740 13200 25746 13212
rect 26326 13172 26332 13184
rect 23676 13144 26332 13172
rect 26326 13132 26332 13144
rect 26384 13132 26390 13184
rect 26605 13175 26663 13181
rect 26605 13141 26617 13175
rect 26651 13172 26663 13175
rect 26970 13172 26976 13184
rect 26651 13144 26976 13172
rect 26651 13141 26663 13144
rect 26605 13135 26663 13141
rect 26970 13132 26976 13144
rect 27028 13132 27034 13184
rect 27540 13172 27568 13271
rect 28902 13268 28908 13320
rect 28960 13308 28966 13320
rect 29733 13311 29791 13317
rect 29733 13308 29745 13311
rect 28960 13280 29745 13308
rect 28960 13268 28966 13280
rect 29733 13277 29745 13280
rect 29779 13277 29791 13311
rect 29733 13271 29791 13277
rect 30009 13311 30067 13317
rect 30009 13277 30021 13311
rect 30055 13308 30067 13311
rect 30190 13308 30196 13320
rect 30055 13280 30196 13308
rect 30055 13277 30067 13280
rect 30009 13271 30067 13277
rect 30190 13268 30196 13280
rect 30248 13268 30254 13320
rect 28629 13243 28687 13249
rect 28629 13209 28641 13243
rect 28675 13240 28687 13243
rect 29638 13240 29644 13252
rect 28675 13212 29644 13240
rect 28675 13209 28687 13212
rect 28629 13203 28687 13209
rect 29638 13200 29644 13212
rect 29696 13200 29702 13252
rect 30561 13243 30619 13249
rect 30561 13209 30573 13243
rect 30607 13209 30619 13243
rect 30668 13240 30696 13348
rect 30938 13243 30996 13249
rect 30938 13240 30950 13243
rect 30668 13212 30950 13240
rect 30561 13203 30619 13209
rect 30938 13209 30950 13212
rect 30984 13209 30996 13243
rect 30938 13203 30996 13209
rect 27614 13172 27620 13184
rect 27540 13144 27620 13172
rect 27614 13132 27620 13144
rect 27672 13132 27678 13184
rect 27801 13175 27859 13181
rect 27801 13141 27813 13175
rect 27847 13172 27859 13175
rect 28718 13172 28724 13184
rect 27847 13144 28724 13172
rect 27847 13141 27859 13144
rect 27801 13135 27859 13141
rect 28718 13132 28724 13144
rect 28776 13132 28782 13184
rect 28810 13132 28816 13184
rect 28868 13181 28874 13184
rect 28868 13175 28887 13181
rect 28875 13141 28887 13175
rect 29546 13172 29552 13184
rect 29507 13144 29552 13172
rect 28868 13135 28887 13141
rect 28868 13132 28874 13135
rect 29546 13132 29552 13144
rect 29604 13132 29610 13184
rect 30576 13172 30604 13203
rect 31018 13172 31024 13184
rect 30576 13144 31024 13172
rect 31018 13132 31024 13144
rect 31076 13132 31082 13184
rect 1104 13082 32016 13104
rect 1104 13030 7288 13082
rect 7340 13030 17592 13082
rect 17644 13030 27896 13082
rect 27948 13030 32016 13082
rect 1104 13008 32016 13030
rect 2133 12971 2191 12977
rect 2133 12937 2145 12971
rect 2179 12968 2191 12971
rect 3510 12968 3516 12980
rect 2179 12940 3516 12968
rect 2179 12937 2191 12940
rect 2133 12931 2191 12937
rect 3510 12928 3516 12940
rect 3568 12928 3574 12980
rect 4617 12971 4675 12977
rect 4617 12968 4629 12971
rect 3896 12940 4629 12968
rect 1486 12900 1492 12912
rect 1447 12872 1492 12900
rect 1486 12860 1492 12872
rect 1544 12860 1550 12912
rect 2866 12900 2872 12912
rect 2608 12872 2872 12900
rect 2314 12832 2320 12844
rect 2275 12804 2320 12832
rect 2314 12792 2320 12804
rect 2372 12792 2378 12844
rect 2608 12841 2636 12872
rect 2866 12860 2872 12872
rect 2924 12860 2930 12912
rect 2976 12872 3740 12900
rect 2593 12835 2651 12841
rect 2593 12801 2605 12835
rect 2639 12801 2651 12835
rect 2593 12795 2651 12801
rect 2774 12792 2780 12844
rect 2832 12832 2838 12844
rect 2976 12832 3004 12872
rect 3712 12841 3740 12872
rect 2832 12804 3004 12832
rect 3421 12835 3479 12841
rect 2832 12792 2838 12804
rect 3421 12801 3433 12835
rect 3467 12801 3479 12835
rect 3421 12795 3479 12801
rect 3697 12835 3755 12841
rect 3697 12801 3709 12835
rect 3743 12801 3755 12835
rect 3697 12795 3755 12801
rect 1302 12724 1308 12776
rect 1360 12764 1366 12776
rect 1360 12736 2360 12764
rect 1360 12724 1366 12736
rect 1673 12699 1731 12705
rect 1673 12665 1685 12699
rect 1719 12696 1731 12699
rect 1854 12696 1860 12708
rect 1719 12668 1860 12696
rect 1719 12665 1731 12668
rect 1673 12659 1731 12665
rect 1854 12656 1860 12668
rect 1912 12656 1918 12708
rect 2332 12696 2360 12736
rect 2406 12724 2412 12776
rect 2464 12764 2470 12776
rect 3436 12764 3464 12795
rect 2464 12736 3464 12764
rect 2464 12724 2470 12736
rect 3896 12696 3924 12940
rect 4617 12937 4629 12940
rect 4663 12937 4675 12971
rect 4798 12968 4804 12980
rect 4759 12940 4804 12968
rect 4617 12931 4675 12937
rect 4798 12928 4804 12940
rect 4856 12928 4862 12980
rect 5169 12971 5227 12977
rect 5169 12937 5181 12971
rect 5215 12968 5227 12971
rect 7558 12968 7564 12980
rect 5215 12940 7564 12968
rect 5215 12937 5227 12940
rect 5169 12931 5227 12937
rect 7558 12928 7564 12940
rect 7616 12928 7622 12980
rect 8021 12971 8079 12977
rect 7668 12940 7972 12968
rect 4062 12860 4068 12912
rect 4120 12900 4126 12912
rect 5261 12903 5319 12909
rect 5261 12900 5273 12903
rect 4120 12872 5273 12900
rect 4120 12860 4126 12872
rect 5261 12869 5273 12872
rect 5307 12900 5319 12903
rect 5350 12900 5356 12912
rect 5307 12872 5356 12900
rect 5307 12869 5319 12872
rect 5261 12863 5319 12869
rect 5350 12860 5356 12872
rect 5408 12860 5414 12912
rect 5828 12872 6500 12900
rect 4338 12832 4344 12844
rect 4299 12804 4344 12832
rect 4338 12792 4344 12804
rect 4396 12792 4402 12844
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 5828 12832 5856 12872
rect 4663 12804 5856 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 5902 12792 5908 12844
rect 5960 12832 5966 12844
rect 6270 12832 6276 12844
rect 5960 12804 6276 12832
rect 5960 12792 5966 12804
rect 6270 12792 6276 12804
rect 6328 12832 6334 12844
rect 6365 12835 6423 12841
rect 6365 12832 6377 12835
rect 6328 12804 6377 12832
rect 6328 12792 6334 12804
rect 6365 12801 6377 12804
rect 6411 12801 6423 12835
rect 6472 12832 6500 12872
rect 7098 12860 7104 12912
rect 7156 12900 7162 12912
rect 7668 12900 7696 12940
rect 7156 12872 7696 12900
rect 7944 12900 7972 12940
rect 8021 12937 8033 12971
rect 8067 12968 8079 12971
rect 8202 12968 8208 12980
rect 8067 12940 8208 12968
rect 8067 12937 8079 12940
rect 8021 12931 8079 12937
rect 8202 12928 8208 12940
rect 8260 12928 8266 12980
rect 8662 12928 8668 12980
rect 8720 12968 8726 12980
rect 14182 12968 14188 12980
rect 8720 12940 14188 12968
rect 8720 12928 8726 12940
rect 14182 12928 14188 12940
rect 14240 12928 14246 12980
rect 14918 12928 14924 12980
rect 14976 12968 14982 12980
rect 20162 12968 20168 12980
rect 14976 12940 20168 12968
rect 14976 12928 14982 12940
rect 20162 12928 20168 12940
rect 20220 12928 20226 12980
rect 20714 12928 20720 12980
rect 20772 12968 20778 12980
rect 25958 12968 25964 12980
rect 20772 12940 25964 12968
rect 20772 12928 20778 12940
rect 25958 12928 25964 12940
rect 26016 12928 26022 12980
rect 26786 12928 26792 12980
rect 26844 12968 26850 12980
rect 26973 12971 27031 12977
rect 26973 12968 26985 12971
rect 26844 12940 26985 12968
rect 26844 12928 26850 12940
rect 26973 12937 26985 12940
rect 27019 12937 27031 12971
rect 29638 12968 29644 12980
rect 29599 12940 29644 12968
rect 26973 12931 27031 12937
rect 29638 12928 29644 12940
rect 29696 12928 29702 12980
rect 11514 12900 11520 12912
rect 7944 12872 11520 12900
rect 7156 12860 7162 12872
rect 11514 12860 11520 12872
rect 11572 12860 11578 12912
rect 14277 12903 14335 12909
rect 14277 12900 14289 12903
rect 11624 12872 14289 12900
rect 7834 12841 7840 12844
rect 7823 12835 7840 12841
rect 7823 12832 7835 12835
rect 6472 12804 7835 12832
rect 6365 12795 6423 12801
rect 7823 12801 7835 12804
rect 7892 12830 7898 12844
rect 8202 12832 8208 12844
rect 7935 12830 8208 12832
rect 7892 12804 8208 12830
rect 7892 12802 7963 12804
rect 7823 12795 7840 12801
rect 7834 12792 7840 12795
rect 7892 12792 7898 12802
rect 8202 12792 8208 12804
rect 8260 12792 8266 12844
rect 8386 12792 8392 12844
rect 8444 12832 8450 12844
rect 8573 12835 8631 12841
rect 8573 12832 8585 12835
rect 8444 12804 8585 12832
rect 8444 12792 8450 12804
rect 8573 12801 8585 12804
rect 8619 12801 8631 12835
rect 8754 12832 8760 12844
rect 8715 12804 8760 12832
rect 8573 12795 8631 12801
rect 8754 12792 8760 12804
rect 8812 12792 8818 12844
rect 9493 12835 9551 12841
rect 9493 12801 9505 12835
rect 9539 12832 9551 12835
rect 9674 12832 9680 12844
rect 9539 12804 9680 12832
rect 9539 12801 9551 12804
rect 9493 12795 9551 12801
rect 9674 12792 9680 12804
rect 9732 12792 9738 12844
rect 9766 12792 9772 12844
rect 9824 12832 9830 12844
rect 10229 12835 10287 12841
rect 9824 12804 9869 12832
rect 9824 12792 9830 12804
rect 10229 12801 10241 12835
rect 10275 12832 10287 12835
rect 10778 12832 10784 12844
rect 10275 12804 10784 12832
rect 10275 12801 10287 12804
rect 10229 12795 10287 12801
rect 10778 12792 10784 12804
rect 10836 12832 10842 12844
rect 11624 12832 11652 12872
rect 14277 12869 14289 12872
rect 14323 12869 14335 12903
rect 14277 12863 14335 12869
rect 15004 12903 15062 12909
rect 15004 12869 15016 12903
rect 15050 12900 15062 12903
rect 15562 12900 15568 12912
rect 15050 12872 15568 12900
rect 15050 12869 15062 12872
rect 15004 12863 15062 12869
rect 15562 12860 15568 12872
rect 15620 12860 15626 12912
rect 16574 12860 16580 12912
rect 16632 12900 16638 12912
rect 18598 12900 18604 12912
rect 16632 12872 17080 12900
rect 16632 12860 16638 12872
rect 10836 12804 11652 12832
rect 11701 12835 11759 12841
rect 10836 12792 10842 12804
rect 11701 12801 11713 12835
rect 11747 12832 11759 12835
rect 12342 12832 12348 12844
rect 11747 12804 12348 12832
rect 11747 12801 11759 12804
rect 11701 12795 11759 12801
rect 12342 12792 12348 12804
rect 12400 12792 12406 12844
rect 12526 12832 12532 12844
rect 12487 12804 12532 12832
rect 12526 12792 12532 12804
rect 12584 12792 12590 12844
rect 12618 12792 12624 12844
rect 12676 12832 12682 12844
rect 12713 12835 12771 12841
rect 12713 12832 12725 12835
rect 12676 12804 12725 12832
rect 12676 12792 12682 12804
rect 12713 12801 12725 12804
rect 12759 12832 12771 12835
rect 13262 12832 13268 12844
rect 12759 12804 13268 12832
rect 12759 12801 12771 12804
rect 12713 12795 12771 12801
rect 13262 12792 13268 12804
rect 13320 12792 13326 12844
rect 13906 12832 13912 12844
rect 13867 12804 13912 12832
rect 13906 12792 13912 12804
rect 13964 12792 13970 12844
rect 14090 12832 14096 12844
rect 14051 12804 14096 12832
rect 14090 12792 14096 12804
rect 14148 12832 14154 12844
rect 14550 12832 14556 12844
rect 14148 12804 14556 12832
rect 14148 12792 14154 12804
rect 14550 12792 14556 12804
rect 14608 12792 14614 12844
rect 14734 12832 14740 12844
rect 14695 12804 14740 12832
rect 14734 12792 14740 12804
rect 14792 12792 14798 12844
rect 16758 12832 16764 12844
rect 16719 12804 16764 12832
rect 16758 12792 16764 12804
rect 16816 12792 16822 12844
rect 17052 12841 17080 12872
rect 17420 12872 18604 12900
rect 16945 12835 17003 12841
rect 16945 12801 16957 12835
rect 16991 12801 17003 12835
rect 16945 12795 17003 12801
rect 17037 12835 17095 12841
rect 17037 12801 17049 12835
rect 17083 12801 17095 12835
rect 17037 12795 17095 12801
rect 3970 12724 3976 12776
rect 4028 12764 4034 12776
rect 5353 12767 5411 12773
rect 5353 12764 5365 12767
rect 4028 12736 5365 12764
rect 4028 12724 4034 12736
rect 5353 12733 5365 12736
rect 5399 12764 5411 12767
rect 5626 12764 5632 12776
rect 5399 12736 5632 12764
rect 5399 12733 5411 12736
rect 5353 12727 5411 12733
rect 5626 12724 5632 12736
rect 5684 12764 5690 12776
rect 6546 12764 6552 12776
rect 5684 12736 6552 12764
rect 5684 12724 5690 12736
rect 6546 12724 6552 12736
rect 6604 12764 6610 12776
rect 6641 12767 6699 12773
rect 6641 12764 6653 12767
rect 6604 12736 6653 12764
rect 6604 12724 6610 12736
rect 6641 12733 6653 12736
rect 6687 12733 6699 12767
rect 6641 12727 6699 12733
rect 7653 12767 7711 12773
rect 7653 12733 7665 12767
rect 7699 12764 7711 12767
rect 8294 12764 8300 12776
rect 7699 12736 8300 12764
rect 7699 12733 7711 12736
rect 7653 12727 7711 12733
rect 8294 12724 8300 12736
rect 8352 12724 8358 12776
rect 10137 12767 10195 12773
rect 10137 12733 10149 12767
rect 10183 12764 10195 12767
rect 11882 12764 11888 12776
rect 10183 12736 11888 12764
rect 10183 12733 10195 12736
rect 10137 12727 10195 12733
rect 11882 12724 11888 12736
rect 11940 12724 11946 12776
rect 11977 12767 12035 12773
rect 11977 12733 11989 12767
rect 12023 12764 12035 12767
rect 13170 12764 13176 12776
rect 12023 12736 13176 12764
rect 12023 12733 12035 12736
rect 11977 12727 12035 12733
rect 13170 12724 13176 12736
rect 13228 12724 13234 12776
rect 16022 12724 16028 12776
rect 16080 12764 16086 12776
rect 16482 12764 16488 12776
rect 16080 12736 16488 12764
rect 16080 12724 16086 12736
rect 16482 12724 16488 12736
rect 16540 12724 16546 12776
rect 16960 12764 16988 12795
rect 17420 12764 17448 12872
rect 18598 12860 18604 12872
rect 18656 12860 18662 12912
rect 18785 12903 18843 12909
rect 18785 12869 18797 12903
rect 18831 12900 18843 12903
rect 19150 12900 19156 12912
rect 18831 12872 19156 12900
rect 18831 12869 18843 12872
rect 18785 12863 18843 12869
rect 19150 12860 19156 12872
rect 19208 12860 19214 12912
rect 19429 12903 19487 12909
rect 19429 12869 19441 12903
rect 19475 12900 19487 12903
rect 19886 12900 19892 12912
rect 19475 12872 19892 12900
rect 19475 12869 19487 12872
rect 19429 12863 19487 12869
rect 19886 12860 19892 12872
rect 19944 12860 19950 12912
rect 22370 12900 22376 12912
rect 20364 12872 22376 12900
rect 17681 12835 17739 12841
rect 17681 12801 17693 12835
rect 17727 12832 17739 12835
rect 17862 12832 17868 12844
rect 17727 12804 17868 12832
rect 17727 12801 17739 12804
rect 17681 12795 17739 12801
rect 17862 12792 17868 12804
rect 17920 12792 17926 12844
rect 17957 12835 18015 12841
rect 17957 12801 17969 12835
rect 18003 12801 18015 12835
rect 18138 12832 18144 12844
rect 18099 12804 18144 12832
rect 17957 12795 18015 12801
rect 16960 12736 17448 12764
rect 17494 12724 17500 12776
rect 17552 12764 17558 12776
rect 17972 12764 18000 12795
rect 18138 12792 18144 12804
rect 18196 12792 18202 12844
rect 19613 12835 19671 12841
rect 19613 12801 19625 12835
rect 19659 12801 19671 12835
rect 20364 12832 20392 12872
rect 22370 12860 22376 12872
rect 22428 12860 22434 12912
rect 24486 12860 24492 12912
rect 24544 12900 24550 12912
rect 24544 12872 25176 12900
rect 24544 12860 24550 12872
rect 20530 12832 20536 12844
rect 19613 12795 19671 12801
rect 19720 12804 20392 12832
rect 20491 12804 20536 12832
rect 17552 12736 18000 12764
rect 17552 12724 17558 12736
rect 2332 12668 3924 12696
rect 4157 12699 4215 12705
rect 4157 12665 4169 12699
rect 4203 12696 4215 12699
rect 16114 12696 16120 12708
rect 4203 12668 13492 12696
rect 16075 12668 16120 12696
rect 4203 12665 4215 12668
rect 4157 12659 4215 12665
rect 2222 12588 2228 12640
rect 2280 12628 2286 12640
rect 3237 12631 3295 12637
rect 3237 12628 3249 12631
rect 2280 12600 3249 12628
rect 2280 12588 2286 12600
rect 3237 12597 3249 12600
rect 3283 12597 3295 12631
rect 3602 12628 3608 12640
rect 3563 12600 3608 12628
rect 3237 12591 3295 12597
rect 3602 12588 3608 12600
rect 3660 12588 3666 12640
rect 5166 12588 5172 12640
rect 5224 12628 5230 12640
rect 7650 12628 7656 12640
rect 5224 12600 7656 12628
rect 5224 12588 5230 12600
rect 7650 12588 7656 12600
rect 7708 12588 7714 12640
rect 9214 12588 9220 12640
rect 9272 12628 9278 12640
rect 9309 12631 9367 12637
rect 9309 12628 9321 12631
rect 9272 12600 9321 12628
rect 9272 12588 9278 12600
rect 9309 12597 9321 12600
rect 9355 12597 9367 12631
rect 9309 12591 9367 12597
rect 9677 12631 9735 12637
rect 9677 12597 9689 12631
rect 9723 12628 9735 12631
rect 10137 12631 10195 12637
rect 10137 12628 10149 12631
rect 9723 12600 10149 12628
rect 9723 12597 9735 12600
rect 9677 12591 9735 12597
rect 10137 12597 10149 12600
rect 10183 12597 10195 12631
rect 10410 12628 10416 12640
rect 10371 12600 10416 12628
rect 10137 12591 10195 12597
rect 10410 12588 10416 12600
rect 10468 12588 10474 12640
rect 11330 12588 11336 12640
rect 11388 12628 11394 12640
rect 11517 12631 11575 12637
rect 11517 12628 11529 12631
rect 11388 12600 11529 12628
rect 11388 12588 11394 12600
rect 11517 12597 11529 12600
rect 11563 12597 11575 12631
rect 13354 12628 13360 12640
rect 13315 12600 13360 12628
rect 11517 12591 11575 12597
rect 13354 12588 13360 12600
rect 13412 12588 13418 12640
rect 13464 12628 13492 12668
rect 16114 12656 16120 12668
rect 16172 12656 16178 12708
rect 16761 12699 16819 12705
rect 16761 12665 16773 12699
rect 16807 12696 16819 12699
rect 19628 12696 19656 12795
rect 16807 12668 18092 12696
rect 16807 12665 16819 12668
rect 16761 12659 16819 12665
rect 16942 12628 16948 12640
rect 13464 12600 16948 12628
rect 16942 12588 16948 12600
rect 17000 12588 17006 12640
rect 17034 12588 17040 12640
rect 17092 12628 17098 12640
rect 17497 12631 17555 12637
rect 17497 12628 17509 12631
rect 17092 12600 17509 12628
rect 17092 12588 17098 12600
rect 17497 12597 17509 12600
rect 17543 12597 17555 12631
rect 18064 12628 18092 12668
rect 18432 12668 19656 12696
rect 18432 12628 18460 12668
rect 18064 12600 18460 12628
rect 18877 12631 18935 12637
rect 17497 12591 17555 12597
rect 18877 12597 18889 12631
rect 18923 12628 18935 12631
rect 19720 12628 19748 12804
rect 20530 12792 20536 12804
rect 20588 12792 20594 12844
rect 21910 12792 21916 12844
rect 21968 12832 21974 12844
rect 22005 12835 22063 12841
rect 22005 12832 22017 12835
rect 21968 12804 22017 12832
rect 21968 12792 21974 12804
rect 22005 12801 22017 12804
rect 22051 12801 22063 12835
rect 22005 12795 22063 12801
rect 23290 12792 23296 12844
rect 23348 12832 23354 12844
rect 23457 12835 23515 12841
rect 23457 12832 23469 12835
rect 23348 12804 23469 12832
rect 23348 12792 23354 12804
rect 23457 12801 23469 12804
rect 23503 12801 23515 12835
rect 25038 12832 25044 12844
rect 24999 12804 25044 12832
rect 23457 12795 23515 12801
rect 25038 12792 25044 12804
rect 25096 12792 25102 12844
rect 25148 12832 25176 12872
rect 25498 12860 25504 12912
rect 25556 12900 25562 12912
rect 27706 12900 27712 12912
rect 25556 12872 26280 12900
rect 25556 12860 25562 12872
rect 25682 12832 25688 12844
rect 25148 12804 25688 12832
rect 25682 12792 25688 12804
rect 25740 12792 25746 12844
rect 25866 12792 25872 12844
rect 25924 12832 25930 12844
rect 26252 12841 26280 12872
rect 26436 12872 27712 12900
rect 26436 12841 26464 12872
rect 27706 12860 27712 12872
rect 27764 12860 27770 12912
rect 28994 12900 29000 12912
rect 28276 12872 29000 12900
rect 25961 12835 26019 12841
rect 25961 12832 25973 12835
rect 25924 12804 25973 12832
rect 25924 12792 25930 12804
rect 25961 12801 25973 12804
rect 26007 12801 26019 12835
rect 25961 12795 26019 12801
rect 26237 12835 26295 12841
rect 26237 12801 26249 12835
rect 26283 12801 26295 12835
rect 26237 12795 26295 12801
rect 26421 12835 26479 12841
rect 26421 12801 26433 12835
rect 26467 12801 26479 12835
rect 26421 12795 26479 12801
rect 27157 12835 27215 12841
rect 27157 12801 27169 12835
rect 27203 12801 27215 12835
rect 27430 12832 27436 12844
rect 27391 12804 27436 12832
rect 27157 12795 27215 12801
rect 19889 12767 19947 12773
rect 19889 12733 19901 12767
rect 19935 12764 19947 12767
rect 20254 12764 20260 12776
rect 19935 12736 20260 12764
rect 19935 12733 19947 12736
rect 19889 12727 19947 12733
rect 20254 12724 20260 12736
rect 20312 12724 20318 12776
rect 20438 12724 20444 12776
rect 20496 12764 20502 12776
rect 20809 12767 20867 12773
rect 20809 12764 20821 12767
rect 20496 12736 20821 12764
rect 20496 12724 20502 12736
rect 20809 12733 20821 12736
rect 20855 12733 20867 12767
rect 20809 12727 20867 12733
rect 21542 12724 21548 12776
rect 21600 12764 21606 12776
rect 21821 12767 21879 12773
rect 21821 12764 21833 12767
rect 21600 12736 21833 12764
rect 21600 12724 21606 12736
rect 21821 12733 21833 12736
rect 21867 12733 21879 12767
rect 21821 12727 21879 12733
rect 23201 12767 23259 12773
rect 23201 12733 23213 12767
rect 23247 12733 23259 12767
rect 24946 12764 24952 12776
rect 23201 12727 23259 12733
rect 24596 12736 24952 12764
rect 20717 12699 20775 12705
rect 20717 12696 20729 12699
rect 19812 12668 20729 12696
rect 19812 12640 19840 12668
rect 20717 12665 20729 12668
rect 20763 12665 20775 12699
rect 20717 12659 20775 12665
rect 21358 12656 21364 12708
rect 21416 12696 21422 12708
rect 23216 12696 23244 12727
rect 21416 12668 23244 12696
rect 21416 12656 21422 12668
rect 18923 12600 19748 12628
rect 18923 12597 18935 12600
rect 18877 12591 18935 12597
rect 19794 12588 19800 12640
rect 19852 12628 19858 12640
rect 20346 12628 20352 12640
rect 19852 12600 19897 12628
rect 20307 12600 20352 12628
rect 19852 12588 19858 12600
rect 20346 12588 20352 12600
rect 20404 12588 20410 12640
rect 20806 12588 20812 12640
rect 20864 12628 20870 12640
rect 21376 12628 21404 12656
rect 20864 12600 21404 12628
rect 22189 12631 22247 12637
rect 20864 12588 20870 12600
rect 22189 12597 22201 12631
rect 22235 12628 22247 12631
rect 22554 12628 22560 12640
rect 22235 12600 22560 12628
rect 22235 12597 22247 12600
rect 22189 12591 22247 12597
rect 22554 12588 22560 12600
rect 22612 12588 22618 12640
rect 23934 12588 23940 12640
rect 23992 12628 23998 12640
rect 24596 12637 24624 12736
rect 24946 12724 24952 12736
rect 25004 12764 25010 12776
rect 25317 12767 25375 12773
rect 25317 12764 25329 12767
rect 25004 12736 25329 12764
rect 25004 12724 25010 12736
rect 25317 12733 25329 12736
rect 25363 12733 25375 12767
rect 25976 12764 26004 12795
rect 26142 12764 26148 12776
rect 25976 12736 26148 12764
rect 25317 12727 25375 12733
rect 26142 12724 26148 12736
rect 26200 12764 26206 12776
rect 27172 12764 27200 12795
rect 27430 12792 27436 12804
rect 27488 12792 27494 12844
rect 27614 12832 27620 12844
rect 27575 12804 27620 12832
rect 27614 12792 27620 12804
rect 27672 12792 27678 12844
rect 28276 12841 28304 12872
rect 28994 12860 29000 12872
rect 29052 12860 29058 12912
rect 28261 12835 28319 12841
rect 28261 12801 28273 12835
rect 28307 12801 28319 12835
rect 28261 12795 28319 12801
rect 28528 12835 28586 12841
rect 28528 12801 28540 12835
rect 28574 12832 28586 12835
rect 29546 12832 29552 12844
rect 28574 12804 29552 12832
rect 28574 12801 28586 12804
rect 28528 12795 28586 12801
rect 29546 12792 29552 12804
rect 29604 12792 29610 12844
rect 30282 12792 30288 12844
rect 30340 12832 30346 12844
rect 30561 12835 30619 12841
rect 30561 12832 30573 12835
rect 30340 12804 30573 12832
rect 30340 12792 30346 12804
rect 30561 12801 30573 12804
rect 30607 12801 30619 12835
rect 30561 12795 30619 12801
rect 30837 12835 30895 12841
rect 30837 12801 30849 12835
rect 30883 12832 30895 12835
rect 30926 12832 30932 12844
rect 30883 12804 30932 12832
rect 30883 12801 30895 12804
rect 30837 12795 30895 12801
rect 30926 12792 30932 12804
rect 30984 12832 30990 12844
rect 31202 12832 31208 12844
rect 30984 12804 31208 12832
rect 30984 12792 30990 12804
rect 31202 12792 31208 12804
rect 31260 12792 31266 12844
rect 26200 12736 27200 12764
rect 26200 12724 26206 12736
rect 29914 12724 29920 12776
rect 29972 12764 29978 12776
rect 30745 12767 30803 12773
rect 30745 12764 30757 12767
rect 29972 12736 30757 12764
rect 29972 12724 29978 12736
rect 30745 12733 30757 12736
rect 30791 12733 30803 12767
rect 30745 12727 30803 12733
rect 25133 12699 25191 12705
rect 25133 12665 25145 12699
rect 25179 12696 25191 12699
rect 27338 12696 27344 12708
rect 25179 12668 27344 12696
rect 25179 12665 25191 12668
rect 25133 12659 25191 12665
rect 27338 12656 27344 12668
rect 27396 12656 27402 12708
rect 24581 12631 24639 12637
rect 24581 12628 24593 12631
rect 23992 12600 24593 12628
rect 23992 12588 23998 12600
rect 24581 12597 24593 12600
rect 24627 12597 24639 12631
rect 24581 12591 24639 12597
rect 25222 12588 25228 12640
rect 25280 12628 25286 12640
rect 25777 12631 25835 12637
rect 25280 12600 25325 12628
rect 25280 12588 25286 12600
rect 25777 12597 25789 12631
rect 25823 12628 25835 12631
rect 25958 12628 25964 12640
rect 25823 12600 25964 12628
rect 25823 12597 25835 12600
rect 25777 12591 25835 12597
rect 25958 12588 25964 12600
rect 26016 12588 26022 12640
rect 30190 12588 30196 12640
rect 30248 12628 30254 12640
rect 30377 12631 30435 12637
rect 30377 12628 30389 12631
rect 30248 12600 30389 12628
rect 30248 12588 30254 12600
rect 30377 12597 30389 12600
rect 30423 12597 30435 12631
rect 30377 12591 30435 12597
rect 1104 12538 32016 12560
rect 1104 12486 2136 12538
rect 2188 12486 12440 12538
rect 12492 12486 22744 12538
rect 22796 12486 32016 12538
rect 1104 12464 32016 12486
rect 2777 12427 2835 12433
rect 2777 12393 2789 12427
rect 2823 12424 2835 12427
rect 2958 12424 2964 12436
rect 2823 12396 2964 12424
rect 2823 12393 2835 12396
rect 2777 12387 2835 12393
rect 2958 12384 2964 12396
rect 3016 12384 3022 12436
rect 3878 12384 3884 12436
rect 3936 12424 3942 12436
rect 5902 12424 5908 12436
rect 3936 12396 5764 12424
rect 5863 12396 5908 12424
rect 3936 12384 3942 12396
rect 3050 12248 3056 12300
rect 3108 12288 3114 12300
rect 3602 12288 3608 12300
rect 3108 12260 3608 12288
rect 3108 12248 3114 12260
rect 3602 12248 3608 12260
rect 3660 12288 3666 12300
rect 4065 12291 4123 12297
rect 4065 12288 4077 12291
rect 3660 12260 4077 12288
rect 3660 12248 3666 12260
rect 4065 12257 4077 12260
rect 4111 12257 4123 12291
rect 5736 12288 5764 12396
rect 5902 12384 5908 12396
rect 5960 12384 5966 12436
rect 6178 12384 6184 12436
rect 6236 12424 6242 12436
rect 6733 12427 6791 12433
rect 6733 12424 6745 12427
rect 6236 12396 6745 12424
rect 6236 12384 6242 12396
rect 6733 12393 6745 12396
rect 6779 12393 6791 12427
rect 6733 12387 6791 12393
rect 7650 12384 7656 12436
rect 7708 12424 7714 12436
rect 8662 12424 8668 12436
rect 7708 12396 8668 12424
rect 7708 12384 7714 12396
rect 8662 12384 8668 12396
rect 8720 12384 8726 12436
rect 9122 12384 9128 12436
rect 9180 12424 9186 12436
rect 13262 12424 13268 12436
rect 9180 12396 13268 12424
rect 9180 12384 9186 12396
rect 13262 12384 13268 12396
rect 13320 12384 13326 12436
rect 13449 12427 13507 12433
rect 13449 12393 13461 12427
rect 13495 12424 13507 12427
rect 13722 12424 13728 12436
rect 13495 12396 13728 12424
rect 13495 12393 13507 12396
rect 13449 12387 13507 12393
rect 13722 12384 13728 12396
rect 13780 12384 13786 12436
rect 14108 12396 15194 12424
rect 6454 12316 6460 12368
rect 6512 12356 6518 12368
rect 6638 12356 6644 12368
rect 6512 12328 6644 12356
rect 6512 12316 6518 12328
rect 6638 12316 6644 12328
rect 6696 12316 6702 12368
rect 7374 12316 7380 12368
rect 7432 12356 7438 12368
rect 7432 12328 8616 12356
rect 7432 12316 7438 12328
rect 8588 12300 8616 12328
rect 11514 12316 11520 12368
rect 11572 12356 11578 12368
rect 14108 12356 14136 12396
rect 11572 12328 14136 12356
rect 15166 12356 15194 12396
rect 15378 12384 15384 12436
rect 15436 12424 15442 12436
rect 17681 12427 17739 12433
rect 15436 12396 17632 12424
rect 15436 12384 15442 12396
rect 16298 12356 16304 12368
rect 15166 12328 16304 12356
rect 11572 12316 11578 12328
rect 16298 12316 16304 12328
rect 16356 12316 16362 12368
rect 6270 12288 6276 12300
rect 5736 12260 6276 12288
rect 4065 12251 4123 12257
rect 6270 12248 6276 12260
rect 6328 12288 6334 12300
rect 8297 12291 8355 12297
rect 6328 12260 8064 12288
rect 6328 12248 6334 12260
rect 1394 12220 1400 12232
rect 1307 12192 1400 12220
rect 1394 12180 1400 12192
rect 1452 12220 1458 12232
rect 4430 12220 4436 12232
rect 1452 12192 4436 12220
rect 1452 12180 1458 12192
rect 4430 12180 4436 12192
rect 4488 12220 4494 12232
rect 4525 12223 4583 12229
rect 4525 12220 4537 12223
rect 4488 12192 4537 12220
rect 4488 12180 4494 12192
rect 4525 12189 4537 12192
rect 4571 12189 4583 12223
rect 6454 12220 6460 12232
rect 6415 12192 6460 12220
rect 4525 12183 4583 12189
rect 6454 12180 6460 12192
rect 6512 12180 6518 12232
rect 6549 12223 6607 12229
rect 6549 12189 6561 12223
rect 6595 12220 6607 12223
rect 6638 12220 6644 12232
rect 6595 12192 6644 12220
rect 6595 12189 6607 12192
rect 6549 12183 6607 12189
rect 6638 12180 6644 12192
rect 6696 12180 6702 12232
rect 7466 12180 7472 12232
rect 7524 12220 7530 12232
rect 7834 12220 7840 12232
rect 7524 12192 7840 12220
rect 7524 12180 7530 12192
rect 7834 12180 7840 12192
rect 7892 12180 7898 12232
rect 8036 12229 8064 12260
rect 8297 12257 8309 12291
rect 8343 12257 8355 12291
rect 8297 12251 8355 12257
rect 8021 12223 8079 12229
rect 8021 12189 8033 12223
rect 8067 12189 8079 12223
rect 8021 12183 8079 12189
rect 1664 12155 1722 12161
rect 1664 12121 1676 12155
rect 1710 12152 1722 12155
rect 2222 12152 2228 12164
rect 1710 12124 2228 12152
rect 1710 12121 1722 12124
rect 1664 12115 1722 12121
rect 2222 12112 2228 12124
rect 2280 12112 2286 12164
rect 2314 12112 2320 12164
rect 2372 12152 2378 12164
rect 2372 12124 2774 12152
rect 2372 12112 2378 12124
rect 2746 12084 2774 12124
rect 3786 12112 3792 12164
rect 3844 12152 3850 12164
rect 3881 12155 3939 12161
rect 3881 12152 3893 12155
rect 3844 12124 3893 12152
rect 3844 12112 3850 12124
rect 3881 12121 3893 12124
rect 3927 12121 3939 12155
rect 3881 12115 3939 12121
rect 4792 12155 4850 12161
rect 4792 12121 4804 12155
rect 4838 12152 4850 12155
rect 4890 12152 4896 12164
rect 4838 12124 4896 12152
rect 4838 12121 4850 12124
rect 4792 12115 4850 12121
rect 4890 12112 4896 12124
rect 4948 12112 4954 12164
rect 5350 12112 5356 12164
rect 5408 12152 5414 12164
rect 8113 12155 8171 12161
rect 8113 12152 8125 12155
rect 5408 12124 8125 12152
rect 5408 12112 5414 12124
rect 8113 12121 8125 12124
rect 8159 12121 8171 12155
rect 8312 12152 8340 12251
rect 8570 12248 8576 12300
rect 8628 12248 8634 12300
rect 8938 12288 8944 12300
rect 8899 12260 8944 12288
rect 8938 12248 8944 12260
rect 8996 12248 9002 12300
rect 13630 12288 13636 12300
rect 13372 12260 13636 12288
rect 9214 12229 9220 12232
rect 9208 12183 9220 12229
rect 9272 12220 9278 12232
rect 10778 12220 10784 12232
rect 9272 12192 9308 12220
rect 10739 12192 10784 12220
rect 9214 12180 9220 12183
rect 9272 12180 9278 12192
rect 10778 12180 10784 12192
rect 10836 12180 10842 12232
rect 11054 12220 11060 12232
rect 11015 12192 11060 12220
rect 11054 12180 11060 12192
rect 11112 12180 11118 12232
rect 12618 12180 12624 12232
rect 12676 12220 12682 12232
rect 13372 12229 13400 12260
rect 13630 12248 13636 12260
rect 13688 12248 13694 12300
rect 15102 12248 15108 12300
rect 15160 12288 15166 12300
rect 16022 12288 16028 12300
rect 15160 12260 16028 12288
rect 15160 12248 15166 12260
rect 16022 12248 16028 12260
rect 16080 12248 16086 12300
rect 12713 12223 12771 12229
rect 12713 12220 12725 12223
rect 12676 12192 12725 12220
rect 12676 12180 12682 12192
rect 12713 12189 12725 12192
rect 12759 12189 12771 12223
rect 12713 12183 12771 12189
rect 13357 12223 13415 12229
rect 13357 12189 13369 12223
rect 13403 12189 13415 12223
rect 13538 12220 13544 12232
rect 13499 12192 13544 12220
rect 13357 12183 13415 12189
rect 13538 12180 13544 12192
rect 13596 12180 13602 12232
rect 13814 12180 13820 12232
rect 13872 12220 13878 12232
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 13872 12192 14105 12220
rect 13872 12180 13878 12192
rect 14093 12189 14105 12192
rect 14139 12220 14151 12223
rect 14734 12220 14740 12232
rect 14139 12192 14740 12220
rect 14139 12189 14151 12192
rect 14093 12183 14151 12189
rect 14734 12180 14740 12192
rect 14792 12220 14798 12232
rect 16301 12223 16359 12229
rect 16301 12220 16313 12223
rect 14792 12192 16313 12220
rect 14792 12180 14798 12192
rect 16301 12189 16313 12192
rect 16347 12189 16359 12223
rect 17604 12220 17632 12396
rect 17681 12393 17693 12427
rect 17727 12424 17739 12427
rect 17954 12424 17960 12436
rect 17727 12396 17960 12424
rect 17727 12393 17739 12396
rect 17681 12387 17739 12393
rect 17954 12384 17960 12396
rect 18012 12424 18018 12436
rect 18138 12424 18144 12436
rect 18012 12396 18144 12424
rect 18012 12384 18018 12396
rect 18138 12384 18144 12396
rect 18196 12384 18202 12436
rect 19334 12384 19340 12436
rect 19392 12424 19398 12436
rect 19613 12427 19671 12433
rect 19392 12396 19564 12424
rect 19392 12384 19398 12396
rect 17770 12316 17776 12368
rect 17828 12356 17834 12368
rect 18966 12356 18972 12368
rect 17828 12328 18972 12356
rect 17828 12316 17834 12328
rect 18966 12316 18972 12328
rect 19024 12316 19030 12368
rect 19536 12356 19564 12396
rect 19613 12393 19625 12427
rect 19659 12424 19671 12427
rect 20530 12424 20536 12436
rect 19659 12396 20536 12424
rect 19659 12393 19671 12396
rect 19613 12387 19671 12393
rect 20530 12384 20536 12396
rect 20588 12384 20594 12436
rect 20898 12384 20904 12436
rect 20956 12424 20962 12436
rect 21634 12424 21640 12436
rect 20956 12396 21640 12424
rect 20956 12384 20962 12396
rect 21634 12384 21640 12396
rect 21692 12384 21698 12436
rect 23290 12384 23296 12436
rect 23348 12424 23354 12436
rect 23385 12427 23443 12433
rect 23385 12424 23397 12427
rect 23348 12396 23397 12424
rect 23348 12384 23354 12396
rect 23385 12393 23397 12396
rect 23431 12393 23443 12427
rect 23385 12387 23443 12393
rect 23474 12384 23480 12436
rect 23532 12424 23538 12436
rect 26145 12427 26203 12433
rect 26145 12424 26157 12427
rect 23532 12396 26157 12424
rect 23532 12384 23538 12396
rect 26145 12393 26157 12396
rect 26191 12424 26203 12427
rect 26510 12424 26516 12436
rect 26191 12396 26516 12424
rect 26191 12393 26203 12396
rect 26145 12387 26203 12393
rect 26510 12384 26516 12396
rect 26568 12384 26574 12436
rect 26712 12396 27660 12424
rect 20714 12356 20720 12368
rect 19536 12328 20720 12356
rect 20714 12316 20720 12328
rect 20772 12316 20778 12368
rect 20993 12359 21051 12365
rect 20993 12325 21005 12359
rect 21039 12356 21051 12359
rect 23753 12359 23811 12365
rect 23753 12356 23765 12359
rect 21039 12328 21956 12356
rect 21039 12325 21051 12328
rect 20993 12319 21051 12325
rect 18693 12291 18751 12297
rect 18693 12257 18705 12291
rect 18739 12288 18751 12291
rect 21928 12288 21956 12328
rect 23676 12328 23765 12356
rect 23676 12300 23704 12328
rect 23753 12325 23765 12328
rect 23799 12325 23811 12359
rect 23753 12319 23811 12325
rect 24118 12316 24124 12368
rect 24176 12356 24182 12368
rect 26712 12356 26740 12396
rect 24176 12328 26740 12356
rect 27632 12356 27660 12396
rect 27706 12384 27712 12436
rect 27764 12424 27770 12436
rect 28074 12424 28080 12436
rect 27764 12396 28080 12424
rect 27764 12384 27770 12396
rect 28074 12384 28080 12396
rect 28132 12384 28138 12436
rect 28718 12424 28724 12436
rect 28679 12396 28724 12424
rect 28718 12384 28724 12396
rect 28776 12384 28782 12436
rect 31018 12384 31024 12436
rect 31076 12424 31082 12436
rect 31297 12427 31355 12433
rect 31297 12424 31309 12427
rect 31076 12396 31309 12424
rect 31076 12384 31082 12396
rect 31297 12393 31309 12396
rect 31343 12393 31355 12427
rect 31297 12387 31355 12393
rect 27632 12328 28212 12356
rect 24176 12316 24182 12328
rect 23106 12288 23112 12300
rect 18739 12260 21864 12288
rect 21928 12260 23112 12288
rect 18739 12257 18751 12260
rect 18693 12251 18751 12257
rect 18509 12223 18567 12229
rect 18509 12220 18521 12223
rect 17604 12192 18521 12220
rect 16301 12183 16359 12189
rect 18509 12189 18521 12192
rect 18555 12189 18567 12223
rect 18509 12183 18567 12189
rect 8312 12124 9444 12152
rect 8113 12115 8171 12121
rect 9416 12096 9444 12124
rect 11238 12112 11244 12164
rect 11296 12152 11302 12164
rect 14338 12155 14396 12161
rect 14338 12152 14350 12155
rect 11296 12124 14350 12152
rect 11296 12112 11302 12124
rect 14338 12121 14350 12124
rect 14384 12121 14396 12155
rect 14338 12115 14396 12121
rect 16568 12155 16626 12161
rect 16568 12121 16580 12155
rect 16614 12152 16626 12155
rect 16850 12152 16856 12164
rect 16614 12124 16856 12152
rect 16614 12121 16626 12124
rect 16568 12115 16626 12121
rect 16850 12112 16856 12124
rect 16908 12112 16914 12164
rect 16942 12112 16948 12164
rect 17000 12152 17006 12164
rect 18322 12152 18328 12164
rect 17000 12124 18328 12152
rect 17000 12112 17006 12124
rect 18322 12112 18328 12124
rect 18380 12112 18386 12164
rect 3694 12084 3700 12096
rect 2746 12056 3700 12084
rect 3694 12044 3700 12056
rect 3752 12044 3758 12096
rect 4706 12044 4712 12096
rect 4764 12084 4770 12096
rect 5718 12084 5724 12096
rect 4764 12056 5724 12084
rect 4764 12044 4770 12056
rect 5718 12044 5724 12056
rect 5776 12044 5782 12096
rect 7006 12044 7012 12096
rect 7064 12084 7070 12096
rect 7466 12084 7472 12096
rect 7064 12056 7472 12084
rect 7064 12044 7070 12056
rect 7466 12044 7472 12056
rect 7524 12044 7530 12096
rect 7650 12084 7656 12096
rect 7611 12056 7656 12084
rect 7650 12044 7656 12056
rect 7708 12044 7714 12096
rect 7834 12044 7840 12096
rect 7892 12084 7898 12096
rect 8754 12084 8760 12096
rect 7892 12056 8760 12084
rect 7892 12044 7898 12056
rect 8754 12044 8760 12056
rect 8812 12044 8818 12096
rect 9398 12044 9404 12096
rect 9456 12084 9462 12096
rect 10321 12087 10379 12093
rect 10321 12084 10333 12087
rect 9456 12056 10333 12084
rect 9456 12044 9462 12056
rect 10321 12053 10333 12056
rect 10367 12053 10379 12087
rect 12802 12084 12808 12096
rect 12763 12056 12808 12084
rect 10321 12047 10379 12053
rect 12802 12044 12808 12056
rect 12860 12044 12866 12096
rect 14550 12044 14556 12096
rect 14608 12084 14614 12096
rect 15473 12087 15531 12093
rect 15473 12084 15485 12087
rect 14608 12056 15485 12084
rect 14608 12044 14614 12056
rect 15473 12053 15485 12056
rect 15519 12053 15531 12087
rect 15473 12047 15531 12053
rect 15930 12044 15936 12096
rect 15988 12084 15994 12096
rect 16758 12084 16764 12096
rect 15988 12056 16764 12084
rect 15988 12044 15994 12056
rect 16758 12044 16764 12056
rect 16816 12084 16822 12096
rect 18414 12084 18420 12096
rect 16816 12056 18420 12084
rect 16816 12044 16822 12056
rect 18414 12044 18420 12056
rect 18472 12044 18478 12096
rect 18524 12084 18552 12183
rect 19150 12180 19156 12232
rect 19208 12220 19214 12232
rect 19702 12220 19708 12232
rect 19208 12192 19708 12220
rect 19208 12180 19214 12192
rect 19702 12180 19708 12192
rect 19760 12220 19766 12232
rect 19797 12223 19855 12229
rect 19797 12220 19809 12223
rect 19760 12192 19809 12220
rect 19760 12180 19766 12192
rect 19797 12189 19809 12192
rect 19843 12189 19855 12223
rect 20070 12220 20076 12232
rect 20031 12192 20076 12220
rect 19797 12183 19855 12189
rect 20070 12180 20076 12192
rect 20128 12180 20134 12232
rect 20254 12180 20260 12232
rect 20312 12220 20318 12232
rect 20530 12220 20536 12232
rect 20312 12192 20536 12220
rect 20312 12180 20318 12192
rect 20530 12180 20536 12192
rect 20588 12180 20594 12232
rect 21450 12220 21456 12232
rect 21411 12192 21456 12220
rect 21450 12180 21456 12192
rect 21508 12180 21514 12232
rect 18966 12112 18972 12164
rect 19024 12152 19030 12164
rect 20088 12152 20116 12180
rect 20809 12155 20867 12161
rect 20809 12152 20821 12155
rect 19024 12124 20116 12152
rect 20640 12124 20821 12152
rect 19024 12112 19030 12124
rect 20640 12084 20668 12124
rect 20809 12121 20821 12124
rect 20855 12152 20867 12155
rect 21358 12152 21364 12164
rect 20855 12124 21364 12152
rect 20855 12121 20867 12124
rect 20809 12115 20867 12121
rect 21358 12112 21364 12124
rect 21416 12112 21422 12164
rect 21836 12152 21864 12260
rect 23106 12248 23112 12260
rect 23164 12288 23170 12300
rect 23474 12288 23480 12300
rect 23164 12260 23480 12288
rect 23164 12248 23170 12260
rect 23474 12248 23480 12260
rect 23532 12248 23538 12300
rect 23658 12248 23664 12300
rect 23716 12248 23722 12300
rect 23860 12260 25084 12288
rect 22554 12220 22560 12232
rect 22515 12192 22560 12220
rect 22554 12180 22560 12192
rect 22612 12180 22618 12232
rect 23566 12220 23572 12232
rect 23527 12192 23572 12220
rect 23566 12180 23572 12192
rect 23624 12180 23630 12232
rect 23860 12229 23888 12260
rect 25056 12232 25084 12260
rect 23845 12223 23903 12229
rect 23845 12189 23857 12223
rect 23891 12189 23903 12223
rect 24946 12220 24952 12232
rect 24907 12192 24952 12220
rect 23845 12183 23903 12189
rect 24946 12180 24952 12192
rect 25004 12180 25010 12232
rect 25038 12180 25044 12232
rect 25096 12220 25102 12232
rect 25133 12223 25191 12229
rect 25133 12220 25145 12223
rect 25096 12192 25145 12220
rect 25096 12180 25102 12192
rect 25133 12189 25145 12192
rect 25179 12189 25191 12223
rect 25133 12183 25191 12189
rect 25225 12223 25283 12229
rect 25225 12189 25237 12223
rect 25271 12189 25283 12223
rect 25958 12220 25964 12232
rect 25919 12192 25964 12220
rect 25225 12183 25283 12189
rect 23658 12152 23664 12164
rect 21836 12124 23664 12152
rect 23658 12112 23664 12124
rect 23716 12112 23722 12164
rect 24026 12112 24032 12164
rect 24084 12152 24090 12164
rect 25240 12152 25268 12183
rect 25958 12180 25964 12192
rect 26016 12180 26022 12232
rect 26237 12223 26295 12229
rect 26237 12189 26249 12223
rect 26283 12189 26295 12223
rect 26694 12220 26700 12232
rect 26655 12192 26700 12220
rect 26237 12183 26295 12189
rect 25406 12152 25412 12164
rect 24084 12124 25412 12152
rect 24084 12112 24090 12124
rect 25406 12112 25412 12124
rect 25464 12112 25470 12164
rect 26252 12152 26280 12183
rect 26694 12180 26700 12192
rect 26752 12180 26758 12232
rect 26970 12229 26976 12232
rect 26964 12183 26976 12229
rect 27028 12220 27034 12232
rect 27028 12192 27064 12220
rect 26970 12180 26976 12183
rect 27028 12180 27034 12192
rect 27614 12152 27620 12164
rect 26252 12124 27620 12152
rect 27614 12112 27620 12124
rect 27672 12152 27678 12164
rect 27982 12152 27988 12164
rect 27672 12124 27988 12152
rect 27672 12112 27678 12124
rect 27982 12112 27988 12124
rect 28040 12152 28046 12164
rect 28184 12152 28212 12328
rect 28994 12248 29000 12300
rect 29052 12288 29058 12300
rect 29917 12291 29975 12297
rect 29917 12288 29929 12291
rect 29052 12260 29929 12288
rect 29052 12248 29058 12260
rect 29917 12257 29929 12260
rect 29963 12257 29975 12291
rect 29917 12251 29975 12257
rect 30190 12229 30196 12232
rect 30184 12183 30196 12229
rect 30248 12220 30254 12232
rect 30248 12192 30284 12220
rect 30190 12180 30196 12183
rect 30248 12180 30254 12192
rect 28537 12155 28595 12161
rect 28537 12152 28549 12155
rect 28040 12124 28120 12152
rect 28184 12124 28549 12152
rect 28040 12112 28046 12124
rect 18524 12056 20668 12084
rect 22649 12087 22707 12093
rect 22649 12053 22661 12087
rect 22695 12084 22707 12087
rect 23382 12084 23388 12096
rect 22695 12056 23388 12084
rect 22695 12053 22707 12056
rect 22649 12047 22707 12053
rect 23382 12044 23388 12056
rect 23440 12044 23446 12096
rect 23566 12044 23572 12096
rect 23624 12084 23630 12096
rect 24302 12084 24308 12096
rect 23624 12056 24308 12084
rect 23624 12044 23630 12056
rect 24302 12044 24308 12056
rect 24360 12044 24366 12096
rect 24762 12084 24768 12096
rect 24723 12056 24768 12084
rect 24762 12044 24768 12056
rect 24820 12044 24826 12096
rect 25777 12087 25835 12093
rect 25777 12053 25789 12087
rect 25823 12084 25835 12087
rect 26786 12084 26792 12096
rect 25823 12056 26792 12084
rect 25823 12053 25835 12056
rect 25777 12047 25835 12053
rect 26786 12044 26792 12056
rect 26844 12044 26850 12096
rect 28092 12093 28120 12124
rect 28537 12121 28549 12124
rect 28583 12152 28595 12155
rect 30834 12152 30840 12164
rect 28583 12124 30840 12152
rect 28583 12121 28595 12124
rect 28537 12115 28595 12121
rect 30834 12112 30840 12124
rect 30892 12112 30898 12164
rect 28077 12087 28135 12093
rect 28077 12053 28089 12087
rect 28123 12053 28135 12087
rect 28077 12047 28135 12053
rect 28166 12044 28172 12096
rect 28224 12084 28230 12096
rect 28737 12087 28795 12093
rect 28737 12084 28749 12087
rect 28224 12056 28749 12084
rect 28224 12044 28230 12056
rect 28737 12053 28749 12056
rect 28783 12053 28795 12087
rect 28737 12047 28795 12053
rect 28905 12087 28963 12093
rect 28905 12053 28917 12087
rect 28951 12084 28963 12087
rect 30006 12084 30012 12096
rect 28951 12056 30012 12084
rect 28951 12053 28963 12056
rect 28905 12047 28963 12053
rect 30006 12044 30012 12056
rect 30064 12044 30070 12096
rect 1104 11994 32016 12016
rect 1104 11942 7288 11994
rect 7340 11942 17592 11994
rect 17644 11942 27896 11994
rect 27948 11942 32016 11994
rect 1104 11920 32016 11942
rect 2498 11840 2504 11892
rect 2556 11880 2562 11892
rect 6733 11883 6791 11889
rect 6733 11880 6745 11883
rect 2556 11852 6745 11880
rect 2556 11840 2562 11852
rect 6733 11849 6745 11852
rect 6779 11880 6791 11883
rect 7929 11883 7987 11889
rect 7929 11880 7941 11883
rect 6779 11852 7941 11880
rect 6779 11849 6791 11852
rect 6733 11843 6791 11849
rect 7929 11849 7941 11852
rect 7975 11849 7987 11883
rect 7929 11843 7987 11849
rect 9950 11840 9956 11892
rect 10008 11880 10014 11892
rect 10873 11883 10931 11889
rect 10873 11880 10885 11883
rect 10008 11852 10885 11880
rect 10008 11840 10014 11852
rect 10873 11849 10885 11852
rect 10919 11880 10931 11883
rect 11146 11880 11152 11892
rect 10919 11852 11152 11880
rect 10919 11849 10931 11852
rect 10873 11843 10931 11849
rect 11146 11840 11152 11852
rect 11204 11840 11210 11892
rect 13170 11880 13176 11892
rect 13131 11852 13176 11880
rect 13170 11840 13176 11852
rect 13228 11880 13234 11892
rect 14001 11883 14059 11889
rect 14001 11880 14013 11883
rect 13228 11852 14013 11880
rect 13228 11840 13234 11852
rect 14001 11849 14013 11852
rect 14047 11849 14059 11883
rect 14001 11843 14059 11849
rect 15473 11883 15531 11889
rect 15473 11849 15485 11883
rect 15519 11849 15531 11883
rect 15473 11843 15531 11849
rect 0 11812 800 11826
rect 1765 11815 1823 11821
rect 0 11784 888 11812
rect 0 11770 800 11784
rect 860 11608 888 11784
rect 1765 11781 1777 11815
rect 1811 11812 1823 11815
rect 2930 11815 2988 11821
rect 2930 11812 2942 11815
rect 1811 11784 2942 11812
rect 1811 11781 1823 11784
rect 1765 11775 1823 11781
rect 2930 11781 2942 11784
rect 2976 11781 2988 11815
rect 2930 11775 2988 11781
rect 3694 11772 3700 11824
rect 3752 11812 3758 11824
rect 6825 11815 6883 11821
rect 6825 11812 6837 11815
rect 3752 11784 6837 11812
rect 3752 11772 3758 11784
rect 6825 11781 6837 11784
rect 6871 11812 6883 11815
rect 8021 11815 8079 11821
rect 8021 11812 8033 11815
rect 6871 11784 8033 11812
rect 6871 11781 6883 11784
rect 6825 11775 6883 11781
rect 8021 11781 8033 11784
rect 8067 11781 8079 11815
rect 8021 11775 8079 11781
rect 10781 11815 10839 11821
rect 10781 11781 10793 11815
rect 10827 11812 10839 11815
rect 10827 11784 12204 11812
rect 10827 11781 10839 11784
rect 10781 11775 10839 11781
rect 1946 11744 1952 11756
rect 1907 11716 1952 11744
rect 1946 11704 1952 11716
rect 2004 11704 2010 11756
rect 4433 11747 4491 11753
rect 4433 11744 4445 11747
rect 2516 11716 4445 11744
rect 1578 11636 1584 11688
rect 1636 11676 1642 11688
rect 2225 11679 2283 11685
rect 2225 11676 2237 11679
rect 1636 11648 2237 11676
rect 1636 11636 1642 11648
rect 2225 11645 2237 11648
rect 2271 11645 2283 11679
rect 2225 11639 2283 11645
rect 768 11580 888 11608
rect 768 11404 796 11580
rect 1762 11568 1768 11620
rect 1820 11608 1826 11620
rect 2516 11608 2544 11716
rect 4433 11713 4445 11716
rect 4479 11713 4491 11747
rect 4433 11707 4491 11713
rect 4522 11704 4528 11756
rect 4580 11744 4586 11756
rect 4801 11747 4859 11753
rect 4801 11744 4813 11747
rect 4580 11716 4813 11744
rect 4580 11704 4586 11716
rect 4801 11713 4813 11716
rect 4847 11713 4859 11747
rect 4801 11707 4859 11713
rect 4982 11704 4988 11756
rect 5040 11744 5046 11756
rect 5077 11747 5135 11753
rect 5077 11744 5089 11747
rect 5040 11716 5089 11744
rect 5040 11704 5046 11716
rect 5077 11713 5089 11716
rect 5123 11713 5135 11747
rect 5077 11707 5135 11713
rect 5261 11747 5319 11753
rect 5261 11713 5273 11747
rect 5307 11744 5319 11747
rect 7190 11744 7196 11756
rect 5307 11716 7196 11744
rect 5307 11713 5319 11716
rect 5261 11707 5319 11713
rect 7190 11704 7196 11716
rect 7248 11704 7254 11756
rect 7558 11704 7564 11756
rect 7616 11744 7622 11756
rect 7926 11744 7932 11756
rect 7616 11716 7932 11744
rect 7616 11704 7622 11716
rect 7926 11704 7932 11716
rect 7984 11704 7990 11756
rect 8662 11704 8668 11756
rect 8720 11744 8726 11756
rect 8757 11747 8815 11753
rect 8757 11744 8769 11747
rect 8720 11716 8769 11744
rect 8720 11704 8726 11716
rect 8757 11713 8769 11716
rect 8803 11713 8815 11747
rect 9398 11744 9404 11756
rect 9359 11716 9404 11744
rect 8757 11707 8815 11713
rect 9398 11704 9404 11716
rect 9456 11704 9462 11756
rect 9766 11704 9772 11756
rect 9824 11744 9830 11756
rect 10134 11744 10140 11756
rect 9824 11716 10140 11744
rect 9824 11704 9830 11716
rect 10134 11704 10140 11716
rect 10192 11704 10198 11756
rect 12066 11753 12072 11756
rect 12060 11744 12072 11753
rect 12027 11716 12072 11744
rect 12060 11707 12072 11716
rect 12066 11704 12072 11707
rect 12124 11704 12130 11756
rect 12176 11744 12204 11784
rect 13262 11772 13268 11824
rect 13320 11812 13326 11824
rect 15488 11812 15516 11843
rect 15838 11840 15844 11892
rect 15896 11880 15902 11892
rect 23658 11880 23664 11892
rect 15896 11852 22094 11880
rect 23619 11852 23664 11880
rect 15896 11840 15902 11852
rect 16850 11812 16856 11824
rect 13320 11784 15516 11812
rect 16811 11784 16856 11812
rect 13320 11772 13326 11784
rect 16850 11772 16856 11784
rect 16908 11772 16914 11824
rect 17494 11772 17500 11824
rect 17552 11812 17558 11824
rect 18966 11812 18972 11824
rect 17552 11784 18972 11812
rect 17552 11772 17558 11784
rect 12618 11744 12624 11756
rect 12176 11716 12624 11744
rect 12618 11704 12624 11716
rect 12676 11704 12682 11756
rect 12802 11704 12808 11756
rect 12860 11744 12866 11756
rect 15289 11747 15347 11753
rect 15289 11744 15301 11747
rect 12860 11716 15301 11744
rect 12860 11704 12866 11716
rect 15289 11713 15301 11716
rect 15335 11713 15347 11747
rect 17034 11744 17040 11756
rect 16995 11716 17040 11744
rect 15289 11707 15347 11713
rect 17034 11704 17040 11716
rect 17092 11704 17098 11756
rect 17221 11747 17279 11753
rect 17221 11713 17233 11747
rect 17267 11744 17279 11747
rect 17678 11744 17684 11756
rect 17267 11716 17684 11744
rect 17267 11713 17279 11716
rect 17221 11707 17279 11713
rect 17678 11704 17684 11716
rect 17736 11704 17742 11756
rect 17862 11704 17868 11756
rect 17920 11744 17926 11756
rect 18708 11753 18736 11784
rect 18966 11772 18972 11784
rect 19024 11772 19030 11824
rect 20162 11812 20168 11824
rect 19352 11784 20168 11812
rect 19352 11753 19380 11784
rect 20162 11772 20168 11784
rect 20220 11772 20226 11824
rect 21358 11772 21364 11824
rect 21416 11812 21422 11824
rect 21913 11815 21971 11821
rect 21913 11812 21925 11815
rect 21416 11784 21925 11812
rect 21416 11772 21422 11784
rect 21913 11781 21925 11784
rect 21959 11781 21971 11815
rect 22066 11812 22094 11852
rect 23658 11840 23664 11852
rect 23716 11880 23722 11892
rect 24489 11883 24547 11889
rect 24489 11880 24501 11883
rect 23716 11852 24501 11880
rect 23716 11840 23722 11852
rect 24489 11849 24501 11852
rect 24535 11849 24547 11883
rect 24489 11843 24547 11849
rect 24762 11840 24768 11892
rect 24820 11880 24826 11892
rect 25241 11883 25299 11889
rect 25241 11880 25253 11883
rect 24820 11852 25253 11880
rect 24820 11840 24826 11852
rect 25241 11849 25253 11852
rect 25287 11849 25299 11883
rect 25241 11843 25299 11849
rect 27433 11883 27491 11889
rect 27433 11849 27445 11883
rect 27479 11880 27491 11883
rect 28166 11880 28172 11892
rect 27479 11852 28172 11880
rect 27479 11849 27491 11852
rect 27433 11843 27491 11849
rect 28166 11840 28172 11852
rect 28224 11840 28230 11892
rect 28902 11880 28908 11892
rect 28863 11852 28908 11880
rect 28902 11840 28908 11852
rect 28960 11840 28966 11892
rect 29546 11840 29552 11892
rect 29604 11840 29610 11892
rect 30282 11880 30288 11892
rect 30243 11852 30288 11880
rect 30282 11840 30288 11852
rect 30340 11840 30346 11892
rect 22066 11784 24532 11812
rect 21913 11775 21971 11781
rect 18417 11747 18475 11753
rect 18417 11744 18429 11747
rect 17920 11716 18429 11744
rect 17920 11704 17926 11716
rect 18417 11713 18429 11716
rect 18463 11713 18475 11747
rect 18417 11707 18475 11713
rect 18693 11747 18751 11753
rect 18693 11713 18705 11747
rect 18739 11713 18751 11747
rect 18693 11707 18751 11713
rect 18877 11747 18935 11753
rect 18877 11713 18889 11747
rect 18923 11744 18935 11747
rect 19337 11747 19395 11753
rect 18923 11716 19288 11744
rect 18923 11713 18935 11716
rect 18877 11707 18935 11713
rect 2682 11676 2688 11688
rect 2643 11648 2688 11676
rect 2682 11636 2688 11648
rect 2740 11636 2746 11688
rect 4614 11676 4620 11688
rect 4080 11648 4620 11676
rect 4080 11617 4108 11648
rect 4614 11636 4620 11648
rect 4672 11636 4678 11688
rect 6086 11636 6092 11688
rect 6144 11676 6150 11688
rect 6638 11676 6644 11688
rect 6144 11648 6644 11676
rect 6144 11636 6150 11648
rect 6638 11636 6644 11648
rect 6696 11636 6702 11688
rect 7009 11679 7067 11685
rect 7009 11645 7021 11679
rect 7055 11676 7067 11679
rect 7098 11676 7104 11688
rect 7055 11648 7104 11676
rect 7055 11645 7067 11648
rect 7009 11639 7067 11645
rect 7098 11636 7104 11648
rect 7156 11636 7162 11688
rect 7834 11636 7840 11688
rect 7892 11676 7898 11688
rect 8205 11679 8263 11685
rect 8205 11676 8217 11679
rect 7892 11648 8217 11676
rect 7892 11636 7898 11648
rect 8205 11645 8217 11648
rect 8251 11676 8263 11679
rect 9677 11679 9735 11685
rect 9677 11676 9689 11679
rect 8251 11648 9689 11676
rect 8251 11645 8263 11648
rect 8205 11639 8263 11645
rect 9677 11645 9689 11648
rect 9723 11676 9735 11679
rect 10318 11676 10324 11688
rect 9723 11648 10324 11676
rect 9723 11645 9735 11648
rect 9677 11639 9735 11645
rect 10318 11636 10324 11648
rect 10376 11636 10382 11688
rect 11790 11676 11796 11688
rect 11751 11648 11796 11676
rect 11790 11636 11796 11648
rect 11848 11636 11854 11688
rect 14093 11679 14151 11685
rect 14093 11645 14105 11679
rect 14139 11645 14151 11679
rect 14274 11676 14280 11688
rect 14235 11648 14280 11676
rect 14093 11639 14151 11645
rect 1820 11580 2544 11608
rect 4065 11611 4123 11617
rect 1820 11568 1826 11580
rect 4065 11577 4077 11611
rect 4111 11577 4123 11611
rect 4065 11571 4123 11577
rect 4433 11611 4491 11617
rect 4433 11577 4445 11611
rect 4479 11608 4491 11611
rect 4479 11580 9674 11608
rect 4479 11577 4491 11580
rect 4433 11571 4491 11577
rect 2133 11543 2191 11549
rect 2133 11509 2145 11543
rect 2179 11540 2191 11543
rect 3050 11540 3056 11552
rect 2179 11512 3056 11540
rect 2179 11509 2191 11512
rect 2133 11503 2191 11509
rect 3050 11500 3056 11512
rect 3108 11500 3114 11552
rect 4617 11543 4675 11549
rect 4617 11509 4629 11543
rect 4663 11540 4675 11543
rect 5258 11540 5264 11552
rect 4663 11512 5264 11540
rect 4663 11509 4675 11512
rect 4617 11503 4675 11509
rect 5258 11500 5264 11512
rect 5316 11500 5322 11552
rect 6178 11500 6184 11552
rect 6236 11540 6242 11552
rect 6365 11543 6423 11549
rect 6365 11540 6377 11543
rect 6236 11512 6377 11540
rect 6236 11500 6242 11512
rect 6365 11509 6377 11512
rect 6411 11509 6423 11543
rect 6365 11503 6423 11509
rect 7561 11543 7619 11549
rect 7561 11509 7573 11543
rect 7607 11540 7619 11543
rect 8294 11540 8300 11552
rect 7607 11512 8300 11540
rect 7607 11509 7619 11512
rect 7561 11503 7619 11509
rect 8294 11500 8300 11512
rect 8352 11500 8358 11552
rect 8849 11543 8907 11549
rect 8849 11509 8861 11543
rect 8895 11540 8907 11543
rect 9122 11540 9128 11552
rect 8895 11512 9128 11540
rect 8895 11509 8907 11512
rect 8849 11503 8907 11509
rect 9122 11500 9128 11512
rect 9180 11500 9186 11552
rect 9646 11540 9674 11580
rect 12894 11568 12900 11620
rect 12952 11608 12958 11620
rect 14108 11608 14136 11639
rect 14274 11636 14280 11648
rect 14332 11636 14338 11688
rect 16114 11636 16120 11688
rect 16172 11676 16178 11688
rect 17313 11679 17371 11685
rect 17313 11676 17325 11679
rect 16172 11648 17325 11676
rect 16172 11636 16178 11648
rect 17313 11645 17325 11648
rect 17359 11645 17371 11679
rect 18432 11676 18460 11707
rect 19150 11676 19156 11688
rect 18432 11648 19156 11676
rect 17313 11639 17371 11645
rect 19150 11636 19156 11648
rect 19208 11636 19214 11688
rect 18506 11608 18512 11620
rect 12952 11580 13768 11608
rect 14108 11580 18512 11608
rect 12952 11568 12958 11580
rect 12986 11540 12992 11552
rect 9646 11512 12992 11540
rect 12986 11500 12992 11512
rect 13044 11500 13050 11552
rect 13630 11540 13636 11552
rect 13591 11512 13636 11540
rect 13630 11500 13636 11512
rect 13688 11500 13694 11552
rect 13740 11540 13768 11580
rect 18506 11568 18512 11580
rect 18564 11568 18570 11620
rect 17310 11540 17316 11552
rect 13740 11512 17316 11540
rect 17310 11500 17316 11512
rect 17368 11500 17374 11552
rect 17494 11500 17500 11552
rect 17552 11540 17558 11552
rect 18233 11543 18291 11549
rect 18233 11540 18245 11543
rect 17552 11512 18245 11540
rect 17552 11500 17558 11512
rect 18233 11509 18245 11512
rect 18279 11509 18291 11543
rect 19260 11540 19288 11716
rect 19337 11713 19349 11747
rect 19383 11713 19395 11747
rect 19337 11707 19395 11713
rect 19604 11747 19662 11753
rect 19604 11713 19616 11747
rect 19650 11744 19662 11747
rect 20346 11744 20352 11756
rect 19650 11716 20352 11744
rect 19650 11713 19662 11716
rect 19604 11707 19662 11713
rect 20346 11704 20352 11716
rect 20404 11704 20410 11756
rect 21928 11744 21956 11775
rect 22741 11747 22799 11753
rect 22741 11744 22753 11747
rect 21928 11716 22753 11744
rect 22741 11713 22753 11716
rect 22787 11713 22799 11747
rect 23566 11744 23572 11756
rect 23527 11716 23572 11744
rect 22741 11707 22799 11713
rect 23566 11704 23572 11716
rect 23624 11704 23630 11756
rect 23793 11747 23851 11753
rect 23793 11744 23805 11747
rect 23768 11713 23805 11744
rect 23839 11713 23851 11747
rect 23934 11744 23940 11756
rect 23895 11716 23940 11744
rect 23768 11707 23851 11713
rect 20622 11636 20628 11688
rect 20680 11676 20686 11688
rect 23385 11679 23443 11685
rect 23385 11676 23397 11679
rect 20680 11648 23397 11676
rect 20680 11636 20686 11648
rect 23385 11645 23397 11648
rect 23431 11645 23443 11679
rect 23385 11639 23443 11645
rect 21634 11568 21640 11620
rect 21692 11608 21698 11620
rect 22094 11608 22100 11620
rect 21692 11580 22100 11608
rect 21692 11568 21698 11580
rect 22094 11568 22100 11580
rect 22152 11568 22158 11620
rect 22925 11611 22983 11617
rect 22925 11577 22937 11611
rect 22971 11608 22983 11611
rect 23014 11608 23020 11620
rect 22971 11580 23020 11608
rect 22971 11577 22983 11580
rect 22925 11571 22983 11577
rect 23014 11568 23020 11580
rect 23072 11568 23078 11620
rect 23198 11568 23204 11620
rect 23256 11608 23262 11620
rect 23768 11608 23796 11707
rect 23934 11704 23940 11716
rect 23992 11704 23998 11756
rect 24397 11747 24455 11753
rect 24397 11744 24409 11747
rect 24136 11716 24409 11744
rect 23256 11580 23796 11608
rect 23256 11568 23262 11580
rect 20438 11540 20444 11552
rect 19260 11512 20444 11540
rect 18233 11503 18291 11509
rect 20438 11500 20444 11512
rect 20496 11500 20502 11552
rect 20622 11500 20628 11552
rect 20680 11540 20686 11552
rect 20717 11543 20775 11549
rect 20717 11540 20729 11543
rect 20680 11512 20729 11540
rect 20680 11500 20686 11512
rect 20717 11509 20729 11512
rect 20763 11509 20775 11543
rect 20717 11503 20775 11509
rect 23290 11500 23296 11552
rect 23348 11540 23354 11552
rect 24136 11540 24164 11716
rect 24397 11713 24409 11716
rect 24443 11713 24455 11747
rect 24504 11744 24532 11784
rect 24578 11772 24584 11824
rect 24636 11812 24642 11824
rect 25041 11815 25099 11821
rect 25041 11812 25053 11815
rect 24636 11784 25053 11812
rect 24636 11772 24642 11784
rect 25041 11781 25053 11784
rect 25087 11781 25099 11815
rect 25041 11775 25099 11781
rect 25406 11772 25412 11824
rect 25464 11812 25470 11824
rect 27801 11815 27859 11821
rect 25464 11784 27752 11812
rect 25464 11772 25470 11784
rect 25961 11747 26019 11753
rect 25961 11744 25973 11747
rect 24504 11716 25973 11744
rect 24397 11707 24455 11713
rect 25961 11713 25973 11716
rect 26007 11713 26019 11747
rect 25961 11707 26019 11713
rect 27617 11747 27675 11753
rect 27617 11713 27629 11747
rect 27663 11713 27675 11747
rect 27724 11744 27752 11784
rect 27801 11781 27813 11815
rect 27847 11812 27859 11815
rect 27982 11812 27988 11824
rect 27847 11784 27988 11812
rect 27847 11781 27859 11784
rect 27801 11775 27859 11781
rect 27982 11772 27988 11784
rect 28040 11772 28046 11824
rect 29564 11812 29592 11840
rect 32320 11812 33120 11826
rect 29564 11784 31754 11812
rect 27893 11747 27951 11753
rect 27893 11744 27905 11747
rect 27724 11716 27905 11744
rect 27617 11707 27675 11713
rect 27893 11713 27905 11716
rect 27939 11713 27951 11747
rect 29086 11744 29092 11756
rect 29047 11716 29092 11744
rect 27893 11707 27951 11713
rect 27632 11676 27660 11707
rect 29086 11704 29092 11716
rect 29144 11704 29150 11756
rect 29362 11744 29368 11756
rect 29323 11716 29368 11744
rect 29362 11704 29368 11716
rect 29420 11704 29426 11756
rect 29549 11747 29607 11753
rect 29549 11713 29561 11747
rect 29595 11744 29607 11747
rect 29638 11744 29644 11756
rect 29595 11716 29644 11744
rect 29595 11713 29607 11716
rect 29549 11707 29607 11713
rect 29638 11704 29644 11716
rect 29696 11704 29702 11756
rect 29730 11704 29736 11756
rect 29788 11744 29794 11756
rect 30469 11747 30527 11753
rect 30469 11744 30481 11747
rect 29788 11716 30481 11744
rect 29788 11704 29794 11716
rect 30469 11713 30481 11716
rect 30515 11713 30527 11747
rect 30469 11707 30527 11713
rect 30745 11747 30803 11753
rect 30745 11713 30757 11747
rect 30791 11713 30803 11747
rect 30745 11707 30803 11713
rect 30929 11747 30987 11753
rect 30929 11713 30941 11747
rect 30975 11744 30987 11747
rect 31018 11744 31024 11756
rect 30975 11716 31024 11744
rect 30975 11713 30987 11716
rect 30929 11707 30987 11713
rect 28074 11676 28080 11688
rect 27632 11648 28080 11676
rect 28074 11636 28080 11648
rect 28132 11636 28138 11688
rect 29380 11676 29408 11704
rect 30760 11676 30788 11707
rect 31018 11704 31024 11716
rect 31076 11704 31082 11756
rect 29380 11648 30788 11676
rect 25409 11611 25467 11617
rect 25409 11577 25421 11611
rect 25455 11608 25467 11611
rect 31294 11608 31300 11620
rect 25455 11580 31300 11608
rect 25455 11577 25467 11580
rect 25409 11571 25467 11577
rect 31294 11568 31300 11580
rect 31352 11568 31358 11620
rect 25222 11540 25228 11552
rect 23348 11512 24164 11540
rect 25183 11512 25228 11540
rect 23348 11500 23354 11512
rect 25222 11500 25228 11512
rect 25280 11500 25286 11552
rect 26050 11540 26056 11552
rect 26011 11512 26056 11540
rect 26050 11500 26056 11512
rect 26108 11500 26114 11552
rect 29086 11500 29092 11552
rect 29144 11540 29150 11552
rect 29730 11540 29736 11552
rect 29144 11512 29736 11540
rect 29144 11500 29150 11512
rect 29730 11500 29736 11512
rect 29788 11500 29794 11552
rect 31726 11540 31754 11784
rect 32232 11784 33120 11812
rect 32232 11676 32260 11784
rect 32320 11770 33120 11784
rect 32232 11648 32352 11676
rect 32324 11540 32352 11648
rect 31726 11512 32352 11540
rect 1104 11450 32016 11472
rect 768 11376 888 11404
rect 1104 11398 2136 11450
rect 2188 11398 12440 11450
rect 12492 11398 22744 11450
rect 22796 11398 32016 11450
rect 1104 11376 32016 11398
rect 860 11336 888 11376
rect 2317 11339 2375 11345
rect 860 11308 1716 11336
rect 1688 11141 1716 11308
rect 2317 11305 2329 11339
rect 2363 11336 2375 11339
rect 2406 11336 2412 11348
rect 2363 11308 2412 11336
rect 2363 11305 2375 11308
rect 2317 11299 2375 11305
rect 2406 11296 2412 11308
rect 2464 11296 2470 11348
rect 3602 11336 3608 11348
rect 2516 11308 3608 11336
rect 1857 11271 1915 11277
rect 1857 11237 1869 11271
rect 1903 11268 1915 11271
rect 2516 11268 2544 11308
rect 3602 11296 3608 11308
rect 3660 11336 3666 11348
rect 4154 11336 4160 11348
rect 3660 11308 4160 11336
rect 3660 11296 3666 11308
rect 4154 11296 4160 11308
rect 4212 11296 4218 11348
rect 5074 11336 5080 11348
rect 5035 11308 5080 11336
rect 5074 11296 5080 11308
rect 5132 11296 5138 11348
rect 7469 11339 7527 11345
rect 7469 11305 7481 11339
rect 7515 11336 7527 11339
rect 12342 11336 12348 11348
rect 7515 11308 12348 11336
rect 7515 11305 7527 11308
rect 7469 11299 7527 11305
rect 12342 11296 12348 11308
rect 12400 11296 12406 11348
rect 12989 11339 13047 11345
rect 12989 11305 13001 11339
rect 13035 11336 13047 11339
rect 13722 11336 13728 11348
rect 13035 11308 13728 11336
rect 13035 11305 13047 11308
rect 12989 11299 13047 11305
rect 13722 11296 13728 11308
rect 13780 11296 13786 11348
rect 15194 11296 15200 11348
rect 15252 11336 15258 11348
rect 15378 11336 15384 11348
rect 15252 11308 15384 11336
rect 15252 11296 15258 11308
rect 15378 11296 15384 11308
rect 15436 11296 15442 11348
rect 17221 11339 17279 11345
rect 17221 11305 17233 11339
rect 17267 11305 17279 11339
rect 17221 11299 17279 11305
rect 5445 11271 5503 11277
rect 5445 11268 5457 11271
rect 1903 11240 2544 11268
rect 2608 11240 5457 11268
rect 1903 11237 1915 11240
rect 1857 11231 1915 11237
rect 2608 11200 2636 11240
rect 5445 11237 5457 11240
rect 5491 11237 5503 11271
rect 8757 11271 8815 11277
rect 8757 11268 8769 11271
rect 5445 11231 5503 11237
rect 7300 11240 8769 11268
rect 3142 11200 3148 11212
rect 1872 11172 2636 11200
rect 2700 11172 3148 11200
rect 1872 11144 1900 11172
rect 1673 11135 1731 11141
rect 1673 11101 1685 11135
rect 1719 11101 1731 11135
rect 1673 11095 1731 11101
rect 1854 11092 1860 11144
rect 1912 11092 1918 11144
rect 2501 11135 2559 11141
rect 2501 11101 2513 11135
rect 2547 11132 2559 11135
rect 2700 11132 2728 11172
rect 3142 11160 3148 11172
rect 3200 11200 3206 11212
rect 4065 11203 4123 11209
rect 4065 11200 4077 11203
rect 3200 11172 4077 11200
rect 3200 11160 3206 11172
rect 4065 11169 4077 11172
rect 4111 11169 4123 11203
rect 5534 11200 5540 11212
rect 5495 11172 5540 11200
rect 4065 11163 4123 11169
rect 5534 11160 5540 11172
rect 5592 11160 5598 11212
rect 6362 11160 6368 11212
rect 6420 11160 6426 11212
rect 2547 11104 2728 11132
rect 2547 11101 2559 11104
rect 2501 11095 2559 11101
rect 2774 11092 2780 11144
rect 2832 11132 2838 11144
rect 2958 11132 2964 11144
rect 2832 11104 2877 11132
rect 2919 11104 2964 11132
rect 2832 11092 2838 11104
rect 2958 11092 2964 11104
rect 3016 11092 3022 11144
rect 3789 11135 3847 11141
rect 3789 11101 3801 11135
rect 3835 11101 3847 11135
rect 3789 11095 3847 11101
rect 2866 11024 2872 11076
rect 2924 11064 2930 11076
rect 3804 11064 3832 11095
rect 4246 11092 4252 11144
rect 4304 11132 4310 11144
rect 4430 11132 4436 11144
rect 4304 11104 4436 11132
rect 4304 11092 4310 11104
rect 4430 11092 4436 11104
rect 4488 11092 4494 11144
rect 5258 11132 5264 11144
rect 5219 11104 5264 11132
rect 5258 11092 5264 11104
rect 5316 11092 5322 11144
rect 7300 11132 7328 11240
rect 8757 11237 8769 11240
rect 8803 11237 8815 11271
rect 8757 11231 8815 11237
rect 8941 11271 8999 11277
rect 8941 11237 8953 11271
rect 8987 11268 8999 11271
rect 9490 11268 9496 11280
rect 8987 11240 9496 11268
rect 8987 11237 8999 11240
rect 8941 11231 8999 11237
rect 9490 11228 9496 11240
rect 9548 11228 9554 11280
rect 12897 11271 12955 11277
rect 12897 11237 12909 11271
rect 12943 11268 12955 11271
rect 13630 11268 13636 11280
rect 12943 11240 13636 11268
rect 12943 11237 12955 11240
rect 12897 11231 12955 11237
rect 13630 11228 13636 11240
rect 13688 11228 13694 11280
rect 17236 11268 17264 11299
rect 17310 11296 17316 11348
rect 17368 11336 17374 11348
rect 19521 11339 19579 11345
rect 17368 11308 18552 11336
rect 17368 11296 17374 11308
rect 17678 11268 17684 11280
rect 17236 11240 17684 11268
rect 17678 11228 17684 11240
rect 17736 11228 17742 11280
rect 18239 11240 18359 11268
rect 7650 11160 7656 11212
rect 7708 11200 7714 11212
rect 9674 11200 9680 11212
rect 7708 11172 9260 11200
rect 9635 11172 9680 11200
rect 7708 11160 7714 11172
rect 5368 11104 7328 11132
rect 5368 11064 5396 11104
rect 7926 11092 7932 11144
rect 7984 11132 7990 11144
rect 8021 11135 8079 11141
rect 8021 11132 8033 11135
rect 7984 11104 8033 11132
rect 7984 11092 7990 11104
rect 8021 11101 8033 11104
rect 8067 11101 8079 11135
rect 8202 11132 8208 11144
rect 8163 11104 8208 11132
rect 8021 11095 8079 11101
rect 8202 11092 8208 11104
rect 8260 11092 8266 11144
rect 9030 11132 9036 11144
rect 8680 11104 9036 11132
rect 6178 11064 6184 11076
rect 2924 11036 5396 11064
rect 6139 11036 6184 11064
rect 2924 11024 2930 11036
rect 6178 11024 6184 11036
rect 6236 11024 6242 11076
rect 6454 11064 6460 11076
rect 6415 11036 6460 11064
rect 6454 11024 6460 11036
rect 6512 11024 6518 11076
rect 6546 11024 6552 11076
rect 6604 11064 6610 11076
rect 6604 11036 6649 11064
rect 6604 11024 6610 11036
rect 6730 11024 6736 11076
rect 6788 11064 6794 11076
rect 6917 11067 6975 11073
rect 6917 11064 6929 11067
rect 6788 11036 6929 11064
rect 6788 11024 6794 11036
rect 6917 11033 6929 11036
rect 6963 11033 6975 11067
rect 6917 11027 6975 11033
rect 7285 11067 7343 11073
rect 7285 11033 7297 11067
rect 7331 11064 7343 11067
rect 8389 11067 8447 11073
rect 8389 11064 8401 11067
rect 7331 11036 8401 11064
rect 7331 11033 7343 11036
rect 7285 11027 7343 11033
rect 8389 11033 8401 11036
rect 8435 11033 8447 11067
rect 8389 11027 8447 11033
rect 2222 10956 2228 11008
rect 2280 10996 2286 11008
rect 5994 10996 6000 11008
rect 2280 10968 6000 10996
rect 2280 10956 2286 10968
rect 5994 10956 6000 10968
rect 6052 10956 6058 11008
rect 7098 10956 7104 11008
rect 7156 10996 7162 11008
rect 7926 10996 7932 11008
rect 7156 10968 7932 10996
rect 7156 10956 7162 10968
rect 7926 10956 7932 10968
rect 7984 10956 7990 11008
rect 8018 10956 8024 11008
rect 8076 10996 8082 11008
rect 8680 10996 8708 11104
rect 9030 11092 9036 11104
rect 9088 11092 9094 11144
rect 9232 11141 9260 11172
rect 9674 11160 9680 11172
rect 9732 11160 9738 11212
rect 10410 11200 10416 11212
rect 10152 11172 10416 11200
rect 9217 11135 9275 11141
rect 9217 11101 9229 11135
rect 9263 11101 9275 11135
rect 9858 11132 9864 11144
rect 9819 11104 9864 11132
rect 9217 11095 9275 11101
rect 9858 11092 9864 11104
rect 9916 11092 9922 11144
rect 10152 11141 10180 11172
rect 10410 11160 10416 11172
rect 10468 11160 10474 11212
rect 12618 11200 12624 11212
rect 11440 11172 12624 11200
rect 10137 11135 10195 11141
rect 10137 11101 10149 11135
rect 10183 11101 10195 11135
rect 10318 11132 10324 11144
rect 10279 11104 10324 11132
rect 10137 11095 10195 11101
rect 10318 11092 10324 11104
rect 10376 11092 10382 11144
rect 11440 11141 11468 11172
rect 12618 11160 12624 11172
rect 12676 11160 12682 11212
rect 12728 11172 12940 11200
rect 11425 11135 11483 11141
rect 11425 11101 11437 11135
rect 11471 11101 11483 11135
rect 11425 11095 11483 11101
rect 11790 11092 11796 11144
rect 11848 11132 11854 11144
rect 12728 11132 12756 11172
rect 11848 11104 12756 11132
rect 12912 11132 12940 11172
rect 12986 11160 12992 11212
rect 13044 11200 13050 11212
rect 17494 11200 17500 11212
rect 13044 11172 14596 11200
rect 13044 11160 13050 11172
rect 14090 11132 14096 11144
rect 12912 11104 14096 11132
rect 11848 11092 11854 11104
rect 14090 11092 14096 11104
rect 14148 11132 14154 11144
rect 14461 11135 14519 11141
rect 14461 11132 14473 11135
rect 14148 11104 14473 11132
rect 14148 11092 14154 11104
rect 14461 11101 14473 11104
rect 14507 11101 14519 11135
rect 14568 11132 14596 11172
rect 17052 11172 17500 11200
rect 17052 11141 17080 11172
rect 17494 11160 17500 11172
rect 17552 11160 17558 11212
rect 18239 11200 18267 11240
rect 18331 11212 18359 11240
rect 17880 11172 18267 11200
rect 14717 11135 14775 11141
rect 14717 11132 14729 11135
rect 14568 11104 14729 11132
rect 14461 11095 14519 11101
rect 14717 11101 14729 11104
rect 14763 11101 14775 11135
rect 14717 11095 14775 11101
rect 17037 11135 17095 11141
rect 17037 11101 17049 11135
rect 17083 11101 17095 11135
rect 17037 11095 17095 11101
rect 17313 11135 17371 11141
rect 17313 11101 17325 11135
rect 17359 11132 17371 11135
rect 17880 11132 17908 11172
rect 18322 11160 18328 11212
rect 18380 11200 18386 11212
rect 18380 11172 18473 11200
rect 18380 11160 18386 11172
rect 17359 11104 17908 11132
rect 18049 11135 18107 11141
rect 18049 11129 18061 11135
rect 17359 11101 17371 11104
rect 17313 11095 17371 11101
rect 17972 11101 18061 11129
rect 18095 11101 18107 11135
rect 8938 11064 8944 11076
rect 8899 11036 8944 11064
rect 8938 11024 8944 11036
rect 8996 11024 9002 11076
rect 9122 11064 9128 11076
rect 9083 11036 9128 11064
rect 9122 11024 9128 11036
rect 9180 11024 9186 11076
rect 11609 11067 11667 11073
rect 11609 11064 11621 11067
rect 9223 11036 11621 11064
rect 8076 10968 8708 10996
rect 8757 10999 8815 11005
rect 8076 10956 8082 10968
rect 8757 10965 8769 10999
rect 8803 10996 8815 10999
rect 9223 10996 9251 11036
rect 11609 11033 11621 11036
rect 11655 11033 11667 11067
rect 11609 11027 11667 11033
rect 12529 11067 12587 11073
rect 12529 11033 12541 11067
rect 12575 11064 12587 11067
rect 12710 11064 12716 11076
rect 12575 11036 12716 11064
rect 12575 11033 12587 11036
rect 12529 11027 12587 11033
rect 12710 11024 12716 11036
rect 12768 11024 12774 11076
rect 17972 11008 18000 11101
rect 18049 11095 18107 11101
rect 18141 11135 18199 11141
rect 18141 11101 18153 11135
rect 18187 11101 18199 11135
rect 18141 11095 18199 11101
rect 18156 11064 18184 11095
rect 18230 11092 18236 11144
rect 18288 11132 18294 11144
rect 18432 11141 18460 11172
rect 18417 11135 18475 11141
rect 18288 11104 18333 11132
rect 18288 11092 18294 11104
rect 18417 11101 18429 11135
rect 18463 11101 18475 11135
rect 18524 11132 18552 11308
rect 19521 11305 19533 11339
rect 19567 11336 19579 11339
rect 21174 11336 21180 11348
rect 19567 11308 21180 11336
rect 19567 11305 19579 11308
rect 19521 11299 19579 11305
rect 21174 11296 21180 11308
rect 21232 11296 21238 11348
rect 24949 11339 25007 11345
rect 24949 11305 24961 11339
rect 24995 11336 25007 11339
rect 28905 11339 28963 11345
rect 24995 11308 28856 11336
rect 24995 11305 25007 11308
rect 24949 11299 25007 11305
rect 22186 11228 22192 11280
rect 22244 11268 22250 11280
rect 23474 11268 23480 11280
rect 22244 11240 23480 11268
rect 22244 11228 22250 11240
rect 23474 11228 23480 11240
rect 23532 11228 23538 11280
rect 28074 11268 28080 11280
rect 28035 11240 28080 11268
rect 28074 11228 28080 11240
rect 28132 11228 28138 11280
rect 28828 11268 28856 11308
rect 28905 11305 28917 11339
rect 28951 11336 28963 11339
rect 29914 11336 29920 11348
rect 28951 11308 29920 11336
rect 28951 11305 28963 11308
rect 28905 11299 28963 11305
rect 29914 11296 29920 11308
rect 29972 11336 29978 11348
rect 31021 11339 31079 11345
rect 31021 11336 31033 11339
rect 29972 11308 31033 11336
rect 29972 11296 29978 11308
rect 31021 11305 31033 11308
rect 31067 11305 31079 11339
rect 31021 11299 31079 11305
rect 29089 11271 29147 11277
rect 29089 11268 29101 11271
rect 28828 11240 29101 11268
rect 29089 11237 29101 11240
rect 29135 11237 29147 11271
rect 29089 11231 29147 11237
rect 29178 11228 29184 11280
rect 29236 11268 29242 11280
rect 29236 11240 30144 11268
rect 29236 11228 29242 11240
rect 20165 11203 20223 11209
rect 20165 11169 20177 11203
rect 20211 11200 20223 11203
rect 20438 11200 20444 11212
rect 20211 11172 20444 11200
rect 20211 11169 20223 11172
rect 20165 11163 20223 11169
rect 20438 11160 20444 11172
rect 20496 11160 20502 11212
rect 20806 11200 20812 11212
rect 20767 11172 20812 11200
rect 20806 11160 20812 11172
rect 20864 11160 20870 11212
rect 21910 11160 21916 11212
rect 21968 11200 21974 11212
rect 29549 11203 29607 11209
rect 29549 11200 29561 11203
rect 21968 11172 24900 11200
rect 21968 11160 21974 11172
rect 19889 11135 19947 11141
rect 19889 11132 19901 11135
rect 18524 11104 19901 11132
rect 18417 11095 18475 11101
rect 19889 11101 19901 11104
rect 19935 11101 19947 11135
rect 19889 11095 19947 11101
rect 19981 11135 20039 11141
rect 19981 11101 19993 11135
rect 20027 11132 20039 11135
rect 20898 11132 20904 11144
rect 20027 11104 20904 11132
rect 20027 11101 20039 11104
rect 19981 11095 20039 11101
rect 20898 11092 20904 11104
rect 20956 11092 20962 11144
rect 22554 11092 22560 11144
rect 22612 11132 22618 11144
rect 22833 11135 22891 11141
rect 22833 11132 22845 11135
rect 22612 11104 22845 11132
rect 22612 11092 22618 11104
rect 22833 11101 22845 11104
rect 22879 11101 22891 11135
rect 22833 11095 22891 11101
rect 23109 11135 23167 11141
rect 23109 11101 23121 11135
rect 23155 11101 23167 11135
rect 23109 11095 23167 11101
rect 18064 11036 18184 11064
rect 18064 11008 18092 11036
rect 18506 11024 18512 11076
rect 18564 11064 18570 11076
rect 21076 11067 21134 11073
rect 18564 11036 21036 11064
rect 18564 11024 18570 11036
rect 8803 10968 9251 10996
rect 8803 10965 8815 10968
rect 8757 10959 8815 10965
rect 15194 10956 15200 11008
rect 15252 10996 15258 11008
rect 15841 10999 15899 11005
rect 15841 10996 15853 10999
rect 15252 10968 15853 10996
rect 15252 10956 15258 10968
rect 15841 10965 15853 10968
rect 15887 10965 15899 10999
rect 15841 10959 15899 10965
rect 16853 10999 16911 11005
rect 16853 10965 16865 10999
rect 16899 10996 16911 10999
rect 17494 10996 17500 11008
rect 16899 10968 17500 10996
rect 16899 10965 16911 10968
rect 16853 10959 16911 10965
rect 17494 10956 17500 10968
rect 17552 10956 17558 11008
rect 17773 10999 17831 11005
rect 17773 10965 17785 10999
rect 17819 10996 17831 10999
rect 17862 10996 17868 11008
rect 17819 10968 17868 10996
rect 17819 10965 17831 10968
rect 17773 10959 17831 10965
rect 17862 10956 17868 10968
rect 17920 10956 17926 11008
rect 17954 10956 17960 11008
rect 18012 10956 18018 11008
rect 18046 10956 18052 11008
rect 18104 10996 18110 11008
rect 19610 10996 19616 11008
rect 18104 10968 19616 10996
rect 18104 10956 18110 10968
rect 19610 10956 19616 10968
rect 19668 10956 19674 11008
rect 21008 10996 21036 11036
rect 21076 11033 21088 11067
rect 21122 11064 21134 11067
rect 21726 11064 21732 11076
rect 21122 11036 21732 11064
rect 21122 11033 21134 11036
rect 21076 11027 21134 11033
rect 21726 11024 21732 11036
rect 21784 11024 21790 11076
rect 22278 11024 22284 11076
rect 22336 11064 22342 11076
rect 22649 11067 22707 11073
rect 22336 11036 22600 11064
rect 22336 11024 22342 11036
rect 22189 10999 22247 11005
rect 22189 10996 22201 10999
rect 21008 10968 22201 10996
rect 22189 10965 22201 10968
rect 22235 10996 22247 10999
rect 22462 10996 22468 11008
rect 22235 10968 22468 10996
rect 22235 10965 22247 10968
rect 22189 10959 22247 10965
rect 22462 10956 22468 10968
rect 22520 10956 22526 11008
rect 22572 10996 22600 11036
rect 22649 11033 22661 11067
rect 22695 11064 22707 11067
rect 22922 11064 22928 11076
rect 22695 11036 22928 11064
rect 22695 11033 22707 11036
rect 22649 11027 22707 11033
rect 22922 11024 22928 11036
rect 22980 11024 22986 11076
rect 23124 11064 23152 11095
rect 23198 11092 23204 11144
rect 23256 11132 23262 11144
rect 24872 11141 24900 11172
rect 28736 11172 29561 11200
rect 23293 11135 23351 11141
rect 23293 11132 23305 11135
rect 23256 11104 23305 11132
rect 23256 11092 23262 11104
rect 23293 11101 23305 11104
rect 23339 11101 23351 11135
rect 23293 11095 23351 11101
rect 24857 11135 24915 11141
rect 24857 11101 24869 11135
rect 24903 11101 24915 11135
rect 25682 11132 25688 11144
rect 25643 11104 25688 11132
rect 24857 11095 24915 11101
rect 25682 11092 25688 11104
rect 25740 11092 25746 11144
rect 25866 11132 25872 11144
rect 25827 11104 25872 11132
rect 25866 11092 25872 11104
rect 25924 11092 25930 11144
rect 25961 11135 26019 11141
rect 25961 11101 25973 11135
rect 26007 11101 26019 11135
rect 26694 11132 26700 11144
rect 26655 11104 26700 11132
rect 25961 11095 26019 11101
rect 23382 11064 23388 11076
rect 23124 11036 23388 11064
rect 23124 10996 23152 11036
rect 23382 11024 23388 11036
rect 23440 11064 23446 11076
rect 25498 11064 25504 11076
rect 23440 11036 24532 11064
rect 25459 11036 25504 11064
rect 23440 11024 23446 11036
rect 22572 10968 23152 10996
rect 23198 10956 23204 11008
rect 23256 10996 23262 11008
rect 24394 10996 24400 11008
rect 23256 10968 24400 10996
rect 23256 10956 23262 10968
rect 24394 10956 24400 10968
rect 24452 10956 24458 11008
rect 24504 10996 24532 11036
rect 25498 11024 25504 11036
rect 25556 11024 25562 11076
rect 25976 11064 26004 11095
rect 26694 11092 26700 11104
rect 26752 11092 26758 11144
rect 26786 11092 26792 11144
rect 26844 11132 26850 11144
rect 28736 11141 28764 11172
rect 29549 11169 29561 11172
rect 29595 11169 29607 11203
rect 29549 11163 29607 11169
rect 30116 11200 30144 11240
rect 31113 11203 31171 11209
rect 31113 11200 31125 11203
rect 30116 11172 31125 11200
rect 26953 11135 27011 11141
rect 26953 11132 26965 11135
rect 26844 11104 26965 11132
rect 26844 11092 26850 11104
rect 26953 11101 26965 11104
rect 26999 11101 27011 11135
rect 26953 11095 27011 11101
rect 28721 11135 28779 11141
rect 28721 11101 28733 11135
rect 28767 11101 28779 11135
rect 28721 11095 28779 11101
rect 28997 11135 29055 11141
rect 28997 11101 29009 11135
rect 29043 11132 29055 11135
rect 29638 11132 29644 11144
rect 29043 11104 29644 11132
rect 29043 11101 29055 11104
rect 28997 11095 29055 11101
rect 29638 11092 29644 11104
rect 29696 11092 29702 11144
rect 29730 11092 29736 11144
rect 29788 11132 29794 11144
rect 30009 11135 30067 11141
rect 29788 11104 29833 11132
rect 29788 11092 29794 11104
rect 30009 11101 30021 11135
rect 30055 11101 30067 11135
rect 30116 11132 30144 11172
rect 31113 11169 31125 11172
rect 31159 11169 31171 11203
rect 31113 11163 31171 11169
rect 30190 11132 30196 11144
rect 30116 11104 30196 11132
rect 30009 11095 30067 11101
rect 27246 11064 27252 11076
rect 25976 11036 27252 11064
rect 27246 11024 27252 11036
rect 27304 11024 27310 11076
rect 28537 11067 28595 11073
rect 28537 11033 28549 11067
rect 28583 11064 28595 11067
rect 29089 11067 29147 11073
rect 28583 11036 29040 11064
rect 28583 11033 28595 11036
rect 28537 11027 28595 11033
rect 29012 11008 29040 11036
rect 29089 11033 29101 11067
rect 29135 11064 29147 11067
rect 29270 11064 29276 11076
rect 29135 11036 29276 11064
rect 29135 11033 29147 11036
rect 29089 11027 29147 11033
rect 29270 11024 29276 11036
rect 29328 11024 29334 11076
rect 29362 11024 29368 11076
rect 29420 11064 29426 11076
rect 30024 11064 30052 11095
rect 30190 11092 30196 11104
rect 30248 11132 30254 11144
rect 30834 11132 30840 11144
rect 30248 11104 30341 11132
rect 30795 11104 30840 11132
rect 30248 11092 30254 11104
rect 30834 11092 30840 11104
rect 30892 11092 30898 11144
rect 29420 11036 30052 11064
rect 29420 11024 29426 11036
rect 29656 11008 29684 11036
rect 30098 11024 30104 11076
rect 30156 11064 30162 11076
rect 30653 11067 30711 11073
rect 30653 11064 30665 11067
rect 30156 11036 30665 11064
rect 30156 11024 30162 11036
rect 30653 11033 30665 11036
rect 30699 11033 30711 11067
rect 30653 11027 30711 11033
rect 25958 10996 25964 11008
rect 24504 10968 25964 10996
rect 25958 10956 25964 10968
rect 26016 10956 26022 11008
rect 28994 10956 29000 11008
rect 29052 10956 29058 11008
rect 29638 10956 29644 11008
rect 29696 10956 29702 11008
rect 1104 10906 32016 10928
rect 1104 10854 7288 10906
rect 7340 10854 17592 10906
rect 17644 10854 27896 10906
rect 27948 10854 32016 10906
rect 1104 10832 32016 10854
rect 2866 10752 2872 10804
rect 2924 10752 2930 10804
rect 5629 10795 5687 10801
rect 5629 10761 5641 10795
rect 5675 10761 5687 10795
rect 6730 10792 6736 10804
rect 6691 10764 6736 10792
rect 5629 10755 5687 10761
rect 1854 10684 1860 10736
rect 1912 10724 1918 10736
rect 2884 10724 2912 10752
rect 1912 10696 2912 10724
rect 1912 10684 1918 10696
rect 4522 10684 4528 10736
rect 4580 10724 4586 10736
rect 5644 10724 5672 10755
rect 6730 10752 6736 10764
rect 6788 10752 6794 10804
rect 8113 10795 8171 10801
rect 8113 10761 8125 10795
rect 8159 10792 8171 10795
rect 8159 10764 8294 10792
rect 8159 10761 8171 10764
rect 8113 10755 8171 10761
rect 7745 10727 7803 10733
rect 7745 10724 7757 10727
rect 4580 10696 4752 10724
rect 5644 10696 7757 10724
rect 4580 10684 4586 10696
rect 1949 10659 2007 10665
rect 1949 10625 1961 10659
rect 1995 10656 2007 10659
rect 2038 10656 2044 10668
rect 1995 10628 2044 10656
rect 1995 10625 2007 10628
rect 1949 10619 2007 10625
rect 2038 10616 2044 10628
rect 2096 10616 2102 10668
rect 2222 10656 2228 10668
rect 2183 10628 2228 10656
rect 2222 10616 2228 10628
rect 2280 10616 2286 10668
rect 2314 10616 2320 10668
rect 2372 10656 2378 10668
rect 4724 10665 4752 10696
rect 7745 10693 7757 10696
rect 7791 10693 7803 10727
rect 7917 10724 7923 10736
rect 7878 10696 7923 10724
rect 7745 10687 7803 10693
rect 7917 10684 7923 10696
rect 7975 10684 7981 10736
rect 8266 10724 8294 10764
rect 8570 10752 8576 10804
rect 8628 10792 8634 10804
rect 14185 10795 14243 10801
rect 14185 10792 14197 10795
rect 8628 10764 14197 10792
rect 8628 10752 8634 10764
rect 14185 10761 14197 10764
rect 14231 10761 14243 10795
rect 14185 10755 14243 10761
rect 15010 10752 15016 10804
rect 15068 10792 15074 10804
rect 15068 10764 16968 10792
rect 15068 10752 15074 10764
rect 8481 10727 8539 10733
rect 8266 10696 8340 10724
rect 3329 10659 3387 10665
rect 3329 10656 3341 10659
rect 2372 10628 3341 10656
rect 2372 10616 2378 10628
rect 3329 10625 3341 10628
rect 3375 10625 3387 10659
rect 3329 10619 3387 10625
rect 4709 10659 4767 10665
rect 4709 10625 4721 10659
rect 4755 10625 4767 10659
rect 4982 10656 4988 10668
rect 4943 10628 4988 10656
rect 4709 10619 4767 10625
rect 1486 10548 1492 10600
rect 1544 10588 1550 10600
rect 1762 10588 1768 10600
rect 1544 10560 1768 10588
rect 1544 10548 1550 10560
rect 1762 10548 1768 10560
rect 1820 10588 1826 10600
rect 2133 10591 2191 10597
rect 2133 10588 2145 10591
rect 1820 10560 2145 10588
rect 1820 10548 1826 10560
rect 2133 10557 2145 10560
rect 2179 10557 2191 10591
rect 2133 10551 2191 10557
rect 3050 10548 3056 10600
rect 3108 10588 3114 10600
rect 3145 10591 3203 10597
rect 3145 10588 3157 10591
rect 3108 10560 3157 10588
rect 3108 10548 3114 10560
rect 3145 10557 3157 10560
rect 3191 10557 3203 10591
rect 3145 10551 3203 10557
rect 3237 10591 3295 10597
rect 3237 10557 3249 10591
rect 3283 10557 3295 10591
rect 3237 10551 3295 10557
rect 3421 10591 3479 10597
rect 3421 10557 3433 10591
rect 3467 10588 3479 10591
rect 4522 10588 4528 10600
rect 3467 10560 4528 10588
rect 3467 10557 3479 10560
rect 3421 10551 3479 10557
rect 2774 10480 2780 10532
rect 2832 10520 2838 10532
rect 3252 10520 3280 10551
rect 4522 10548 4528 10560
rect 4580 10548 4586 10600
rect 4724 10588 4752 10619
rect 4982 10616 4988 10628
rect 5040 10616 5046 10668
rect 5169 10659 5227 10665
rect 5169 10625 5181 10659
rect 5215 10656 5227 10659
rect 5626 10656 5632 10668
rect 5215 10628 5632 10656
rect 5215 10625 5227 10628
rect 5169 10619 5227 10625
rect 5626 10616 5632 10628
rect 5684 10616 5690 10668
rect 5813 10659 5871 10665
rect 5813 10625 5825 10659
rect 5859 10656 5871 10659
rect 5994 10656 6000 10668
rect 5859 10628 6000 10656
rect 5859 10625 5871 10628
rect 5813 10619 5871 10625
rect 5994 10616 6000 10628
rect 6052 10616 6058 10668
rect 7006 10616 7012 10668
rect 7064 10656 7070 10668
rect 7101 10659 7159 10665
rect 7101 10656 7113 10659
rect 7064 10628 7113 10656
rect 7064 10616 7070 10628
rect 7101 10625 7113 10628
rect 7147 10656 7159 10659
rect 7650 10656 7656 10668
rect 7147 10628 7656 10656
rect 7147 10625 7159 10628
rect 7101 10619 7159 10625
rect 7650 10616 7656 10628
rect 7708 10616 7714 10668
rect 8110 10616 8116 10668
rect 8168 10656 8174 10668
rect 8205 10659 8263 10665
rect 8205 10656 8217 10659
rect 8168 10628 8217 10656
rect 8168 10616 8174 10628
rect 8205 10625 8217 10628
rect 8251 10625 8263 10659
rect 8312 10656 8340 10696
rect 8481 10693 8493 10727
rect 8527 10724 8539 10727
rect 10134 10724 10140 10736
rect 8527 10696 10140 10724
rect 8527 10693 8539 10696
rect 8481 10687 8539 10693
rect 10134 10684 10140 10696
rect 10192 10684 10198 10736
rect 10229 10727 10287 10733
rect 10229 10693 10241 10727
rect 10275 10724 10287 10727
rect 10275 10696 11744 10724
rect 10275 10693 10287 10696
rect 10229 10687 10287 10693
rect 8570 10656 8576 10668
rect 8312 10628 8576 10656
rect 8205 10619 8263 10625
rect 8570 10616 8576 10628
rect 8628 10616 8634 10668
rect 8665 10659 8723 10665
rect 8665 10625 8677 10659
rect 8711 10625 8723 10659
rect 8665 10619 8723 10625
rect 9309 10659 9367 10665
rect 9309 10625 9321 10659
rect 9355 10625 9367 10659
rect 9490 10656 9496 10668
rect 9451 10628 9496 10656
rect 9309 10619 9367 10625
rect 4798 10588 4804 10600
rect 4724 10560 4804 10588
rect 4798 10548 4804 10560
rect 4856 10548 4862 10600
rect 7190 10588 7196 10600
rect 4908 10560 7196 10588
rect 2832 10492 3280 10520
rect 2832 10480 2838 10492
rect 3602 10480 3608 10532
rect 3660 10520 3666 10532
rect 4908 10520 4936 10560
rect 7190 10548 7196 10560
rect 7248 10548 7254 10600
rect 7285 10591 7343 10597
rect 7285 10557 7297 10591
rect 7331 10557 7343 10591
rect 7285 10551 7343 10557
rect 7837 10591 7895 10597
rect 7837 10557 7849 10591
rect 7883 10588 7895 10591
rect 8481 10591 8539 10597
rect 8481 10588 8493 10591
rect 7883 10560 8493 10588
rect 7883 10557 7895 10560
rect 7837 10551 7895 10557
rect 8481 10557 8493 10560
rect 8527 10557 8539 10591
rect 8481 10551 8539 10557
rect 3660 10492 4936 10520
rect 3660 10480 3666 10492
rect 6914 10480 6920 10532
rect 6972 10520 6978 10532
rect 7300 10520 7328 10551
rect 8680 10520 8708 10619
rect 9324 10588 9352 10619
rect 9490 10616 9496 10628
rect 9548 10616 9554 10668
rect 9858 10616 9864 10668
rect 9916 10656 9922 10668
rect 11716 10665 11744 10696
rect 12618 10684 12624 10736
rect 12676 10724 12682 10736
rect 13265 10727 13323 10733
rect 13265 10724 13277 10727
rect 12676 10696 13277 10724
rect 12676 10684 12682 10696
rect 13265 10693 13277 10696
rect 13311 10693 13323 10727
rect 13265 10687 13323 10693
rect 13354 10684 13360 10736
rect 13412 10724 13418 10736
rect 13725 10727 13783 10733
rect 13725 10724 13737 10727
rect 13412 10696 13737 10724
rect 13412 10684 13418 10696
rect 13725 10693 13737 10696
rect 13771 10724 13783 10727
rect 15841 10727 15899 10733
rect 15841 10724 15853 10727
rect 13771 10696 15853 10724
rect 13771 10693 13783 10696
rect 13725 10687 13783 10693
rect 15841 10693 15853 10696
rect 15887 10724 15899 10727
rect 15930 10724 15936 10736
rect 15887 10696 15936 10724
rect 15887 10693 15899 10696
rect 15841 10687 15899 10693
rect 15930 10684 15936 10696
rect 15988 10684 15994 10736
rect 10413 10659 10471 10665
rect 10413 10656 10425 10659
rect 9916 10628 10425 10656
rect 9916 10616 9922 10628
rect 10244 10600 10272 10628
rect 10413 10625 10425 10628
rect 10459 10625 10471 10659
rect 10413 10619 10471 10625
rect 10689 10659 10747 10665
rect 10689 10625 10701 10659
rect 10735 10625 10747 10659
rect 10689 10619 10747 10625
rect 10873 10659 10931 10665
rect 10873 10625 10885 10659
rect 10919 10656 10931 10659
rect 10965 10659 11023 10665
rect 10965 10656 10977 10659
rect 10919 10628 10977 10656
rect 10919 10625 10931 10628
rect 10873 10619 10931 10625
rect 10965 10625 10977 10628
rect 11011 10625 11023 10659
rect 10965 10619 11023 10625
rect 11701 10659 11759 10665
rect 11701 10625 11713 10659
rect 11747 10625 11759 10659
rect 11701 10619 11759 10625
rect 9674 10588 9680 10600
rect 9324 10560 9680 10588
rect 9674 10548 9680 10560
rect 9732 10548 9738 10600
rect 10226 10548 10232 10600
rect 10284 10548 10290 10600
rect 10704 10588 10732 10619
rect 12986 10616 12992 10668
rect 13044 10656 13050 10668
rect 13081 10659 13139 10665
rect 13081 10656 13093 10659
rect 13044 10628 13093 10656
rect 13044 10616 13050 10628
rect 13081 10625 13093 10628
rect 13127 10625 13139 10659
rect 13081 10619 13139 10625
rect 14642 10616 14648 10668
rect 14700 10656 14706 10668
rect 15013 10659 15071 10665
rect 15013 10656 15025 10659
rect 14700 10628 15025 10656
rect 14700 10616 14706 10628
rect 15013 10625 15025 10628
rect 15059 10625 15071 10659
rect 15194 10656 15200 10668
rect 15155 10628 15200 10656
rect 15013 10619 15071 10625
rect 11054 10588 11060 10600
rect 10704 10560 11060 10588
rect 11054 10548 11060 10560
rect 11112 10588 11118 10600
rect 11882 10588 11888 10600
rect 11112 10560 11888 10588
rect 11112 10548 11118 10560
rect 11882 10548 11888 10560
rect 11940 10548 11946 10600
rect 11977 10591 12035 10597
rect 11977 10557 11989 10591
rect 12023 10557 12035 10591
rect 15028 10588 15056 10619
rect 15194 10616 15200 10628
rect 15252 10616 15258 10668
rect 16022 10656 16028 10668
rect 15983 10628 16028 10656
rect 16022 10616 16028 10628
rect 16080 10616 16086 10668
rect 16114 10616 16120 10668
rect 16172 10656 16178 10668
rect 16853 10659 16911 10665
rect 16172 10628 16217 10656
rect 16172 10616 16178 10628
rect 16853 10625 16865 10659
rect 16899 10625 16911 10659
rect 16940 10656 16968 10764
rect 17862 10752 17868 10804
rect 17920 10792 17926 10804
rect 18414 10792 18420 10804
rect 17920 10764 18420 10792
rect 17920 10752 17926 10764
rect 18414 10752 18420 10764
rect 18472 10752 18478 10804
rect 20257 10795 20315 10801
rect 20257 10761 20269 10795
rect 20303 10792 20315 10795
rect 20533 10795 20591 10801
rect 20533 10792 20545 10795
rect 20303 10764 20545 10792
rect 20303 10761 20315 10764
rect 20257 10755 20315 10761
rect 20533 10761 20545 10764
rect 20579 10761 20591 10795
rect 20533 10755 20591 10761
rect 20898 10752 20904 10804
rect 20956 10792 20962 10804
rect 20956 10764 21772 10792
rect 20956 10752 20962 10764
rect 17954 10724 17960 10736
rect 17144 10696 17960 10724
rect 17144 10665 17172 10696
rect 17954 10684 17960 10696
rect 18012 10684 18018 10736
rect 19058 10684 19064 10736
rect 19116 10724 19122 10736
rect 19426 10724 19432 10736
rect 19116 10696 19432 10724
rect 19116 10684 19122 10696
rect 19426 10684 19432 10696
rect 19484 10724 19490 10736
rect 20073 10727 20131 10733
rect 20073 10724 20085 10727
rect 19484 10696 20085 10724
rect 19484 10684 19490 10696
rect 20073 10693 20085 10696
rect 20119 10693 20131 10727
rect 20622 10724 20628 10736
rect 20073 10687 20131 10693
rect 20180 10696 20628 10724
rect 17037 10659 17095 10665
rect 17037 10656 17049 10659
rect 16940 10628 17049 10656
rect 16853 10619 16911 10625
rect 17037 10625 17049 10628
rect 17083 10625 17095 10659
rect 17037 10619 17095 10625
rect 17129 10659 17187 10665
rect 17129 10625 17141 10659
rect 17175 10625 17187 10659
rect 17129 10619 17187 10625
rect 16666 10588 16672 10600
rect 15028 10560 15516 10588
rect 16627 10560 16672 10588
rect 11977 10551 12035 10557
rect 6972 10492 7328 10520
rect 8036 10492 8708 10520
rect 8941 10523 8999 10529
rect 6972 10480 6978 10492
rect 1762 10452 1768 10464
rect 1723 10424 1768 10452
rect 1762 10412 1768 10424
rect 1820 10412 1826 10464
rect 2961 10455 3019 10461
rect 2961 10421 2973 10455
rect 3007 10452 3019 10455
rect 4430 10452 4436 10464
rect 3007 10424 4436 10452
rect 3007 10421 3019 10424
rect 2961 10415 3019 10421
rect 4430 10412 4436 10424
rect 4488 10412 4494 10464
rect 4525 10455 4583 10461
rect 4525 10421 4537 10455
rect 4571 10452 4583 10455
rect 5074 10452 5080 10464
rect 4571 10424 5080 10452
rect 4571 10421 4583 10424
rect 4525 10415 4583 10421
rect 5074 10412 5080 10424
rect 5132 10412 5138 10464
rect 5718 10412 5724 10464
rect 5776 10452 5782 10464
rect 7742 10452 7748 10464
rect 5776 10424 7748 10452
rect 5776 10412 5782 10424
rect 7742 10412 7748 10424
rect 7800 10412 7806 10464
rect 7929 10455 7987 10461
rect 7929 10421 7941 10455
rect 7975 10452 7987 10455
rect 8036 10452 8064 10492
rect 8941 10489 8953 10523
rect 8987 10520 8999 10523
rect 9582 10520 9588 10532
rect 8987 10492 9588 10520
rect 8987 10489 8999 10492
rect 8941 10483 8999 10489
rect 9582 10480 9588 10492
rect 9640 10480 9646 10532
rect 10318 10480 10324 10532
rect 10376 10520 10382 10532
rect 11992 10520 12020 10551
rect 10376 10492 12020 10520
rect 14093 10523 14151 10529
rect 10376 10480 10382 10492
rect 14093 10489 14105 10523
rect 14139 10520 14151 10523
rect 14274 10520 14280 10532
rect 14139 10492 14280 10520
rect 14139 10489 14151 10492
rect 14093 10483 14151 10489
rect 14274 10480 14280 10492
rect 14332 10520 14338 10532
rect 15381 10523 15439 10529
rect 15381 10520 15393 10523
rect 14332 10492 15393 10520
rect 14332 10480 14338 10492
rect 15381 10489 15393 10492
rect 15427 10489 15439 10523
rect 15381 10483 15439 10489
rect 7975 10424 8064 10452
rect 7975 10421 7987 10424
rect 7929 10415 7987 10421
rect 8662 10412 8668 10464
rect 8720 10452 8726 10464
rect 10965 10455 11023 10461
rect 10965 10452 10977 10455
rect 8720 10424 10977 10452
rect 8720 10412 8726 10424
rect 10965 10421 10977 10424
rect 11011 10452 11023 10455
rect 11146 10452 11152 10464
rect 11011 10424 11152 10452
rect 11011 10421 11023 10424
rect 10965 10415 11023 10421
rect 11146 10412 11152 10424
rect 11204 10412 11210 10464
rect 11514 10452 11520 10464
rect 11475 10424 11520 10452
rect 11514 10412 11520 10424
rect 11572 10412 11578 10464
rect 11885 10455 11943 10461
rect 11885 10421 11897 10455
rect 11931 10452 11943 10455
rect 11974 10452 11980 10464
rect 11931 10424 11980 10452
rect 11931 10421 11943 10424
rect 11885 10415 11943 10421
rect 11974 10412 11980 10424
rect 12032 10412 12038 10464
rect 15488 10452 15516 10560
rect 16666 10548 16672 10560
rect 16724 10548 16730 10600
rect 15841 10523 15899 10529
rect 15841 10489 15853 10523
rect 15887 10520 15899 10523
rect 16868 10520 16896 10619
rect 17494 10616 17500 10668
rect 17552 10656 17558 10668
rect 18121 10659 18179 10665
rect 18121 10656 18133 10659
rect 17552 10628 18133 10656
rect 17552 10616 17558 10628
rect 18121 10625 18133 10628
rect 18167 10625 18179 10659
rect 18121 10619 18179 10625
rect 19705 10659 19763 10665
rect 19705 10625 19717 10659
rect 19751 10656 19763 10659
rect 20180 10656 20208 10696
rect 20622 10684 20628 10696
rect 20680 10724 20686 10736
rect 21085 10727 21143 10733
rect 21085 10724 21097 10727
rect 20680 10696 21097 10724
rect 20680 10684 20686 10696
rect 21085 10693 21097 10696
rect 21131 10693 21143 10727
rect 21744 10724 21772 10764
rect 22094 10752 22100 10804
rect 22152 10792 22158 10804
rect 22554 10792 22560 10804
rect 22152 10764 22560 10792
rect 22152 10752 22158 10764
rect 22554 10752 22560 10764
rect 22612 10792 22618 10804
rect 23753 10795 23811 10801
rect 22612 10764 23704 10792
rect 22612 10752 22618 10764
rect 23477 10727 23535 10733
rect 21744 10696 23336 10724
rect 21085 10687 21143 10693
rect 19751 10628 20208 10656
rect 20533 10659 20591 10665
rect 19751 10625 19763 10628
rect 19705 10619 19763 10625
rect 20533 10625 20545 10659
rect 20579 10656 20591 10659
rect 20901 10659 20959 10665
rect 20901 10656 20913 10659
rect 20579 10628 20913 10656
rect 20579 10625 20591 10628
rect 20533 10619 20591 10625
rect 20901 10625 20913 10628
rect 20947 10625 20959 10659
rect 20901 10619 20959 10625
rect 21174 10616 21180 10668
rect 21232 10656 21238 10668
rect 22005 10659 22063 10665
rect 21232 10628 21277 10656
rect 21232 10616 21238 10628
rect 22005 10625 22017 10659
rect 22051 10656 22063 10659
rect 22094 10656 22100 10668
rect 22051 10628 22100 10656
rect 22051 10625 22063 10628
rect 22005 10619 22063 10625
rect 22094 10616 22100 10628
rect 22152 10616 22158 10668
rect 22278 10616 22284 10668
rect 22336 10656 22342 10668
rect 22462 10656 22468 10668
rect 22336 10628 22381 10656
rect 22423 10628 22468 10656
rect 22336 10616 22342 10628
rect 22462 10616 22468 10628
rect 22520 10616 22526 10668
rect 23198 10656 23204 10668
rect 22940 10628 23204 10656
rect 17678 10548 17684 10600
rect 17736 10588 17742 10600
rect 17865 10591 17923 10597
rect 17865 10588 17877 10591
rect 17736 10560 17877 10588
rect 17736 10548 17742 10560
rect 17865 10557 17877 10560
rect 17911 10557 17923 10591
rect 17865 10551 17923 10557
rect 19334 10548 19340 10600
rect 19392 10588 19398 10600
rect 22940 10588 22968 10628
rect 23198 10616 23204 10628
rect 23256 10616 23262 10668
rect 23308 10656 23336 10696
rect 23477 10693 23489 10727
rect 23523 10724 23535 10727
rect 23676 10724 23704 10764
rect 23753 10761 23765 10795
rect 23799 10792 23811 10795
rect 23934 10792 23940 10804
rect 23799 10764 23940 10792
rect 23799 10761 23811 10764
rect 23753 10755 23811 10761
rect 23934 10752 23940 10764
rect 23992 10752 23998 10804
rect 25501 10795 25559 10801
rect 25501 10761 25513 10795
rect 25547 10792 25559 10795
rect 25682 10792 25688 10804
rect 25547 10764 25688 10792
rect 25547 10761 25559 10764
rect 25501 10755 25559 10761
rect 25682 10752 25688 10764
rect 25740 10752 25746 10804
rect 26142 10752 26148 10804
rect 26200 10752 26206 10804
rect 28077 10795 28135 10801
rect 28077 10761 28089 10795
rect 28123 10792 28135 10795
rect 29822 10792 29828 10804
rect 28123 10764 29828 10792
rect 28123 10761 28135 10764
rect 28077 10755 28135 10761
rect 29822 10752 29828 10764
rect 29880 10752 29886 10804
rect 30101 10795 30159 10801
rect 30101 10761 30113 10795
rect 30147 10792 30159 10795
rect 30190 10792 30196 10804
rect 30147 10764 30196 10792
rect 30147 10761 30159 10764
rect 30101 10755 30159 10761
rect 30190 10752 30196 10764
rect 30248 10752 30254 10804
rect 30561 10795 30619 10801
rect 30561 10761 30573 10795
rect 30607 10792 30619 10795
rect 30834 10792 30840 10804
rect 30607 10764 30840 10792
rect 30607 10761 30619 10764
rect 30561 10755 30619 10761
rect 30834 10752 30840 10764
rect 30892 10752 30898 10804
rect 24026 10724 24032 10736
rect 23523 10696 23612 10724
rect 23676 10696 24032 10724
rect 23523 10693 23535 10696
rect 23477 10687 23535 10693
rect 23584 10656 23612 10696
rect 24026 10684 24032 10696
rect 24084 10684 24090 10736
rect 26160 10724 26188 10752
rect 25700 10696 27200 10724
rect 23750 10656 23756 10668
rect 23308 10628 23500 10656
rect 23584 10628 23756 10656
rect 23106 10588 23112 10600
rect 19392 10560 22968 10588
rect 23067 10560 23112 10588
rect 19392 10548 19398 10560
rect 23106 10548 23112 10560
rect 23164 10548 23170 10600
rect 23290 10548 23296 10600
rect 23348 10588 23354 10600
rect 23385 10591 23443 10597
rect 23385 10588 23397 10591
rect 23348 10560 23397 10588
rect 23348 10548 23354 10560
rect 23385 10557 23397 10560
rect 23431 10557 23443 10591
rect 23472 10588 23500 10628
rect 23750 10616 23756 10628
rect 23808 10616 23814 10668
rect 23842 10616 23848 10668
rect 23900 10656 23906 10668
rect 25700 10665 25728 10696
rect 24397 10659 24455 10665
rect 24397 10656 24409 10659
rect 23900 10628 24409 10656
rect 23900 10616 23906 10628
rect 24397 10625 24409 10628
rect 24443 10625 24455 10659
rect 24397 10619 24455 10625
rect 25685 10659 25743 10665
rect 25685 10625 25697 10659
rect 25731 10625 25743 10659
rect 25685 10619 25743 10625
rect 25958 10616 25964 10668
rect 26016 10660 26022 10668
rect 26016 10656 26087 10660
rect 26145 10659 26203 10665
rect 26016 10628 26109 10656
rect 26016 10616 26022 10628
rect 23594 10591 23652 10597
rect 23594 10588 23606 10591
rect 23472 10560 23606 10588
rect 23385 10551 23443 10557
rect 23594 10557 23606 10560
rect 23640 10557 23652 10591
rect 23594 10551 23652 10557
rect 24673 10591 24731 10597
rect 24673 10557 24685 10591
rect 24719 10588 24731 10591
rect 26059 10588 26087 10628
rect 26145 10625 26157 10659
rect 26191 10656 26203 10659
rect 26234 10656 26240 10668
rect 26191 10628 26240 10656
rect 26191 10625 26203 10628
rect 26145 10619 26203 10625
rect 26234 10616 26240 10628
rect 26292 10616 26298 10668
rect 27172 10665 27200 10696
rect 27246 10684 27252 10736
rect 27304 10724 27310 10736
rect 28994 10733 29000 10736
rect 28988 10724 29000 10733
rect 27304 10696 27660 10724
rect 28955 10696 29000 10724
rect 27304 10684 27310 10696
rect 27157 10659 27215 10665
rect 27157 10625 27169 10659
rect 27203 10625 27215 10659
rect 27430 10656 27436 10668
rect 27391 10628 27436 10656
rect 27157 10619 27215 10625
rect 27430 10616 27436 10628
rect 27488 10616 27494 10668
rect 27632 10665 27660 10696
rect 28988 10687 29000 10696
rect 28994 10684 29000 10687
rect 29052 10684 29058 10736
rect 29178 10684 29184 10736
rect 29236 10684 29242 10736
rect 29638 10684 29644 10736
rect 29696 10724 29702 10736
rect 29696 10696 31064 10724
rect 29696 10684 29702 10696
rect 27617 10659 27675 10665
rect 27617 10625 27629 10659
rect 27663 10625 27675 10659
rect 27617 10619 27675 10625
rect 28261 10659 28319 10665
rect 28261 10625 28273 10659
rect 28307 10625 28319 10659
rect 29196 10656 29224 10684
rect 28261 10619 28319 10625
rect 28736 10628 29224 10656
rect 27448 10588 27476 10616
rect 24719 10560 25912 10588
rect 26059 10560 27476 10588
rect 24719 10557 24731 10560
rect 24673 10551 24731 10557
rect 20717 10523 20775 10529
rect 15887 10492 16896 10520
rect 18984 10492 20576 10520
rect 15887 10489 15899 10492
rect 15841 10483 15899 10489
rect 18984 10452 19012 10492
rect 15488 10424 19012 10452
rect 19245 10455 19303 10461
rect 19245 10421 19257 10455
rect 19291 10452 19303 10455
rect 20073 10455 20131 10461
rect 20073 10452 20085 10455
rect 19291 10424 20085 10452
rect 19291 10421 19303 10424
rect 19245 10415 19303 10421
rect 20073 10421 20085 10424
rect 20119 10452 20131 10455
rect 20438 10452 20444 10464
rect 20119 10424 20444 10452
rect 20119 10421 20131 10424
rect 20073 10415 20131 10421
rect 20438 10412 20444 10424
rect 20496 10412 20502 10464
rect 20548 10452 20576 10492
rect 20717 10489 20729 10523
rect 20763 10520 20775 10523
rect 24946 10520 24952 10532
rect 20763 10492 24952 10520
rect 20763 10489 20775 10492
rect 20717 10483 20775 10489
rect 24946 10480 24952 10492
rect 25004 10480 25010 10532
rect 25884 10520 25912 10560
rect 27522 10548 27528 10600
rect 27580 10588 27586 10600
rect 28276 10588 28304 10619
rect 28736 10597 28764 10628
rect 29730 10616 29736 10668
rect 29788 10656 29794 10668
rect 31036 10665 31064 10696
rect 30745 10659 30803 10665
rect 30745 10656 30757 10659
rect 29788 10628 30757 10656
rect 29788 10616 29794 10628
rect 30745 10625 30757 10628
rect 30791 10625 30803 10659
rect 30745 10619 30803 10625
rect 31021 10659 31079 10665
rect 31021 10625 31033 10659
rect 31067 10625 31079 10659
rect 31202 10656 31208 10668
rect 31163 10628 31208 10656
rect 31021 10619 31079 10625
rect 31202 10616 31208 10628
rect 31260 10616 31266 10668
rect 27580 10560 28304 10588
rect 28721 10591 28779 10597
rect 27580 10548 27586 10560
rect 28721 10557 28733 10591
rect 28767 10557 28779 10591
rect 28721 10551 28779 10557
rect 26234 10520 26240 10532
rect 25884 10492 26240 10520
rect 26234 10480 26240 10492
rect 26292 10480 26298 10532
rect 21542 10452 21548 10464
rect 20548 10424 21548 10452
rect 21542 10412 21548 10424
rect 21600 10412 21606 10464
rect 21818 10452 21824 10464
rect 21779 10424 21824 10452
rect 21818 10412 21824 10424
rect 21876 10412 21882 10464
rect 24210 10452 24216 10464
rect 24171 10424 24216 10452
rect 24210 10412 24216 10424
rect 24268 10412 24274 10464
rect 24581 10455 24639 10461
rect 24581 10421 24593 10455
rect 24627 10452 24639 10455
rect 25866 10452 25872 10464
rect 24627 10424 25872 10452
rect 24627 10421 24639 10424
rect 24581 10415 24639 10421
rect 25866 10412 25872 10424
rect 25924 10412 25930 10464
rect 26326 10412 26332 10464
rect 26384 10452 26390 10464
rect 26973 10455 27031 10461
rect 26973 10452 26985 10455
rect 26384 10424 26985 10452
rect 26384 10412 26390 10424
rect 26973 10421 26985 10424
rect 27019 10421 27031 10455
rect 26973 10415 27031 10421
rect 1104 10362 32016 10384
rect 1104 10310 2136 10362
rect 2188 10310 12440 10362
rect 12492 10310 22744 10362
rect 22796 10310 32016 10362
rect 1104 10288 32016 10310
rect 1118 10208 1124 10260
rect 1176 10248 1182 10260
rect 1176 10220 2360 10248
rect 1176 10208 1182 10220
rect 2332 10180 2360 10220
rect 3050 10208 3056 10260
rect 3108 10248 3114 10260
rect 3878 10248 3884 10260
rect 3108 10220 3884 10248
rect 3108 10208 3114 10220
rect 3878 10208 3884 10220
rect 3936 10208 3942 10260
rect 3988 10220 5212 10248
rect 3988 10180 4016 10220
rect 2332 10152 4016 10180
rect 5184 10112 5212 10220
rect 5442 10208 5448 10260
rect 5500 10248 5506 10260
rect 5537 10251 5595 10257
rect 5537 10248 5549 10251
rect 5500 10220 5549 10248
rect 5500 10208 5506 10220
rect 5537 10217 5549 10220
rect 5583 10217 5595 10251
rect 5537 10211 5595 10217
rect 6454 10208 6460 10260
rect 6512 10248 6518 10260
rect 6733 10251 6791 10257
rect 6733 10248 6745 10251
rect 6512 10220 6745 10248
rect 6512 10208 6518 10220
rect 6733 10217 6745 10220
rect 6779 10217 6791 10251
rect 6733 10211 6791 10217
rect 7193 10251 7251 10257
rect 7193 10217 7205 10251
rect 7239 10248 7251 10251
rect 7239 10220 8156 10248
rect 7239 10217 7251 10220
rect 7193 10211 7251 10217
rect 6270 10140 6276 10192
rect 6328 10180 6334 10192
rect 6549 10183 6607 10189
rect 6549 10180 6561 10183
rect 6328 10152 6561 10180
rect 6328 10140 6334 10152
rect 6549 10149 6561 10152
rect 6595 10149 6607 10183
rect 6549 10143 6607 10149
rect 7650 10140 7656 10192
rect 7708 10180 7714 10192
rect 7837 10183 7895 10189
rect 7837 10180 7849 10183
rect 7708 10152 7849 10180
rect 7708 10140 7714 10152
rect 7837 10149 7849 10152
rect 7883 10149 7895 10183
rect 8128 10180 8156 10220
rect 8202 10208 8208 10260
rect 8260 10248 8266 10260
rect 8389 10251 8447 10257
rect 8260 10220 8305 10248
rect 8260 10208 8266 10220
rect 8389 10217 8401 10251
rect 8435 10248 8447 10251
rect 8938 10248 8944 10260
rect 8435 10220 8944 10248
rect 8435 10217 8447 10220
rect 8389 10211 8447 10217
rect 8938 10208 8944 10220
rect 8996 10208 9002 10260
rect 11146 10248 11152 10260
rect 9784 10220 10732 10248
rect 11107 10220 11152 10248
rect 9784 10180 9812 10220
rect 8128 10152 9812 10180
rect 10704 10180 10732 10220
rect 11146 10208 11152 10220
rect 11204 10208 11210 10260
rect 13078 10208 13084 10260
rect 13136 10248 13142 10260
rect 13173 10251 13231 10257
rect 13173 10248 13185 10251
rect 13136 10220 13185 10248
rect 13136 10208 13142 10220
rect 13173 10217 13185 10220
rect 13219 10217 13231 10251
rect 13173 10211 13231 10217
rect 16022 10208 16028 10260
rect 16080 10248 16086 10260
rect 18049 10251 18107 10257
rect 16080 10220 17954 10248
rect 16080 10208 16086 10220
rect 11238 10180 11244 10192
rect 10704 10152 11244 10180
rect 7837 10143 7895 10149
rect 11238 10140 11244 10152
rect 11296 10140 11302 10192
rect 16666 10140 16672 10192
rect 16724 10140 16730 10192
rect 17926 10180 17954 10220
rect 18049 10217 18061 10251
rect 18095 10248 18107 10251
rect 18322 10248 18328 10260
rect 18095 10220 18328 10248
rect 18095 10217 18107 10220
rect 18049 10211 18107 10217
rect 18322 10208 18328 10220
rect 18380 10208 18386 10260
rect 21269 10251 21327 10257
rect 21269 10217 21281 10251
rect 21315 10248 21327 10251
rect 23842 10248 23848 10260
rect 21315 10220 23848 10248
rect 21315 10217 21327 10220
rect 21269 10211 21327 10217
rect 23842 10208 23848 10220
rect 23900 10208 23906 10260
rect 24026 10208 24032 10260
rect 24084 10248 24090 10260
rect 25958 10248 25964 10260
rect 24084 10220 25964 10248
rect 24084 10208 24090 10220
rect 25958 10208 25964 10220
rect 26016 10208 26022 10260
rect 27246 10208 27252 10260
rect 27304 10248 27310 10260
rect 27617 10251 27675 10257
rect 27617 10248 27629 10251
rect 27304 10220 27629 10248
rect 27304 10208 27310 10220
rect 27617 10217 27629 10220
rect 27663 10217 27675 10251
rect 31202 10248 31208 10260
rect 31163 10220 31208 10248
rect 27617 10211 27675 10217
rect 31202 10208 31208 10220
rect 31260 10208 31266 10260
rect 18506 10180 18512 10192
rect 17926 10152 18512 10180
rect 18506 10140 18512 10152
rect 18564 10180 18570 10192
rect 18601 10183 18659 10189
rect 18601 10180 18613 10183
rect 18564 10152 18613 10180
rect 18564 10140 18570 10152
rect 18601 10149 18613 10152
rect 18647 10149 18659 10183
rect 18601 10143 18659 10149
rect 20257 10183 20315 10189
rect 20257 10149 20269 10183
rect 20303 10149 20315 10183
rect 21910 10180 21916 10192
rect 20257 10143 20315 10149
rect 20732 10152 21916 10180
rect 9214 10112 9220 10124
rect 5184 10084 9220 10112
rect 9214 10072 9220 10084
rect 9272 10072 9278 10124
rect 14274 10072 14280 10124
rect 14332 10112 14338 10124
rect 16301 10115 16359 10121
rect 16301 10112 16313 10115
rect 14332 10084 16313 10112
rect 14332 10072 14338 10084
rect 16301 10081 16313 10084
rect 16347 10081 16359 10115
rect 16684 10112 16712 10140
rect 20272 10112 20300 10143
rect 16684 10084 16804 10112
rect 16301 10075 16359 10081
rect 1397 10047 1455 10053
rect 1397 10013 1409 10047
rect 1443 10044 1455 10047
rect 2682 10044 2688 10056
rect 1443 10016 2688 10044
rect 1443 10013 1455 10016
rect 1397 10007 1455 10013
rect 2682 10004 2688 10016
rect 2740 10044 2746 10056
rect 4154 10044 4160 10056
rect 2740 10016 4160 10044
rect 2740 10004 2746 10016
rect 4154 10004 4160 10016
rect 4212 10004 4218 10056
rect 5994 10004 6000 10056
rect 6052 10044 6058 10056
rect 6730 10044 6736 10056
rect 6052 10016 6736 10044
rect 6052 10004 6058 10016
rect 6730 10004 6736 10016
rect 6788 10044 6794 10056
rect 7374 10044 7380 10056
rect 6788 10016 7236 10044
rect 7335 10016 7380 10044
rect 6788 10004 6794 10016
rect 0 9976 800 9990
rect 1664 9979 1722 9985
rect 0 9948 888 9976
rect 0 9934 800 9948
rect 860 9840 888 9948
rect 1664 9945 1676 9979
rect 1710 9976 1722 9979
rect 1762 9976 1768 9988
rect 1710 9948 1768 9976
rect 1710 9945 1722 9948
rect 1664 9939 1722 9945
rect 1762 9936 1768 9948
rect 1820 9936 1826 9988
rect 4424 9979 4482 9985
rect 4424 9945 4436 9979
rect 4470 9976 4482 9979
rect 6273 9979 6331 9985
rect 4470 9948 6040 9976
rect 4470 9945 4482 9948
rect 4424 9939 4482 9945
rect 6012 9920 6040 9948
rect 6273 9945 6285 9979
rect 6319 9976 6331 9979
rect 7098 9976 7104 9988
rect 6319 9948 7104 9976
rect 6319 9945 6331 9948
rect 6273 9939 6331 9945
rect 7098 9936 7104 9948
rect 7156 9936 7162 9988
rect 7208 9976 7236 10016
rect 7374 10004 7380 10016
rect 7432 10004 7438 10056
rect 9769 10047 9827 10053
rect 7852 10016 9251 10044
rect 7852 9976 7880 10016
rect 7208 9948 7880 9976
rect 8205 9979 8263 9985
rect 8205 9945 8217 9979
rect 8251 9976 8263 9979
rect 8386 9976 8392 9988
rect 8251 9948 8392 9976
rect 8251 9945 8263 9948
rect 8205 9939 8263 9945
rect 8386 9936 8392 9948
rect 8444 9936 8450 9988
rect 8754 9936 8760 9988
rect 8812 9976 8818 9988
rect 8938 9976 8944 9988
rect 8812 9948 8944 9976
rect 8812 9936 8818 9948
rect 8938 9936 8944 9948
rect 8996 9976 9002 9988
rect 9125 9979 9183 9985
rect 9125 9976 9137 9979
rect 8996 9948 9137 9976
rect 8996 9936 9002 9948
rect 9125 9945 9137 9948
rect 9171 9945 9183 9979
rect 9223 9976 9251 10016
rect 9769 10013 9781 10047
rect 9815 10044 9827 10047
rect 11790 10044 11796 10056
rect 9815 10016 11796 10044
rect 9815 10013 9827 10016
rect 9769 10007 9827 10013
rect 11790 10004 11796 10016
rect 11848 10004 11854 10056
rect 16669 10047 16727 10053
rect 16669 10044 16681 10047
rect 16040 10016 16681 10044
rect 9858 9976 9864 9988
rect 9223 9948 9864 9976
rect 9125 9939 9183 9945
rect 9858 9936 9864 9948
rect 9916 9936 9922 9988
rect 10036 9979 10094 9985
rect 10036 9945 10048 9979
rect 10082 9976 10094 9979
rect 11514 9976 11520 9988
rect 10082 9948 11520 9976
rect 10082 9945 10094 9948
rect 10036 9939 10094 9945
rect 11514 9936 11520 9948
rect 11572 9936 11578 9988
rect 12066 9985 12072 9988
rect 12060 9939 12072 9985
rect 12124 9976 12130 9988
rect 14458 9976 14464 9988
rect 12124 9948 12160 9976
rect 14419 9948 14464 9976
rect 12066 9936 12072 9939
rect 12124 9936 12130 9948
rect 14458 9936 14464 9948
rect 14516 9936 14522 9988
rect 2222 9868 2228 9920
rect 2280 9908 2286 9920
rect 2777 9911 2835 9917
rect 2777 9908 2789 9911
rect 2280 9880 2789 9908
rect 2280 9868 2286 9880
rect 2777 9877 2789 9880
rect 2823 9877 2835 9911
rect 2777 9871 2835 9877
rect 3418 9868 3424 9920
rect 3476 9908 3482 9920
rect 3786 9908 3792 9920
rect 3476 9880 3792 9908
rect 3476 9868 3482 9880
rect 3786 9868 3792 9880
rect 3844 9868 3850 9920
rect 5994 9868 6000 9920
rect 6052 9868 6058 9920
rect 7190 9868 7196 9920
rect 7248 9908 7254 9920
rect 8294 9908 8300 9920
rect 7248 9880 8300 9908
rect 7248 9868 7254 9880
rect 8294 9868 8300 9880
rect 8352 9868 8358 9920
rect 8846 9868 8852 9920
rect 8904 9908 8910 9920
rect 9217 9911 9275 9917
rect 9217 9908 9229 9911
rect 8904 9880 9229 9908
rect 8904 9868 8910 9880
rect 9217 9877 9229 9880
rect 9263 9877 9275 9911
rect 9217 9871 9275 9877
rect 14090 9868 14096 9920
rect 14148 9908 14154 9920
rect 15749 9911 15807 9917
rect 15749 9908 15761 9911
rect 14148 9880 15761 9908
rect 14148 9868 14154 9880
rect 15749 9877 15761 9880
rect 15795 9908 15807 9911
rect 16040 9908 16068 10016
rect 16669 10013 16681 10016
rect 16715 10013 16727 10047
rect 16776 10044 16804 10084
rect 17926 10084 20300 10112
rect 16925 10047 16983 10053
rect 16925 10044 16937 10047
rect 16776 10016 16937 10044
rect 16669 10007 16727 10013
rect 16925 10013 16937 10016
rect 16971 10013 16983 10047
rect 16925 10007 16983 10013
rect 16301 9979 16359 9985
rect 16301 9945 16313 9979
rect 16347 9976 16359 9979
rect 17926 9976 17954 10084
rect 18322 10004 18328 10056
rect 18380 10044 18386 10056
rect 18509 10047 18567 10053
rect 18509 10044 18521 10047
rect 18380 10016 18521 10044
rect 18380 10004 18386 10016
rect 18509 10013 18521 10016
rect 18555 10013 18567 10047
rect 18509 10007 18567 10013
rect 18598 10004 18604 10056
rect 18656 10044 18662 10056
rect 20073 10047 20131 10053
rect 20073 10044 20085 10047
rect 18656 10016 20085 10044
rect 18656 10004 18662 10016
rect 20073 10013 20085 10016
rect 20119 10044 20131 10047
rect 20732 10044 20760 10152
rect 21910 10140 21916 10152
rect 21968 10140 21974 10192
rect 20806 10072 20812 10124
rect 20864 10112 20870 10124
rect 22005 10115 22063 10121
rect 22005 10112 22017 10115
rect 20864 10084 22017 10112
rect 20864 10072 20870 10084
rect 22005 10081 22017 10084
rect 22051 10081 22063 10115
rect 22005 10075 22063 10081
rect 20119 10016 20760 10044
rect 20119 10013 20131 10016
rect 20073 10007 20131 10013
rect 21082 10004 21088 10056
rect 21140 10044 21146 10056
rect 21269 10047 21327 10053
rect 21269 10044 21281 10047
rect 21140 10016 21281 10044
rect 21140 10004 21146 10016
rect 21269 10013 21281 10016
rect 21315 10013 21327 10047
rect 21269 10007 21327 10013
rect 21545 10047 21603 10053
rect 21545 10013 21557 10047
rect 21591 10044 21603 10047
rect 21634 10044 21640 10056
rect 21591 10016 21640 10044
rect 21591 10013 21603 10016
rect 21545 10007 21603 10013
rect 21634 10004 21640 10016
rect 21692 10004 21698 10056
rect 23658 10044 23664 10056
rect 22204 10016 23664 10044
rect 19334 9976 19340 9988
rect 16347 9948 17954 9976
rect 19295 9948 19340 9976
rect 16347 9945 16359 9948
rect 16301 9939 16359 9945
rect 19334 9936 19340 9948
rect 19392 9936 19398 9988
rect 21453 9979 21511 9985
rect 21453 9945 21465 9979
rect 21499 9976 21511 9979
rect 22204 9976 22232 10016
rect 23658 10004 23664 10016
rect 23716 10004 23722 10056
rect 24397 10047 24455 10053
rect 24397 10013 24409 10047
rect 24443 10044 24455 10047
rect 26237 10047 26295 10053
rect 26237 10044 26249 10047
rect 24443 10016 26249 10044
rect 24443 10013 24455 10016
rect 24397 10007 24455 10013
rect 26237 10013 26249 10016
rect 26283 10044 26295 10047
rect 26786 10044 26792 10056
rect 26283 10016 26792 10044
rect 26283 10013 26295 10016
rect 26237 10007 26295 10013
rect 26786 10004 26792 10016
rect 26844 10004 26850 10056
rect 27522 10004 27528 10056
rect 27580 10044 27586 10056
rect 28813 10047 28871 10053
rect 28813 10044 28825 10047
rect 27580 10016 28825 10044
rect 27580 10004 27586 10016
rect 28813 10013 28825 10016
rect 28859 10013 28871 10047
rect 28813 10007 28871 10013
rect 29178 10004 29184 10056
rect 29236 10044 29242 10056
rect 30098 10053 30104 10056
rect 29825 10047 29883 10053
rect 29825 10044 29837 10047
rect 29236 10016 29837 10044
rect 29236 10004 29242 10016
rect 29825 10013 29837 10016
rect 29871 10013 29883 10047
rect 30092 10044 30104 10053
rect 30059 10016 30104 10044
rect 29825 10007 29883 10013
rect 30092 10007 30104 10016
rect 30098 10004 30104 10007
rect 30156 10004 30162 10056
rect 21499 9948 22232 9976
rect 22272 9979 22330 9985
rect 21499 9945 21511 9948
rect 21453 9939 21511 9945
rect 22272 9945 22284 9979
rect 22318 9976 22330 9979
rect 22646 9976 22652 9988
rect 22318 9948 22652 9976
rect 22318 9945 22330 9948
rect 22272 9939 22330 9945
rect 22646 9936 22652 9948
rect 22704 9936 22710 9988
rect 23290 9936 23296 9988
rect 23348 9976 23354 9988
rect 23348 9948 23500 9976
rect 23348 9936 23354 9948
rect 15795 9880 16068 9908
rect 15795 9877 15807 9880
rect 15749 9871 15807 9877
rect 16114 9868 16120 9920
rect 16172 9908 16178 9920
rect 19429 9911 19487 9917
rect 19429 9908 19441 9911
rect 16172 9880 19441 9908
rect 16172 9868 16178 9880
rect 19429 9877 19441 9880
rect 19475 9908 19487 9911
rect 19518 9908 19524 9920
rect 19475 9880 19524 9908
rect 19475 9877 19487 9880
rect 19429 9871 19487 9877
rect 19518 9868 19524 9880
rect 19576 9868 19582 9920
rect 22462 9868 22468 9920
rect 22520 9908 22526 9920
rect 23106 9908 23112 9920
rect 22520 9880 23112 9908
rect 22520 9868 22526 9880
rect 23106 9868 23112 9880
rect 23164 9908 23170 9920
rect 23385 9911 23443 9917
rect 23385 9908 23397 9911
rect 23164 9880 23397 9908
rect 23164 9868 23170 9880
rect 23385 9877 23397 9880
rect 23431 9877 23443 9911
rect 23472 9908 23500 9948
rect 24210 9936 24216 9988
rect 24268 9976 24274 9988
rect 24642 9979 24700 9985
rect 24642 9976 24654 9979
rect 24268 9948 24654 9976
rect 24268 9936 24274 9948
rect 24642 9945 24654 9948
rect 24688 9945 24700 9979
rect 24642 9939 24700 9945
rect 26142 9936 26148 9988
rect 26200 9976 26206 9988
rect 26482 9979 26540 9985
rect 26482 9976 26494 9979
rect 26200 9948 26494 9976
rect 26200 9936 26206 9948
rect 26482 9945 26494 9948
rect 26528 9945 26540 9979
rect 32320 9976 33120 9990
rect 26482 9939 26540 9945
rect 26589 9948 33120 9976
rect 25777 9911 25835 9917
rect 25777 9908 25789 9911
rect 23472 9880 25789 9908
rect 23385 9871 23443 9877
rect 25777 9877 25789 9880
rect 25823 9877 25835 9911
rect 25777 9871 25835 9877
rect 26234 9868 26240 9920
rect 26292 9908 26298 9920
rect 26589 9908 26617 9948
rect 32320 9934 33120 9948
rect 26292 9880 26617 9908
rect 26292 9868 26298 9880
rect 28534 9868 28540 9920
rect 28592 9908 28598 9920
rect 28629 9911 28687 9917
rect 28629 9908 28641 9911
rect 28592 9880 28641 9908
rect 28592 9868 28598 9880
rect 28629 9877 28641 9880
rect 28675 9908 28687 9911
rect 29086 9908 29092 9920
rect 28675 9880 29092 9908
rect 28675 9877 28687 9880
rect 28629 9871 28687 9877
rect 29086 9868 29092 9880
rect 29144 9868 29150 9920
rect 768 9812 888 9840
rect 1104 9818 32016 9840
rect 768 9704 796 9812
rect 1104 9766 7288 9818
rect 7340 9766 17592 9818
rect 17644 9766 27896 9818
rect 27948 9766 32016 9818
rect 1104 9744 32016 9766
rect 3694 9704 3700 9716
rect 768 9676 3700 9704
rect 3694 9664 3700 9676
rect 3752 9664 3758 9716
rect 3878 9664 3884 9716
rect 3936 9704 3942 9716
rect 5537 9707 5595 9713
rect 5537 9704 5549 9707
rect 3936 9676 5549 9704
rect 3936 9664 3942 9676
rect 5537 9673 5549 9676
rect 5583 9704 5595 9707
rect 6638 9704 6644 9716
rect 5583 9676 6644 9704
rect 5583 9673 5595 9676
rect 5537 9667 5595 9673
rect 6638 9664 6644 9676
rect 6696 9664 6702 9716
rect 7650 9664 7656 9716
rect 7708 9704 7714 9716
rect 7708 9676 8984 9704
rect 7708 9664 7714 9676
rect 1489 9639 1547 9645
rect 1489 9605 1501 9639
rect 1535 9636 1547 9639
rect 1762 9636 1768 9648
rect 1535 9608 1768 9636
rect 1535 9605 1547 9608
rect 1489 9599 1547 9605
rect 1762 9596 1768 9608
rect 1820 9636 1826 9648
rect 2314 9636 2320 9648
rect 1820 9608 2320 9636
rect 1820 9596 1826 9608
rect 2314 9596 2320 9608
rect 2372 9596 2378 9648
rect 4706 9636 4712 9648
rect 3528 9608 4712 9636
rect 1394 9568 1400 9580
rect 1355 9540 1400 9568
rect 1394 9528 1400 9540
rect 1452 9528 1458 9580
rect 2041 9571 2099 9577
rect 2041 9537 2053 9571
rect 2087 9568 2099 9571
rect 2222 9568 2228 9580
rect 2087 9540 2228 9568
rect 2087 9537 2099 9540
rect 2041 9531 2099 9537
rect 2222 9528 2228 9540
rect 2280 9528 2286 9580
rect 2682 9568 2688 9580
rect 2332 9540 2688 9568
rect 2332 9512 2360 9540
rect 2682 9528 2688 9540
rect 2740 9528 2746 9580
rect 3528 9577 3556 9608
rect 4706 9596 4712 9608
rect 4764 9596 4770 9648
rect 4890 9636 4896 9648
rect 4851 9608 4896 9636
rect 4890 9596 4896 9608
rect 4948 9596 4954 9648
rect 5184 9608 6684 9636
rect 3513 9571 3571 9577
rect 3513 9537 3525 9571
rect 3559 9537 3571 9571
rect 3513 9531 3571 9537
rect 4065 9571 4123 9577
rect 4065 9537 4077 9571
rect 4111 9568 4123 9571
rect 4522 9568 4528 9580
rect 4111 9540 4528 9568
rect 4111 9537 4123 9540
rect 4065 9531 4123 9537
rect 4522 9528 4528 9540
rect 4580 9528 4586 9580
rect 5074 9568 5080 9580
rect 5035 9540 5080 9568
rect 5074 9528 5080 9540
rect 5132 9528 5138 9580
rect 2314 9500 2320 9512
rect 2275 9472 2320 9500
rect 2314 9460 2320 9472
rect 2372 9460 2378 9512
rect 2406 9460 2412 9512
rect 2464 9500 2470 9512
rect 4157 9503 4215 9509
rect 4157 9500 4169 9503
rect 2464 9472 4169 9500
rect 2464 9460 2470 9472
rect 4157 9469 4169 9472
rect 4203 9469 4215 9503
rect 5184 9500 5212 9608
rect 5353 9571 5411 9577
rect 5353 9537 5365 9571
rect 5399 9568 5411 9571
rect 5718 9568 5724 9580
rect 5399 9540 5724 9568
rect 5399 9537 5411 9540
rect 5353 9531 5411 9537
rect 5718 9528 5724 9540
rect 5776 9568 5782 9580
rect 6546 9568 6552 9580
rect 5776 9540 6552 9568
rect 5776 9528 5782 9540
rect 6546 9528 6552 9540
rect 6604 9528 6610 9580
rect 6656 9568 6684 9608
rect 6822 9596 6828 9648
rect 6880 9636 6886 9648
rect 7193 9639 7251 9645
rect 7193 9636 7205 9639
rect 6880 9608 7205 9636
rect 6880 9596 6886 9608
rect 7193 9605 7205 9608
rect 7239 9605 7251 9639
rect 7193 9599 7251 9605
rect 8018 9596 8024 9648
rect 8076 9636 8082 9648
rect 8297 9639 8355 9645
rect 8297 9636 8309 9639
rect 8076 9608 8309 9636
rect 8076 9596 8082 9608
rect 8297 9605 8309 9608
rect 8343 9605 8355 9639
rect 8297 9599 8355 9605
rect 8386 9596 8392 9648
rect 8444 9636 8450 9648
rect 8757 9639 8815 9645
rect 8757 9636 8769 9639
rect 8444 9608 8769 9636
rect 8444 9596 8450 9608
rect 8757 9605 8769 9608
rect 8803 9605 8815 9639
rect 8757 9599 8815 9605
rect 8849 9639 8907 9645
rect 8849 9605 8861 9639
rect 8895 9636 8907 9639
rect 8956 9636 8984 9676
rect 9030 9664 9036 9716
rect 9088 9704 9094 9716
rect 9125 9707 9183 9713
rect 9125 9704 9137 9707
rect 9088 9676 9137 9704
rect 9088 9664 9094 9676
rect 9125 9673 9137 9676
rect 9171 9673 9183 9707
rect 9125 9667 9183 9673
rect 9214 9664 9220 9716
rect 9272 9704 9278 9716
rect 9272 9676 22600 9704
rect 9272 9664 9278 9676
rect 8895 9608 8984 9636
rect 9140 9608 9444 9636
rect 8895 9605 8907 9608
rect 8849 9599 8907 9605
rect 7101 9571 7159 9577
rect 7101 9568 7113 9571
rect 6656 9540 7113 9568
rect 7101 9537 7113 9540
rect 7147 9537 7159 9571
rect 8662 9568 8668 9580
rect 7101 9531 7159 9537
rect 7208 9540 8668 9568
rect 7208 9500 7236 9540
rect 8662 9528 8668 9540
rect 8720 9528 8726 9580
rect 7374 9500 7380 9512
rect 4157 9463 4215 9469
rect 5092 9472 5212 9500
rect 5460 9472 7236 9500
rect 7335 9472 7380 9500
rect 3602 9432 3608 9444
rect 3563 9404 3608 9432
rect 3602 9392 3608 9404
rect 3660 9392 3666 9444
rect 3970 9392 3976 9444
rect 4028 9432 4034 9444
rect 5092 9432 5120 9472
rect 5460 9432 5488 9472
rect 7374 9460 7380 9472
rect 7432 9460 7438 9512
rect 7558 9460 7564 9512
rect 7616 9500 7622 9512
rect 8389 9503 8447 9509
rect 8389 9500 8401 9503
rect 7616 9472 8401 9500
rect 7616 9460 7622 9472
rect 8389 9469 8401 9472
rect 8435 9469 8447 9503
rect 8389 9463 8447 9469
rect 8573 9503 8631 9509
rect 8573 9469 8585 9503
rect 8619 9500 8631 9503
rect 8754 9500 8760 9512
rect 8619 9472 8760 9500
rect 8619 9469 8631 9472
rect 8573 9463 8631 9469
rect 8754 9460 8760 9472
rect 8812 9460 8818 9512
rect 8849 9503 8907 9509
rect 8849 9469 8861 9503
rect 8895 9500 8907 9503
rect 9140 9500 9168 9608
rect 9416 9509 9444 9608
rect 9582 9596 9588 9648
rect 9640 9636 9646 9648
rect 13906 9636 13912 9648
rect 9640 9608 13912 9636
rect 9640 9596 9646 9608
rect 13906 9596 13912 9608
rect 13964 9596 13970 9648
rect 14366 9645 14372 9648
rect 14360 9599 14372 9645
rect 14424 9636 14430 9648
rect 21910 9636 21916 9648
rect 14424 9608 14460 9636
rect 14568 9608 21916 9636
rect 14366 9596 14372 9599
rect 14424 9596 14430 9608
rect 9674 9528 9680 9580
rect 9732 9528 9738 9580
rect 10689 9571 10747 9577
rect 10689 9537 10701 9571
rect 10735 9568 10747 9571
rect 10961 9571 11019 9577
rect 10735 9540 10824 9568
rect 10735 9537 10747 9540
rect 10689 9531 10747 9537
rect 10796 9534 10824 9540
rect 10961 9564 10973 9571
rect 11007 9564 11019 9571
rect 8895 9472 9168 9500
rect 9309 9503 9367 9509
rect 8895 9469 8907 9472
rect 8849 9463 8907 9469
rect 9309 9469 9321 9503
rect 9355 9469 9367 9503
rect 9309 9463 9367 9469
rect 9401 9503 9459 9509
rect 9401 9469 9413 9503
rect 9447 9469 9459 9503
rect 9401 9463 9459 9469
rect 9493 9503 9551 9509
rect 9493 9469 9505 9503
rect 9539 9469 9551 9503
rect 9493 9463 9551 9469
rect 9585 9503 9643 9509
rect 9585 9469 9597 9503
rect 9631 9500 9643 9503
rect 9692 9500 9720 9528
rect 10796 9512 10916 9534
rect 10961 9531 10968 9564
rect 10962 9512 10968 9531
rect 11020 9512 11026 9564
rect 11146 9528 11152 9580
rect 11204 9568 11210 9580
rect 11517 9571 11575 9577
rect 11517 9568 11529 9571
rect 11204 9540 11529 9568
rect 11204 9528 11210 9540
rect 11517 9537 11529 9540
rect 11563 9537 11575 9571
rect 11517 9531 11575 9537
rect 11606 9528 11612 9580
rect 11664 9568 11670 9580
rect 11701 9571 11759 9577
rect 11701 9568 11713 9571
rect 11664 9540 11713 9568
rect 11664 9528 11670 9540
rect 11701 9537 11713 9540
rect 11747 9537 11759 9571
rect 11701 9531 11759 9537
rect 11882 9528 11888 9580
rect 11940 9568 11946 9580
rect 11977 9571 12035 9577
rect 11977 9568 11989 9571
rect 11940 9540 11989 9568
rect 11940 9528 11946 9540
rect 11977 9537 11989 9540
rect 12023 9537 12035 9571
rect 12158 9568 12164 9580
rect 12119 9540 12164 9568
rect 11977 9531 12035 9537
rect 12158 9528 12164 9540
rect 12216 9528 12222 9580
rect 12986 9528 12992 9580
rect 13044 9568 13050 9580
rect 13265 9571 13323 9577
rect 13265 9568 13277 9571
rect 13044 9540 13277 9568
rect 13044 9528 13050 9540
rect 13265 9537 13277 9540
rect 13311 9537 13323 9571
rect 14090 9568 14096 9580
rect 14051 9540 14096 9568
rect 13265 9531 13323 9537
rect 14090 9528 14096 9540
rect 14148 9528 14154 9580
rect 14568 9568 14596 9608
rect 21910 9596 21916 9608
rect 21968 9596 21974 9648
rect 22572 9636 22600 9676
rect 22646 9664 22652 9716
rect 22704 9704 22710 9716
rect 22741 9707 22799 9713
rect 22741 9704 22753 9707
rect 22704 9676 22753 9704
rect 22704 9664 22710 9676
rect 22741 9673 22753 9676
rect 22787 9673 22799 9707
rect 26234 9704 26240 9716
rect 22741 9667 22799 9673
rect 22940 9676 26240 9704
rect 22940 9636 22968 9676
rect 26234 9664 26240 9676
rect 26292 9664 26298 9716
rect 26329 9707 26387 9713
rect 26329 9673 26341 9707
rect 26375 9704 26387 9707
rect 26418 9704 26424 9716
rect 26375 9676 26424 9704
rect 26375 9673 26387 9676
rect 26329 9667 26387 9673
rect 26418 9664 26424 9676
rect 26476 9664 26482 9716
rect 26694 9664 26700 9716
rect 26752 9704 26758 9716
rect 26752 9676 27660 9704
rect 26752 9664 26758 9676
rect 22572 9608 22968 9636
rect 23014 9596 23020 9648
rect 23072 9636 23078 9648
rect 24118 9636 24124 9648
rect 23072 9608 24124 9636
rect 23072 9596 23078 9608
rect 24118 9596 24124 9608
rect 24176 9596 24182 9648
rect 24489 9639 24547 9645
rect 24489 9605 24501 9639
rect 24535 9636 24547 9639
rect 24854 9636 24860 9648
rect 24535 9608 24860 9636
rect 24535 9605 24547 9608
rect 24489 9599 24547 9605
rect 24854 9596 24860 9608
rect 24912 9596 24918 9648
rect 25216 9639 25274 9645
rect 25216 9605 25228 9639
rect 25262 9636 25274 9639
rect 25498 9636 25504 9648
rect 25262 9608 25504 9636
rect 25262 9605 25274 9608
rect 25216 9599 25274 9605
rect 25498 9596 25504 9608
rect 25556 9596 25562 9648
rect 27632 9636 27660 9676
rect 29086 9636 29092 9648
rect 27632 9608 29092 9636
rect 14200 9540 14596 9568
rect 10318 9500 10324 9512
rect 9631 9472 10324 9500
rect 9631 9469 9643 9472
rect 9585 9463 9643 9469
rect 4028 9404 5120 9432
rect 5184 9404 5488 9432
rect 5537 9435 5595 9441
rect 4028 9392 4034 9404
rect 1946 9324 1952 9376
rect 2004 9364 2010 9376
rect 5184 9364 5212 9404
rect 5537 9401 5549 9435
rect 5583 9432 5595 9435
rect 6733 9435 6791 9441
rect 5583 9404 6408 9432
rect 5583 9401 5595 9404
rect 5537 9395 5595 9401
rect 2004 9336 5212 9364
rect 5261 9367 5319 9373
rect 2004 9324 2010 9336
rect 5261 9333 5273 9367
rect 5307 9364 5319 9367
rect 6270 9364 6276 9376
rect 5307 9336 6276 9364
rect 5307 9333 5319 9336
rect 5261 9327 5319 9333
rect 6270 9324 6276 9336
rect 6328 9324 6334 9376
rect 6380 9364 6408 9404
rect 6733 9401 6745 9435
rect 6779 9432 6791 9435
rect 9030 9432 9036 9444
rect 6779 9404 9036 9432
rect 6779 9401 6791 9404
rect 6733 9395 6791 9401
rect 9030 9392 9036 9404
rect 9088 9392 9094 9444
rect 7650 9364 7656 9376
rect 6380 9336 7656 9364
rect 7650 9324 7656 9336
rect 7708 9324 7714 9376
rect 7929 9367 7987 9373
rect 7929 9333 7941 9367
rect 7975 9364 7987 9367
rect 8570 9364 8576 9376
rect 7975 9336 8576 9364
rect 7975 9333 7987 9336
rect 7929 9327 7987 9333
rect 8570 9324 8576 9336
rect 8628 9324 8634 9376
rect 8757 9367 8815 9373
rect 8757 9333 8769 9367
rect 8803 9364 8815 9367
rect 9324 9364 9352 9463
rect 9508 9376 9536 9463
rect 10318 9460 10324 9472
rect 10376 9460 10382 9512
rect 10796 9506 10876 9512
rect 10870 9460 10876 9506
rect 10928 9460 10934 9512
rect 14200 9500 14228 9540
rect 14642 9528 14648 9580
rect 14700 9568 14706 9580
rect 16114 9568 16120 9580
rect 14700 9540 15148 9568
rect 16075 9540 16120 9568
rect 14700 9528 14706 9540
rect 12406 9472 14228 9500
rect 15120 9500 15148 9540
rect 16114 9528 16120 9540
rect 16172 9528 16178 9580
rect 16206 9528 16212 9580
rect 16264 9568 16270 9580
rect 16853 9571 16911 9577
rect 16853 9568 16865 9571
rect 16264 9540 16865 9568
rect 16264 9528 16270 9540
rect 16853 9537 16865 9540
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 17494 9528 17500 9580
rect 17552 9568 17558 9580
rect 17770 9568 17776 9580
rect 17552 9540 17776 9568
rect 17552 9528 17558 9540
rect 17770 9528 17776 9540
rect 17828 9528 17834 9580
rect 17862 9528 17868 9580
rect 17920 9568 17926 9580
rect 18233 9571 18291 9577
rect 18233 9568 18245 9571
rect 17920 9540 18245 9568
rect 17920 9528 17926 9540
rect 18233 9537 18245 9540
rect 18279 9537 18291 9571
rect 18414 9568 18420 9580
rect 18375 9540 18420 9568
rect 18233 9531 18291 9537
rect 18414 9528 18420 9540
rect 18472 9528 18478 9580
rect 19334 9568 19340 9580
rect 18616 9540 19340 9568
rect 17129 9503 17187 9509
rect 17129 9500 17141 9503
rect 15120 9472 17141 9500
rect 9674 9392 9680 9444
rect 9732 9432 9738 9444
rect 12406 9432 12434 9472
rect 17129 9469 17141 9472
rect 17175 9469 17187 9503
rect 18138 9500 18144 9512
rect 17129 9463 17187 9469
rect 17236 9472 18144 9500
rect 9732 9404 12434 9432
rect 13541 9435 13599 9441
rect 9732 9392 9738 9404
rect 13541 9401 13553 9435
rect 13587 9432 13599 9435
rect 13998 9432 14004 9444
rect 13587 9404 14004 9432
rect 13587 9401 13599 9404
rect 13541 9395 13599 9401
rect 13998 9392 14004 9404
rect 14056 9392 14062 9444
rect 15102 9392 15108 9444
rect 15160 9432 15166 9444
rect 15933 9435 15991 9441
rect 15933 9432 15945 9435
rect 15160 9404 15945 9432
rect 15160 9392 15166 9404
rect 15933 9401 15945 9404
rect 15979 9401 15991 9435
rect 17236 9432 17264 9472
rect 18138 9460 18144 9472
rect 18196 9460 18202 9512
rect 18325 9503 18383 9509
rect 18325 9469 18337 9503
rect 18371 9500 18383 9503
rect 18506 9500 18512 9512
rect 18371 9472 18512 9500
rect 18371 9469 18383 9472
rect 18325 9463 18383 9469
rect 18506 9460 18512 9472
rect 18564 9460 18570 9512
rect 15933 9395 15991 9401
rect 16040 9404 17264 9432
rect 8803 9336 9352 9364
rect 8803 9333 8815 9336
rect 8757 9327 8815 9333
rect 9490 9324 9496 9376
rect 9548 9324 9554 9376
rect 10505 9367 10563 9373
rect 10505 9333 10517 9367
rect 10551 9364 10563 9367
rect 10594 9364 10600 9376
rect 10551 9336 10600 9364
rect 10551 9333 10563 9336
rect 10505 9327 10563 9333
rect 10594 9324 10600 9336
rect 10652 9324 10658 9376
rect 10873 9367 10931 9373
rect 10873 9333 10885 9367
rect 10919 9364 10931 9367
rect 11238 9364 11244 9376
rect 10919 9336 11244 9364
rect 10919 9333 10931 9336
rect 10873 9327 10931 9333
rect 11238 9324 11244 9336
rect 11296 9364 11302 9376
rect 11974 9364 11980 9376
rect 11296 9336 11980 9364
rect 11296 9324 11302 9336
rect 11974 9324 11980 9336
rect 12032 9324 12038 9376
rect 13078 9324 13084 9376
rect 13136 9364 13142 9376
rect 15473 9367 15531 9373
rect 15473 9364 15485 9367
rect 13136 9336 15485 9364
rect 13136 9324 13142 9336
rect 15473 9333 15485 9336
rect 15519 9333 15531 9367
rect 15473 9327 15531 9333
rect 15746 9324 15752 9376
rect 15804 9364 15810 9376
rect 16040 9364 16068 9404
rect 17770 9392 17776 9444
rect 17828 9432 17834 9444
rect 18616 9432 18644 9540
rect 19334 9528 19340 9540
rect 19392 9528 19398 9580
rect 20349 9571 20407 9577
rect 20349 9537 20361 9571
rect 20395 9537 20407 9571
rect 20349 9531 20407 9537
rect 18690 9460 18696 9512
rect 18748 9500 18754 9512
rect 18969 9503 19027 9509
rect 18969 9500 18981 9503
rect 18748 9472 18981 9500
rect 18748 9460 18754 9472
rect 18969 9469 18981 9472
rect 19015 9469 19027 9503
rect 18969 9463 19027 9469
rect 19150 9460 19156 9512
rect 19208 9500 19214 9512
rect 20254 9500 20260 9512
rect 19208 9472 20260 9500
rect 19208 9460 19214 9472
rect 20254 9460 20260 9472
rect 20312 9500 20318 9512
rect 20364 9500 20392 9531
rect 20530 9528 20536 9580
rect 20588 9568 20594 9580
rect 20625 9571 20683 9577
rect 20625 9568 20637 9571
rect 20588 9540 20637 9568
rect 20588 9528 20594 9540
rect 20625 9537 20637 9540
rect 20671 9537 20683 9571
rect 20625 9531 20683 9537
rect 20809 9571 20867 9577
rect 20809 9537 20821 9571
rect 20855 9568 20867 9571
rect 21266 9568 21272 9580
rect 20855 9540 21272 9568
rect 20855 9537 20867 9540
rect 20809 9531 20867 9537
rect 21266 9528 21272 9540
rect 21324 9528 21330 9580
rect 21818 9528 21824 9580
rect 21876 9568 21882 9580
rect 22005 9571 22063 9577
rect 22005 9568 22017 9571
rect 21876 9540 22017 9568
rect 21876 9528 21882 9540
rect 22005 9537 22017 9540
rect 22051 9537 22063 9571
rect 22005 9531 22063 9537
rect 22281 9571 22339 9577
rect 22281 9537 22293 9571
rect 22327 9568 22339 9571
rect 22462 9568 22468 9580
rect 22327 9540 22468 9568
rect 22327 9537 22339 9540
rect 22281 9531 22339 9537
rect 22462 9528 22468 9540
rect 22520 9528 22526 9580
rect 22925 9571 22983 9577
rect 22925 9537 22937 9571
rect 22971 9537 22983 9571
rect 22925 9531 22983 9537
rect 23201 9571 23259 9577
rect 23201 9537 23213 9571
rect 23247 9568 23259 9571
rect 23290 9568 23296 9580
rect 23247 9540 23296 9568
rect 23247 9537 23259 9540
rect 23201 9531 23259 9537
rect 22094 9500 22100 9512
rect 20312 9472 22100 9500
rect 20312 9460 20318 9472
rect 22094 9460 22100 9472
rect 22152 9460 22158 9512
rect 22940 9444 22968 9531
rect 23290 9528 23296 9540
rect 23348 9528 23354 9580
rect 24305 9571 24363 9577
rect 24305 9537 24317 9571
rect 24351 9568 24363 9571
rect 25038 9568 25044 9580
rect 24351 9540 25044 9568
rect 24351 9537 24363 9540
rect 24305 9531 24363 9537
rect 25038 9528 25044 9540
rect 25096 9568 25102 9580
rect 25590 9568 25596 9580
rect 25096 9540 25596 9568
rect 25096 9528 25102 9540
rect 25590 9528 25596 9540
rect 25648 9528 25654 9580
rect 25774 9528 25780 9580
rect 25832 9568 25838 9580
rect 27632 9577 27660 9608
rect 29086 9596 29092 9608
rect 29144 9596 29150 9648
rect 27157 9571 27215 9577
rect 27157 9568 27169 9571
rect 25832 9540 27169 9568
rect 25832 9528 25838 9540
rect 27157 9537 27169 9540
rect 27203 9537 27215 9571
rect 27157 9531 27215 9537
rect 27617 9571 27675 9577
rect 27617 9537 27629 9571
rect 27663 9537 27675 9571
rect 27617 9531 27675 9537
rect 27706 9528 27712 9580
rect 27764 9568 27770 9580
rect 27873 9571 27931 9577
rect 27873 9568 27885 9571
rect 27764 9540 27885 9568
rect 27764 9528 27770 9540
rect 27873 9537 27885 9540
rect 27919 9537 27931 9571
rect 27873 9531 27931 9537
rect 29270 9528 29276 9580
rect 29328 9568 29334 9580
rect 29457 9571 29515 9577
rect 29457 9568 29469 9571
rect 29328 9540 29469 9568
rect 29328 9528 29334 9540
rect 29457 9537 29469 9540
rect 29503 9537 29515 9571
rect 29457 9531 29515 9537
rect 30006 9528 30012 9580
rect 30064 9568 30070 9580
rect 31297 9571 31355 9577
rect 31297 9568 31309 9571
rect 30064 9540 31309 9568
rect 30064 9528 30070 9540
rect 31297 9537 31309 9540
rect 31343 9537 31355 9571
rect 31297 9531 31355 9537
rect 24857 9503 24915 9509
rect 24857 9469 24869 9503
rect 24903 9500 24915 9503
rect 24949 9503 25007 9509
rect 24949 9500 24961 9503
rect 24903 9472 24961 9500
rect 24903 9469 24915 9472
rect 24857 9463 24915 9469
rect 24949 9469 24961 9472
rect 24995 9469 25007 9503
rect 24949 9463 25007 9469
rect 29638 9460 29644 9512
rect 29696 9500 29702 9512
rect 29733 9503 29791 9509
rect 29733 9500 29745 9503
rect 29696 9472 29745 9500
rect 29696 9460 29702 9472
rect 29733 9469 29745 9472
rect 29779 9469 29791 9503
rect 29733 9463 29791 9469
rect 17828 9404 18644 9432
rect 17828 9392 17834 9404
rect 19058 9392 19064 9444
rect 19116 9432 19122 9444
rect 19245 9435 19303 9441
rect 19245 9432 19257 9435
rect 19116 9404 19257 9432
rect 19116 9392 19122 9404
rect 19245 9401 19257 9404
rect 19291 9401 19303 9435
rect 19245 9395 19303 9401
rect 19518 9392 19524 9444
rect 19576 9432 19582 9444
rect 20622 9432 20628 9444
rect 19576 9404 20628 9432
rect 19576 9392 19582 9404
rect 20622 9392 20628 9404
rect 20680 9392 20686 9444
rect 21726 9392 21732 9444
rect 21784 9432 21790 9444
rect 21821 9435 21879 9441
rect 21821 9432 21833 9435
rect 21784 9404 21833 9432
rect 21784 9392 21790 9404
rect 21821 9401 21833 9404
rect 21867 9401 21879 9435
rect 21821 9395 21879 9401
rect 22922 9392 22928 9444
rect 22980 9392 22986 9444
rect 23566 9392 23572 9444
rect 23624 9432 23630 9444
rect 24673 9435 24731 9441
rect 24673 9432 24685 9435
rect 23624 9404 24685 9432
rect 23624 9392 23630 9404
rect 24673 9401 24685 9404
rect 24719 9401 24731 9435
rect 24673 9395 24731 9401
rect 25884 9404 27108 9432
rect 15804 9336 16068 9364
rect 15804 9324 15810 9336
rect 16298 9324 16304 9376
rect 16356 9364 16362 9376
rect 16669 9367 16727 9373
rect 16669 9364 16681 9367
rect 16356 9336 16681 9364
rect 16356 9324 16362 9336
rect 16669 9333 16681 9336
rect 16715 9333 16727 9367
rect 17034 9364 17040 9376
rect 16995 9336 17040 9364
rect 16669 9327 16727 9333
rect 17034 9324 17040 9336
rect 17092 9324 17098 9376
rect 17954 9364 17960 9376
rect 17915 9336 17960 9364
rect 17954 9324 17960 9336
rect 18012 9324 18018 9376
rect 18138 9324 18144 9376
rect 18196 9364 18202 9376
rect 19429 9367 19487 9373
rect 19429 9364 19441 9367
rect 18196 9336 19441 9364
rect 18196 9324 18202 9336
rect 19429 9333 19441 9336
rect 19475 9333 19487 9367
rect 19429 9327 19487 9333
rect 19610 9324 19616 9376
rect 19668 9364 19674 9376
rect 20165 9367 20223 9373
rect 20165 9364 20177 9367
rect 19668 9336 20177 9364
rect 19668 9324 19674 9336
rect 20165 9333 20177 9336
rect 20211 9333 20223 9367
rect 20165 9327 20223 9333
rect 22189 9367 22247 9373
rect 22189 9333 22201 9367
rect 22235 9364 22247 9367
rect 23109 9367 23167 9373
rect 23109 9364 23121 9367
rect 22235 9336 23121 9364
rect 22235 9333 22247 9336
rect 22189 9327 22247 9333
rect 23109 9333 23121 9336
rect 23155 9364 23167 9367
rect 23198 9364 23204 9376
rect 23155 9336 23204 9364
rect 23155 9333 23167 9336
rect 23109 9327 23167 9333
rect 23198 9324 23204 9336
rect 23256 9324 23262 9376
rect 23290 9324 23296 9376
rect 23348 9364 23354 9376
rect 23750 9364 23756 9376
rect 23348 9336 23756 9364
rect 23348 9324 23354 9336
rect 23750 9324 23756 9336
rect 23808 9324 23814 9376
rect 24118 9324 24124 9376
rect 24176 9364 24182 9376
rect 25884 9364 25912 9404
rect 24176 9336 25912 9364
rect 24176 9324 24182 9336
rect 25958 9324 25964 9376
rect 26016 9364 26022 9376
rect 26973 9367 27031 9373
rect 26973 9364 26985 9367
rect 26016 9336 26985 9364
rect 26016 9324 26022 9336
rect 26973 9333 26985 9336
rect 27019 9333 27031 9367
rect 27080 9364 27108 9404
rect 28626 9392 28632 9444
rect 28684 9432 28690 9444
rect 30926 9432 30932 9444
rect 28684 9404 30932 9432
rect 28684 9392 28690 9404
rect 30926 9392 30932 9404
rect 30984 9392 30990 9444
rect 28350 9364 28356 9376
rect 27080 9336 28356 9364
rect 26973 9327 27031 9333
rect 28350 9324 28356 9336
rect 28408 9324 28414 9376
rect 28994 9364 29000 9376
rect 28955 9336 29000 9364
rect 28994 9324 29000 9336
rect 29052 9324 29058 9376
rect 31110 9364 31116 9376
rect 31071 9336 31116 9364
rect 31110 9324 31116 9336
rect 31168 9324 31174 9376
rect 1104 9274 32016 9296
rect 1104 9222 2136 9274
rect 2188 9222 12440 9274
rect 12492 9222 22744 9274
rect 22796 9222 32016 9274
rect 1104 9200 32016 9222
rect 3326 9120 3332 9172
rect 3384 9160 3390 9172
rect 3878 9160 3884 9172
rect 3384 9132 3884 9160
rect 3384 9120 3390 9132
rect 3878 9120 3884 9132
rect 3936 9120 3942 9172
rect 4157 9163 4215 9169
rect 4157 9129 4169 9163
rect 4203 9160 4215 9163
rect 4433 9163 4491 9169
rect 4433 9160 4445 9163
rect 4203 9132 4445 9160
rect 4203 9129 4215 9132
rect 4157 9123 4215 9129
rect 4433 9129 4445 9132
rect 4479 9129 4491 9163
rect 4433 9123 4491 9129
rect 5537 9163 5595 9169
rect 5537 9129 5549 9163
rect 5583 9160 5595 9163
rect 7558 9160 7564 9172
rect 5583 9132 7564 9160
rect 5583 9129 5595 9132
rect 5537 9123 5595 9129
rect 7558 9120 7564 9132
rect 7616 9120 7622 9172
rect 8205 9163 8263 9169
rect 8205 9129 8217 9163
rect 8251 9160 8263 9163
rect 8251 9132 13860 9160
rect 8251 9129 8263 9132
rect 8205 9123 8263 9129
rect 2590 9052 2596 9104
rect 2648 9092 2654 9104
rect 9674 9092 9680 9104
rect 2648 9064 9680 9092
rect 2648 9052 2654 9064
rect 9674 9052 9680 9064
rect 9732 9052 9738 9104
rect 11514 9052 11520 9104
rect 11572 9092 11578 9104
rect 11885 9095 11943 9101
rect 11885 9092 11897 9095
rect 11572 9064 11897 9092
rect 11572 9052 11578 9064
rect 11885 9061 11897 9064
rect 11931 9092 11943 9095
rect 12158 9092 12164 9104
rect 11931 9064 12164 9092
rect 11931 9061 11943 9064
rect 11885 9055 11943 9061
rect 12158 9052 12164 9064
rect 12216 9052 12222 9104
rect 12989 9095 13047 9101
rect 12989 9061 13001 9095
rect 13035 9092 13047 9095
rect 13078 9092 13084 9104
rect 13035 9064 13084 9092
rect 13035 9061 13047 9064
rect 12989 9055 13047 9061
rect 13078 9052 13084 9064
rect 13136 9052 13142 9104
rect 13832 9092 13860 9132
rect 13998 9120 14004 9172
rect 14056 9160 14062 9172
rect 17770 9160 17776 9172
rect 14056 9132 17776 9160
rect 14056 9120 14062 9132
rect 17770 9120 17776 9132
rect 17828 9120 17834 9172
rect 17954 9120 17960 9172
rect 18012 9160 18018 9172
rect 24946 9160 24952 9172
rect 18012 9132 24952 9160
rect 18012 9120 18018 9132
rect 24946 9120 24952 9132
rect 25004 9160 25010 9172
rect 25133 9163 25191 9169
rect 25133 9160 25145 9163
rect 25004 9132 25145 9160
rect 25004 9120 25010 9132
rect 25133 9129 25145 9132
rect 25179 9129 25191 9163
rect 26142 9160 26148 9172
rect 26103 9132 26148 9160
rect 25133 9123 25191 9129
rect 26142 9120 26148 9132
rect 26200 9120 26206 9172
rect 27433 9163 27491 9169
rect 27433 9129 27445 9163
rect 27479 9160 27491 9163
rect 27706 9160 27712 9172
rect 27479 9132 27712 9160
rect 27479 9129 27491 9132
rect 27433 9123 27491 9129
rect 27706 9120 27712 9132
rect 27764 9120 27770 9172
rect 27801 9163 27859 9169
rect 27801 9129 27813 9163
rect 27847 9160 27859 9163
rect 28258 9160 28264 9172
rect 27847 9132 28264 9160
rect 27847 9129 27859 9132
rect 27801 9123 27859 9129
rect 28258 9120 28264 9132
rect 28316 9120 28322 9172
rect 28350 9120 28356 9172
rect 28408 9160 28414 9172
rect 30469 9163 30527 9169
rect 30469 9160 30481 9163
rect 28408 9132 30481 9160
rect 28408 9120 28414 9132
rect 30469 9129 30481 9132
rect 30515 9129 30527 9163
rect 30469 9123 30527 9129
rect 14366 9092 14372 9104
rect 13832 9064 14372 9092
rect 14366 9052 14372 9064
rect 14424 9052 14430 9104
rect 17497 9095 17555 9101
rect 17497 9061 17509 9095
rect 17543 9092 17555 9095
rect 18230 9092 18236 9104
rect 17543 9064 18236 9092
rect 17543 9061 17555 9064
rect 17497 9055 17555 9061
rect 18230 9052 18236 9064
rect 18288 9052 18294 9104
rect 18417 9095 18475 9101
rect 18417 9061 18429 9095
rect 18463 9092 18475 9095
rect 19702 9092 19708 9104
rect 18463 9064 19708 9092
rect 18463 9061 18475 9064
rect 18417 9055 18475 9061
rect 2222 8984 2228 9036
rect 2280 9024 2286 9036
rect 2501 9027 2559 9033
rect 2501 9024 2513 9027
rect 2280 8996 2513 9024
rect 2280 8984 2286 8996
rect 2501 8993 2513 8996
rect 2547 8993 2559 9027
rect 2501 8987 2559 8993
rect 2961 9027 3019 9033
rect 2961 8993 2973 9027
rect 3007 9024 3019 9027
rect 5537 9027 5595 9033
rect 5537 9024 5549 9027
rect 3007 8996 5549 9024
rect 3007 8993 3019 8996
rect 2961 8987 3019 8993
rect 5537 8993 5549 8996
rect 5583 8993 5595 9027
rect 5537 8987 5595 8993
rect 5626 8984 5632 9036
rect 5684 9024 5690 9036
rect 6365 9027 6423 9033
rect 6365 9024 6377 9027
rect 5684 8996 6377 9024
rect 5684 8984 5690 8996
rect 6365 8993 6377 8996
rect 6411 8993 6423 9027
rect 6365 8987 6423 8993
rect 8110 8984 8116 9036
rect 8168 9024 8174 9036
rect 10505 9027 10563 9033
rect 10505 9024 10517 9027
rect 8168 8996 10517 9024
rect 8168 8984 8174 8996
rect 10505 8993 10517 8996
rect 10551 8993 10563 9027
rect 10505 8987 10563 8993
rect 12621 9027 12679 9033
rect 12621 8993 12633 9027
rect 12667 9024 12679 9027
rect 12710 9024 12716 9036
rect 12667 8996 12716 9024
rect 12667 8993 12679 8996
rect 12621 8987 12679 8993
rect 12710 8984 12716 8996
rect 12768 9024 12774 9036
rect 13538 9024 13544 9036
rect 12768 8996 13544 9024
rect 12768 8984 12774 8996
rect 13538 8984 13544 8996
rect 13596 8984 13602 9036
rect 14090 8984 14096 9036
rect 14148 9024 14154 9036
rect 14645 9027 14703 9033
rect 14645 9024 14657 9027
rect 14148 8996 14657 9024
rect 14148 8984 14154 8996
rect 14645 8993 14657 8996
rect 14691 8993 14703 9027
rect 14645 8987 14703 8993
rect 15930 8984 15936 9036
rect 15988 9024 15994 9036
rect 16945 9027 17003 9033
rect 16945 9024 16957 9027
rect 15988 8996 16957 9024
rect 15988 8984 15994 8996
rect 16945 8993 16957 8996
rect 16991 8993 17003 9027
rect 18432 9024 18460 9055
rect 19702 9052 19708 9064
rect 19760 9052 19766 9104
rect 21266 9052 21272 9104
rect 21324 9092 21330 9104
rect 21637 9095 21695 9101
rect 21637 9092 21649 9095
rect 21324 9064 21649 9092
rect 21324 9052 21330 9064
rect 21637 9061 21649 9064
rect 21683 9092 21695 9095
rect 21683 9064 22416 9092
rect 21683 9061 21695 9064
rect 21637 9055 21695 9061
rect 19610 9024 19616 9036
rect 16945 8987 17003 8993
rect 17328 8996 18460 9024
rect 19536 8996 19616 9024
rect 1670 8916 1676 8968
rect 1728 8956 1734 8968
rect 2317 8959 2375 8965
rect 2317 8956 2329 8959
rect 1728 8928 2329 8956
rect 1728 8916 1734 8928
rect 2317 8925 2329 8928
rect 2363 8956 2375 8959
rect 2363 8928 3188 8956
rect 2363 8925 2375 8928
rect 2317 8919 2375 8925
rect 2409 8891 2467 8897
rect 2409 8857 2421 8891
rect 2455 8888 2467 8891
rect 2961 8891 3019 8897
rect 2961 8888 2973 8891
rect 2455 8860 2973 8888
rect 2455 8857 2467 8860
rect 2409 8851 2467 8857
rect 2961 8857 2973 8860
rect 3007 8857 3019 8891
rect 3160 8888 3188 8928
rect 3234 8916 3240 8968
rect 3292 8956 3298 8968
rect 3789 8959 3847 8965
rect 3789 8956 3801 8959
rect 3292 8928 3801 8956
rect 3292 8916 3298 8928
rect 3789 8925 3801 8928
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 4890 8916 4896 8968
rect 4948 8956 4954 8968
rect 4985 8959 5043 8965
rect 4985 8956 4997 8959
rect 4948 8928 4997 8956
rect 4948 8916 4954 8928
rect 4985 8925 4997 8928
rect 5031 8925 5043 8959
rect 5258 8956 5264 8968
rect 5219 8928 5264 8956
rect 4985 8919 5043 8925
rect 5258 8916 5264 8928
rect 5316 8916 5322 8968
rect 5442 8956 5448 8968
rect 5403 8928 5448 8956
rect 5442 8916 5448 8928
rect 5500 8916 5506 8968
rect 6089 8959 6147 8965
rect 6089 8956 6101 8959
rect 5552 8928 6101 8956
rect 4062 8888 4068 8900
rect 3160 8860 4068 8888
rect 2961 8851 3019 8857
rect 4062 8848 4068 8860
rect 4120 8848 4126 8900
rect 4801 8891 4859 8897
rect 4801 8857 4813 8891
rect 4847 8888 4859 8891
rect 5552 8888 5580 8928
rect 6089 8925 6101 8928
rect 6135 8925 6147 8959
rect 6089 8919 6147 8925
rect 6270 8916 6276 8968
rect 6328 8956 6334 8968
rect 6914 8956 6920 8968
rect 6328 8928 6421 8956
rect 6875 8928 6920 8956
rect 6328 8916 6334 8928
rect 6914 8916 6920 8928
rect 6972 8916 6978 8968
rect 7098 8916 7104 8968
rect 7156 8956 7162 8968
rect 7193 8959 7251 8965
rect 7193 8956 7205 8959
rect 7156 8928 7205 8956
rect 7156 8916 7162 8928
rect 7193 8925 7205 8928
rect 7239 8925 7251 8959
rect 7193 8919 7251 8925
rect 8389 8959 8447 8965
rect 8389 8925 8401 8959
rect 8435 8956 8447 8959
rect 8757 8959 8815 8965
rect 8757 8956 8769 8959
rect 8435 8928 8769 8956
rect 8435 8925 8447 8928
rect 8389 8919 8447 8925
rect 8757 8925 8769 8928
rect 8803 8925 8815 8959
rect 9214 8956 9220 8968
rect 9175 8928 9220 8956
rect 8757 8919 8815 8925
rect 9214 8916 9220 8928
rect 9272 8916 9278 8968
rect 9309 8959 9367 8965
rect 9309 8925 9321 8959
rect 9355 8925 9367 8959
rect 9309 8919 9367 8925
rect 9493 8959 9551 8965
rect 9493 8925 9505 8959
rect 9539 8925 9551 8959
rect 9493 8919 9551 8925
rect 4847 8860 5580 8888
rect 5905 8891 5963 8897
rect 4847 8857 4859 8860
rect 4801 8851 4859 8857
rect 5905 8857 5917 8891
rect 5951 8888 5963 8891
rect 5994 8888 6000 8900
rect 5951 8860 6000 8888
rect 5951 8857 5963 8860
rect 5905 8851 5963 8857
rect 5994 8848 6000 8860
rect 6052 8848 6058 8900
rect 6288 8888 6316 8916
rect 6638 8888 6644 8900
rect 6288 8860 6644 8888
rect 6638 8848 6644 8860
rect 6696 8888 6702 8900
rect 6696 8860 8156 8888
rect 6696 8848 6702 8860
rect 1946 8820 1952 8832
rect 1907 8792 1952 8820
rect 1946 8780 1952 8792
rect 2004 8780 2010 8832
rect 3050 8780 3056 8832
rect 3108 8820 3114 8832
rect 4157 8823 4215 8829
rect 4157 8820 4169 8823
rect 3108 8792 4169 8820
rect 3108 8780 3114 8792
rect 4157 8789 4169 8792
rect 4203 8789 4215 8823
rect 4338 8820 4344 8832
rect 4299 8792 4344 8820
rect 4157 8783 4215 8789
rect 4338 8780 4344 8792
rect 4396 8780 4402 8832
rect 4433 8823 4491 8829
rect 4433 8789 4445 8823
rect 4479 8820 4491 8823
rect 7466 8820 7472 8832
rect 4479 8792 7472 8820
rect 4479 8789 4491 8792
rect 4433 8783 4491 8789
rect 7466 8780 7472 8792
rect 7524 8820 7530 8832
rect 8018 8820 8024 8832
rect 7524 8792 8024 8820
rect 7524 8780 7530 8792
rect 8018 8780 8024 8792
rect 8076 8780 8082 8832
rect 8128 8820 8156 8860
rect 8294 8848 8300 8900
rect 8352 8888 8358 8900
rect 9324 8888 9352 8919
rect 8352 8860 9352 8888
rect 9508 8888 9536 8919
rect 9582 8916 9588 8968
rect 9640 8956 9646 8968
rect 9953 8959 10011 8965
rect 9953 8956 9965 8959
rect 9640 8928 9965 8956
rect 9640 8916 9646 8928
rect 9953 8925 9965 8928
rect 9999 8925 10011 8959
rect 9953 8919 10011 8925
rect 10594 8916 10600 8968
rect 10652 8956 10658 8968
rect 10761 8959 10819 8965
rect 10761 8956 10773 8959
rect 10652 8928 10773 8956
rect 10652 8916 10658 8928
rect 10761 8925 10773 8928
rect 10807 8925 10819 8959
rect 10761 8919 10819 8925
rect 14912 8959 14970 8965
rect 14912 8925 14924 8959
rect 14958 8956 14970 8959
rect 16298 8956 16304 8968
rect 14958 8928 16304 8956
rect 14958 8925 14970 8928
rect 14912 8919 14970 8925
rect 16298 8916 16304 8928
rect 16356 8916 16362 8968
rect 16574 8916 16580 8968
rect 16632 8956 16638 8968
rect 16669 8959 16727 8965
rect 16669 8956 16681 8959
rect 16632 8928 16681 8956
rect 16632 8916 16638 8928
rect 16669 8925 16681 8928
rect 16715 8925 16727 8959
rect 16669 8919 16727 8925
rect 16853 8959 16911 8965
rect 16853 8925 16865 8959
rect 16899 8956 16911 8959
rect 17034 8956 17040 8968
rect 16899 8928 17040 8956
rect 16899 8925 16911 8928
rect 16853 8919 16911 8925
rect 17034 8916 17040 8928
rect 17092 8956 17098 8968
rect 17328 8956 17356 8996
rect 17092 8928 17356 8956
rect 17405 8959 17463 8965
rect 17092 8916 17098 8928
rect 17405 8925 17417 8959
rect 17451 8956 17463 8959
rect 17494 8956 17500 8968
rect 17451 8928 17500 8956
rect 17451 8925 17463 8928
rect 17405 8919 17463 8925
rect 17494 8916 17500 8928
rect 17552 8916 17558 8968
rect 17589 8959 17647 8965
rect 17589 8925 17601 8959
rect 17635 8956 17647 8959
rect 17862 8956 17868 8968
rect 17635 8928 17868 8956
rect 17635 8925 17647 8928
rect 17589 8919 17647 8925
rect 17862 8916 17868 8928
rect 17920 8916 17926 8968
rect 18230 8956 18236 8968
rect 18191 8928 18236 8956
rect 18230 8916 18236 8928
rect 18288 8916 18294 8968
rect 18506 8916 18512 8968
rect 18564 8956 18570 8968
rect 19536 8965 19564 8996
rect 19610 8984 19616 8996
rect 19668 8984 19674 9036
rect 21542 8984 21548 9036
rect 21600 9024 21606 9036
rect 21818 9024 21824 9036
rect 21600 8996 21824 9024
rect 21600 8984 21606 8996
rect 21818 8984 21824 8996
rect 21876 8984 21882 9036
rect 22388 9024 22416 9064
rect 22462 9052 22468 9104
rect 22520 9092 22526 9104
rect 23109 9095 23167 9101
rect 23109 9092 23121 9095
rect 22520 9064 23121 9092
rect 22520 9052 22526 9064
rect 23109 9061 23121 9064
rect 23155 9061 23167 9095
rect 23109 9055 23167 9061
rect 23198 9052 23204 9104
rect 23256 9092 23262 9104
rect 25866 9092 25872 9104
rect 23256 9064 25872 9092
rect 23256 9052 23262 9064
rect 25866 9052 25872 9064
rect 25924 9092 25930 9104
rect 26513 9095 26571 9101
rect 26513 9092 26525 9095
rect 25924 9064 26525 9092
rect 25924 9052 25930 9064
rect 26513 9061 26525 9064
rect 26559 9061 26571 9095
rect 28074 9092 28080 9104
rect 26513 9055 26571 9061
rect 26620 9064 28080 9092
rect 26620 9033 26648 9064
rect 28074 9052 28080 9064
rect 28132 9052 28138 9104
rect 29270 9052 29276 9104
rect 29328 9092 29334 9104
rect 29328 9064 30052 9092
rect 29328 9052 29334 9064
rect 26605 9027 26663 9033
rect 22388 8996 26096 9024
rect 19521 8959 19579 8965
rect 18564 8928 18609 8956
rect 18564 8916 18570 8928
rect 19521 8925 19533 8959
rect 19567 8925 19579 8959
rect 19702 8956 19708 8968
rect 19663 8928 19708 8956
rect 19521 8919 19579 8925
rect 19702 8916 19708 8928
rect 19760 8916 19766 8968
rect 19797 8959 19855 8965
rect 19797 8925 19809 8959
rect 19843 8956 19855 8959
rect 20073 8959 20131 8965
rect 20073 8956 20085 8959
rect 19843 8928 20085 8956
rect 19843 8925 19855 8928
rect 19797 8919 19855 8925
rect 20073 8925 20085 8928
rect 20119 8925 20131 8959
rect 20073 8919 20131 8925
rect 20162 8916 20168 8968
rect 20220 8956 20226 8968
rect 20257 8959 20315 8965
rect 20257 8956 20269 8959
rect 20220 8928 20269 8956
rect 20220 8916 20226 8928
rect 20257 8925 20269 8928
rect 20303 8925 20315 8959
rect 20257 8919 20315 8925
rect 21082 8916 21088 8968
rect 21140 8956 21146 8968
rect 23109 8959 23167 8965
rect 23109 8956 23121 8959
rect 21140 8928 23121 8956
rect 21140 8916 21146 8928
rect 23109 8925 23121 8928
rect 23155 8925 23167 8959
rect 23109 8919 23167 8925
rect 23198 8916 23204 8968
rect 23256 8956 23262 8968
rect 23385 8959 23443 8965
rect 23385 8956 23397 8959
rect 23256 8928 23397 8956
rect 23256 8916 23262 8928
rect 23385 8925 23397 8928
rect 23431 8925 23443 8959
rect 23385 8919 23443 8925
rect 11698 8888 11704 8900
rect 9508 8860 11704 8888
rect 8352 8848 8358 8860
rect 11698 8848 11704 8860
rect 11756 8848 11762 8900
rect 18138 8888 18144 8900
rect 11808 8860 12434 8888
rect 8478 8820 8484 8832
rect 8128 8792 8484 8820
rect 8478 8780 8484 8792
rect 8536 8780 8542 8832
rect 8757 8823 8815 8829
rect 8757 8789 8769 8823
rect 8803 8820 8815 8823
rect 11808 8820 11836 8860
rect 8803 8792 11836 8820
rect 12406 8820 12434 8860
rect 13004 8860 18144 8888
rect 13004 8820 13032 8860
rect 18138 8848 18144 8860
rect 18196 8848 18202 8900
rect 19337 8891 19395 8897
rect 19337 8857 19349 8891
rect 19383 8888 19395 8891
rect 20502 8891 20560 8897
rect 20502 8888 20514 8891
rect 19383 8860 20514 8888
rect 19383 8857 19395 8860
rect 19337 8851 19395 8857
rect 20502 8857 20514 8860
rect 20548 8857 20560 8891
rect 22278 8888 22284 8900
rect 22239 8860 22284 8888
rect 20502 8851 20560 8857
rect 22278 8848 22284 8860
rect 22336 8848 22342 8900
rect 22646 8888 22652 8900
rect 22559 8860 22652 8888
rect 22646 8848 22652 8860
rect 22704 8888 22710 8900
rect 22833 8891 22891 8897
rect 22833 8888 22845 8891
rect 22704 8860 22845 8888
rect 22704 8848 22710 8860
rect 22833 8857 22845 8860
rect 22879 8857 22891 8891
rect 22833 8851 22891 8857
rect 24854 8848 24860 8900
rect 24912 8888 24918 8900
rect 24949 8891 25007 8897
rect 24949 8888 24961 8891
rect 24912 8860 24961 8888
rect 24912 8848 24918 8860
rect 24949 8857 24961 8860
rect 24995 8857 25007 8891
rect 26068 8888 26096 8996
rect 26605 8993 26617 9027
rect 26651 8993 26663 9027
rect 28353 9027 28411 9033
rect 28353 9024 28365 9027
rect 26605 8987 26663 8993
rect 27632 8996 28365 9024
rect 26326 8956 26332 8968
rect 26287 8928 26332 8956
rect 26326 8916 26332 8928
rect 26384 8916 26390 8968
rect 27632 8965 27660 8996
rect 28353 8993 28365 8996
rect 28399 8993 28411 9027
rect 29638 9024 29644 9036
rect 28353 8987 28411 8993
rect 28828 8996 29644 9024
rect 27617 8959 27675 8965
rect 27617 8925 27629 8959
rect 27663 8925 27675 8959
rect 27617 8919 27675 8925
rect 27893 8959 27951 8965
rect 27893 8925 27905 8959
rect 27939 8925 27951 8959
rect 28534 8956 28540 8968
rect 28495 8928 28540 8956
rect 27893 8919 27951 8925
rect 27908 8888 27936 8919
rect 28534 8916 28540 8928
rect 28592 8916 28598 8968
rect 28828 8965 28856 8996
rect 29638 8984 29644 8996
rect 29696 8984 29702 9036
rect 30024 9033 30052 9064
rect 30009 9027 30067 9033
rect 30009 8993 30021 9027
rect 30055 8993 30067 9027
rect 30009 8987 30067 8993
rect 28813 8959 28871 8965
rect 28813 8925 28825 8959
rect 28859 8925 28871 8959
rect 28813 8919 28871 8925
rect 28994 8916 29000 8968
rect 29052 8956 29058 8968
rect 29733 8959 29791 8965
rect 29052 8928 29145 8956
rect 29052 8916 29058 8928
rect 29733 8925 29745 8959
rect 29779 8925 29791 8959
rect 29733 8919 29791 8925
rect 29917 8959 29975 8965
rect 29917 8925 29929 8959
rect 29963 8956 29975 8959
rect 30653 8959 30711 8965
rect 29963 8928 30512 8956
rect 29963 8925 29975 8928
rect 29917 8919 29975 8925
rect 26068 8860 27936 8888
rect 24949 8851 25007 8857
rect 12406 8792 13032 8820
rect 13081 8823 13139 8829
rect 8803 8789 8815 8792
rect 8757 8783 8815 8789
rect 13081 8789 13093 8823
rect 13127 8820 13139 8823
rect 13630 8820 13636 8832
rect 13127 8792 13636 8820
rect 13127 8789 13139 8792
rect 13081 8783 13139 8789
rect 13630 8780 13636 8792
rect 13688 8780 13694 8832
rect 13906 8780 13912 8832
rect 13964 8820 13970 8832
rect 15746 8820 15752 8832
rect 13964 8792 15752 8820
rect 13964 8780 13970 8792
rect 15746 8780 15752 8792
rect 15804 8780 15810 8832
rect 15930 8780 15936 8832
rect 15988 8820 15994 8832
rect 16025 8823 16083 8829
rect 16025 8820 16037 8823
rect 15988 8792 16037 8820
rect 15988 8780 15994 8792
rect 16025 8789 16037 8792
rect 16071 8789 16083 8823
rect 16482 8820 16488 8832
rect 16443 8792 16488 8820
rect 16025 8783 16083 8789
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 18049 8823 18107 8829
rect 18049 8789 18061 8823
rect 18095 8820 18107 8823
rect 18322 8820 18328 8832
rect 18095 8792 18328 8820
rect 18095 8789 18107 8792
rect 18049 8783 18107 8789
rect 18322 8780 18328 8792
rect 18380 8780 18386 8832
rect 19426 8780 19432 8832
rect 19484 8820 19490 8832
rect 19978 8820 19984 8832
rect 19484 8792 19984 8820
rect 19484 8780 19490 8792
rect 19978 8780 19984 8792
rect 20036 8780 20042 8832
rect 20073 8823 20131 8829
rect 20073 8789 20085 8823
rect 20119 8820 20131 8823
rect 20714 8820 20720 8832
rect 20119 8792 20720 8820
rect 20119 8789 20131 8792
rect 20073 8783 20131 8789
rect 20714 8780 20720 8792
rect 20772 8780 20778 8832
rect 23014 8780 23020 8832
rect 23072 8820 23078 8832
rect 23293 8823 23351 8829
rect 23072 8792 23117 8820
rect 23072 8780 23078 8792
rect 23293 8789 23305 8823
rect 23339 8820 23351 8823
rect 23750 8820 23756 8832
rect 23339 8792 23756 8820
rect 23339 8789 23351 8792
rect 23293 8783 23351 8789
rect 23750 8780 23756 8792
rect 23808 8780 23814 8832
rect 25038 8780 25044 8832
rect 25096 8820 25102 8832
rect 25149 8823 25207 8829
rect 25149 8820 25161 8823
rect 25096 8792 25161 8820
rect 25096 8780 25102 8792
rect 25149 8789 25161 8792
rect 25195 8789 25207 8823
rect 25149 8783 25207 8789
rect 25317 8823 25375 8829
rect 25317 8789 25329 8823
rect 25363 8820 25375 8823
rect 25958 8820 25964 8832
rect 25363 8792 25964 8820
rect 25363 8789 25375 8792
rect 25317 8783 25375 8789
rect 25958 8780 25964 8792
rect 26016 8780 26022 8832
rect 27338 8780 27344 8832
rect 27396 8820 27402 8832
rect 29012 8820 29040 8916
rect 29748 8888 29776 8919
rect 30374 8888 30380 8900
rect 29748 8860 30380 8888
rect 30374 8848 30380 8860
rect 30432 8848 30438 8900
rect 30484 8888 30512 8928
rect 30653 8925 30665 8959
rect 30699 8956 30711 8959
rect 30926 8956 30932 8968
rect 30699 8928 30932 8956
rect 30699 8925 30711 8928
rect 30653 8919 30711 8925
rect 30926 8916 30932 8928
rect 30984 8916 30990 8968
rect 31294 8956 31300 8968
rect 31255 8928 31300 8956
rect 31294 8916 31300 8928
rect 31352 8916 31358 8968
rect 31386 8888 31392 8900
rect 30484 8860 31392 8888
rect 31386 8848 31392 8860
rect 31444 8848 31450 8900
rect 27396 8792 29040 8820
rect 29549 8823 29607 8829
rect 27396 8780 27402 8792
rect 29549 8789 29561 8823
rect 29595 8820 29607 8823
rect 29822 8820 29828 8832
rect 29595 8792 29828 8820
rect 29595 8789 29607 8792
rect 29549 8783 29607 8789
rect 29822 8780 29828 8792
rect 29880 8780 29886 8832
rect 30650 8780 30656 8832
rect 30708 8820 30714 8832
rect 31113 8823 31171 8829
rect 31113 8820 31125 8823
rect 30708 8792 31125 8820
rect 30708 8780 30714 8792
rect 31113 8789 31125 8792
rect 31159 8789 31171 8823
rect 31113 8783 31171 8789
rect 1104 8730 32016 8752
rect 1104 8678 7288 8730
rect 7340 8678 17592 8730
rect 17644 8678 27896 8730
rect 27948 8678 32016 8730
rect 1104 8656 32016 8678
rect 4338 8616 4344 8628
rect 1872 8588 4344 8616
rect 1872 8557 1900 8588
rect 4338 8576 4344 8588
rect 4396 8576 4402 8628
rect 5534 8616 5540 8628
rect 5495 8588 5540 8616
rect 5534 8576 5540 8588
rect 5592 8576 5598 8628
rect 5644 8588 6684 8616
rect 1857 8551 1915 8557
rect 1857 8517 1869 8551
rect 1903 8517 1915 8551
rect 1857 8511 1915 8517
rect 1946 8508 1952 8560
rect 2004 8548 2010 8560
rect 3053 8551 3111 8557
rect 2004 8520 2176 8548
rect 2004 8508 2010 8520
rect 1762 8440 1768 8492
rect 1820 8480 1826 8492
rect 2148 8489 2176 8520
rect 3053 8517 3065 8551
rect 3099 8548 3111 8551
rect 3421 8551 3479 8557
rect 3421 8548 3433 8551
rect 3099 8520 3433 8548
rect 3099 8517 3111 8520
rect 3053 8511 3111 8517
rect 3421 8517 3433 8520
rect 3467 8517 3479 8551
rect 3421 8511 3479 8517
rect 3602 8508 3608 8560
rect 3660 8548 3666 8560
rect 5644 8548 5672 8588
rect 3660 8520 5672 8548
rect 6656 8548 6684 8588
rect 6914 8576 6920 8628
rect 6972 8616 6978 8628
rect 7745 8619 7803 8625
rect 7745 8616 7757 8619
rect 6972 8588 7757 8616
rect 6972 8576 6978 8588
rect 7745 8585 7757 8588
rect 7791 8585 7803 8619
rect 7745 8579 7803 8585
rect 8205 8619 8263 8625
rect 8205 8585 8217 8619
rect 8251 8616 8263 8619
rect 8294 8616 8300 8628
rect 8251 8588 8300 8616
rect 8251 8585 8263 8588
rect 8205 8579 8263 8585
rect 8294 8576 8300 8588
rect 8352 8576 8358 8628
rect 8570 8616 8576 8628
rect 8531 8588 8576 8616
rect 8570 8576 8576 8588
rect 8628 8576 8634 8628
rect 8662 8576 8668 8628
rect 8720 8616 8726 8628
rect 19288 8616 19294 8628
rect 8720 8588 19294 8616
rect 8720 8576 8726 8588
rect 19288 8576 19294 8588
rect 19346 8576 19352 8628
rect 19978 8576 19984 8628
rect 20036 8616 20042 8628
rect 31110 8616 31116 8628
rect 20036 8588 31116 8616
rect 20036 8576 20042 8588
rect 31110 8576 31116 8588
rect 31168 8576 31174 8628
rect 9674 8548 9680 8560
rect 6656 8520 6776 8548
rect 3660 8508 3666 8520
rect 2041 8483 2099 8489
rect 2041 8480 2053 8483
rect 1820 8452 2053 8480
rect 1820 8440 1826 8452
rect 2041 8449 2053 8452
rect 2087 8449 2099 8483
rect 2041 8443 2099 8449
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8449 2191 8483
rect 2133 8443 2191 8449
rect 2961 8483 3019 8489
rect 2961 8449 2973 8483
rect 3007 8480 3019 8483
rect 3326 8480 3332 8492
rect 3007 8452 3332 8480
rect 3007 8449 3019 8452
rect 2961 8443 3019 8449
rect 3326 8440 3332 8452
rect 3384 8480 3390 8492
rect 3970 8480 3976 8492
rect 3384 8452 3976 8480
rect 3384 8440 3390 8452
rect 3970 8440 3976 8452
rect 4028 8440 4034 8492
rect 4154 8480 4160 8492
rect 4115 8452 4160 8480
rect 4154 8440 4160 8452
rect 4212 8440 4218 8492
rect 4424 8483 4482 8489
rect 4424 8449 4436 8483
rect 4470 8470 4482 8483
rect 6270 8480 6276 8492
rect 4520 8470 6276 8480
rect 4470 8452 6276 8470
rect 4470 8449 4548 8452
rect 4424 8443 4548 8449
rect 4439 8442 4548 8443
rect 6270 8440 6276 8452
rect 6328 8440 6334 8492
rect 6454 8440 6460 8492
rect 6512 8480 6518 8492
rect 6621 8483 6679 8489
rect 6621 8480 6633 8483
rect 6512 8452 6633 8480
rect 6512 8440 6518 8452
rect 6621 8449 6633 8452
rect 6667 8449 6679 8483
rect 6748 8480 6776 8520
rect 8220 8520 9680 8548
rect 8220 8480 8248 8520
rect 9674 8508 9680 8520
rect 9732 8508 9738 8560
rect 9769 8551 9827 8557
rect 9769 8517 9781 8551
rect 9815 8548 9827 8551
rect 9858 8548 9864 8560
rect 9815 8520 9864 8548
rect 9815 8517 9827 8520
rect 9769 8511 9827 8517
rect 9858 8508 9864 8520
rect 9916 8508 9922 8560
rect 9968 8520 10732 8548
rect 6748 8452 8248 8480
rect 6621 8443 6679 8449
rect 8938 8440 8944 8492
rect 8996 8480 9002 8492
rect 9968 8480 9996 8520
rect 10594 8480 10600 8492
rect 8996 8452 9996 8480
rect 10555 8452 10600 8480
rect 8996 8440 9002 8452
rect 10594 8440 10600 8452
rect 10652 8440 10658 8492
rect 10704 8480 10732 8520
rect 10778 8508 10784 8560
rect 10836 8548 10842 8560
rect 11609 8551 11667 8557
rect 11609 8548 11621 8551
rect 10836 8520 11621 8548
rect 10836 8508 10842 8520
rect 11609 8517 11621 8520
rect 11655 8517 11667 8551
rect 14090 8548 14096 8560
rect 11609 8511 11667 8517
rect 13004 8520 14096 8548
rect 13004 8489 13032 8520
rect 14090 8508 14096 8520
rect 14148 8508 14154 8560
rect 16482 8508 16488 8560
rect 16540 8548 16546 8560
rect 16914 8551 16972 8557
rect 16914 8548 16926 8551
rect 16540 8520 16926 8548
rect 16540 8508 16546 8520
rect 16914 8517 16926 8520
rect 16960 8517 16972 8551
rect 16914 8511 16972 8517
rect 17034 8508 17040 8560
rect 17092 8508 17098 8560
rect 17494 8508 17500 8560
rect 17552 8548 17558 8560
rect 18690 8548 18696 8560
rect 17552 8520 18696 8548
rect 17552 8508 17558 8520
rect 18690 8508 18696 8520
rect 18748 8508 18754 8560
rect 18874 8508 18880 8560
rect 18932 8548 18938 8560
rect 21821 8551 21879 8557
rect 21821 8548 21833 8551
rect 18932 8520 21833 8548
rect 18932 8508 18938 8520
rect 21821 8517 21833 8520
rect 21867 8517 21879 8551
rect 21821 8511 21879 8517
rect 22554 8508 22560 8560
rect 22612 8548 22618 8560
rect 22612 8520 22784 8548
rect 22612 8508 22618 8520
rect 12345 8483 12403 8489
rect 12345 8480 12357 8483
rect 10704 8452 12357 8480
rect 12345 8449 12357 8452
rect 12391 8449 12403 8483
rect 12345 8443 12403 8449
rect 12989 8483 13047 8489
rect 12989 8449 13001 8483
rect 13035 8449 13047 8483
rect 12989 8443 13047 8449
rect 13256 8483 13314 8489
rect 13256 8449 13268 8483
rect 13302 8480 13314 8483
rect 15654 8480 15660 8492
rect 13302 8452 15660 8480
rect 13302 8449 13314 8452
rect 13256 8443 13314 8449
rect 15654 8440 15660 8452
rect 15712 8440 15718 8492
rect 17052 8480 17080 8508
rect 16500 8452 17080 8480
rect 2314 8372 2320 8424
rect 2372 8412 2378 8424
rect 3234 8412 3240 8424
rect 2372 8384 2774 8412
rect 3195 8384 3240 8412
rect 2372 8372 2378 8384
rect 1857 8347 1915 8353
rect 1857 8313 1869 8347
rect 1903 8344 1915 8347
rect 2406 8344 2412 8356
rect 1903 8316 2412 8344
rect 1903 8313 1915 8316
rect 1857 8307 1915 8313
rect 2406 8304 2412 8316
rect 2464 8304 2470 8356
rect 2746 8344 2774 8384
rect 3234 8372 3240 8384
rect 3292 8372 3298 8424
rect 5994 8372 6000 8424
rect 6052 8412 6058 8424
rect 6365 8415 6423 8421
rect 6365 8412 6377 8415
rect 6052 8384 6377 8412
rect 6052 8372 6058 8384
rect 6365 8381 6377 8384
rect 6411 8381 6423 8415
rect 6365 8375 6423 8381
rect 8202 8372 8208 8424
rect 8260 8412 8266 8424
rect 8665 8415 8723 8421
rect 8665 8412 8677 8415
rect 8260 8384 8677 8412
rect 8260 8372 8266 8384
rect 8665 8381 8677 8384
rect 8711 8381 8723 8415
rect 8665 8375 8723 8381
rect 8849 8415 8907 8421
rect 8849 8381 8861 8415
rect 8895 8412 8907 8415
rect 9401 8415 9459 8421
rect 9401 8412 9413 8415
rect 8895 8384 9413 8412
rect 8895 8381 8907 8384
rect 8849 8375 8907 8381
rect 9401 8381 9413 8384
rect 9447 8412 9459 8415
rect 10873 8415 10931 8421
rect 10873 8412 10885 8415
rect 9447 8384 10885 8412
rect 9447 8381 9459 8384
rect 9401 8375 9459 8381
rect 10873 8381 10885 8384
rect 10919 8412 10931 8415
rect 10962 8412 10968 8424
rect 10919 8384 10968 8412
rect 10919 8381 10931 8384
rect 10873 8375 10931 8381
rect 10962 8372 10968 8384
rect 11020 8372 11026 8424
rect 11238 8412 11244 8424
rect 11072 8384 11244 8412
rect 3252 8344 3280 8372
rect 2746 8316 3280 8344
rect 3421 8347 3479 8353
rect 3421 8313 3433 8347
rect 3467 8344 3479 8347
rect 3970 8344 3976 8356
rect 3467 8316 3976 8344
rect 3467 8313 3479 8316
rect 3421 8307 3479 8313
rect 3970 8304 3976 8316
rect 4028 8304 4034 8356
rect 7650 8304 7656 8356
rect 7708 8344 7714 8356
rect 9306 8344 9312 8356
rect 7708 8316 9312 8344
rect 7708 8304 7714 8316
rect 9306 8304 9312 8316
rect 9364 8304 9370 8356
rect 9953 8347 10011 8353
rect 9953 8344 9965 8347
rect 9416 8316 9965 8344
rect 2590 8276 2596 8288
rect 2551 8248 2596 8276
rect 2590 8236 2596 8248
rect 2648 8236 2654 8288
rect 2682 8236 2688 8288
rect 2740 8276 2746 8288
rect 4890 8276 4896 8288
rect 2740 8248 4896 8276
rect 2740 8236 2746 8248
rect 4890 8236 4896 8248
rect 4948 8236 4954 8288
rect 5074 8236 5080 8288
rect 5132 8276 5138 8288
rect 6638 8276 6644 8288
rect 5132 8248 6644 8276
rect 5132 8236 5138 8248
rect 6638 8236 6644 8248
rect 6696 8236 6702 8288
rect 9122 8236 9128 8288
rect 9180 8276 9186 8288
rect 9416 8276 9444 8316
rect 9953 8313 9965 8316
rect 9999 8313 10011 8347
rect 9953 8307 10011 8313
rect 10413 8347 10471 8353
rect 10413 8313 10425 8347
rect 10459 8344 10471 8347
rect 10502 8344 10508 8356
rect 10459 8316 10508 8344
rect 10459 8313 10471 8316
rect 10413 8307 10471 8313
rect 10502 8304 10508 8316
rect 10560 8304 10566 8356
rect 10781 8347 10839 8353
rect 10781 8313 10793 8347
rect 10827 8344 10839 8347
rect 11072 8344 11100 8384
rect 11238 8372 11244 8384
rect 11296 8412 11302 8424
rect 12529 8415 12587 8421
rect 12529 8412 12541 8415
rect 11296 8384 12541 8412
rect 11296 8372 11302 8384
rect 12529 8381 12541 8384
rect 12575 8381 12587 8415
rect 15289 8415 15347 8421
rect 12529 8375 12587 8381
rect 14200 8384 15240 8412
rect 11793 8347 11851 8353
rect 11793 8344 11805 8347
rect 10827 8316 11100 8344
rect 11164 8316 11805 8344
rect 10827 8313 10839 8316
rect 10781 8307 10839 8313
rect 9766 8276 9772 8288
rect 9180 8248 9444 8276
rect 9727 8248 9772 8276
rect 9180 8236 9186 8248
rect 9766 8236 9772 8248
rect 9824 8236 9830 8288
rect 10134 8236 10140 8288
rect 10192 8276 10198 8288
rect 11164 8276 11192 8316
rect 11793 8313 11805 8316
rect 11839 8313 11851 8347
rect 14200 8344 14228 8384
rect 14366 8344 14372 8356
rect 11793 8307 11851 8313
rect 13924 8316 14228 8344
rect 14279 8316 14372 8344
rect 10192 8248 11192 8276
rect 10192 8236 10198 8248
rect 13354 8236 13360 8288
rect 13412 8276 13418 8288
rect 13924 8276 13952 8316
rect 14366 8304 14372 8316
rect 14424 8344 14430 8356
rect 14642 8344 14648 8356
rect 14424 8316 14648 8344
rect 14424 8304 14430 8316
rect 14642 8304 14648 8316
rect 14700 8304 14706 8356
rect 15212 8344 15240 8384
rect 15289 8381 15301 8415
rect 15335 8412 15347 8415
rect 15378 8412 15384 8424
rect 15335 8384 15384 8412
rect 15335 8381 15347 8384
rect 15289 8375 15347 8381
rect 15378 8372 15384 8384
rect 15436 8372 15442 8424
rect 15565 8415 15623 8421
rect 15565 8381 15577 8415
rect 15611 8412 15623 8415
rect 16500 8412 16528 8452
rect 18230 8440 18236 8492
rect 18288 8480 18294 8492
rect 18969 8483 19027 8489
rect 18969 8480 18981 8483
rect 18288 8452 18981 8480
rect 18288 8440 18294 8452
rect 18969 8449 18981 8452
rect 19015 8449 19027 8483
rect 18969 8443 19027 8449
rect 19150 8440 19156 8492
rect 19208 8480 19214 8492
rect 19429 8483 19487 8489
rect 19208 8452 19253 8480
rect 19208 8440 19214 8452
rect 19429 8449 19441 8483
rect 19475 8480 19487 8483
rect 19625 8483 19683 8489
rect 19475 8452 19555 8480
rect 19475 8449 19487 8452
rect 19429 8443 19487 8449
rect 16666 8412 16672 8424
rect 15611 8384 16528 8412
rect 16627 8384 16672 8412
rect 15611 8381 15623 8384
rect 15565 8375 15623 8381
rect 16666 8372 16672 8384
rect 16724 8372 16730 8424
rect 19527 8412 19555 8452
rect 19625 8449 19637 8483
rect 19671 8480 19683 8483
rect 19794 8480 19800 8492
rect 19671 8452 19800 8480
rect 19671 8449 19683 8452
rect 19625 8443 19683 8449
rect 19794 8440 19800 8452
rect 19852 8440 19858 8492
rect 20254 8480 20260 8492
rect 20215 8452 20260 8480
rect 20254 8440 20260 8452
rect 20312 8440 20318 8492
rect 20530 8480 20536 8492
rect 20443 8452 20536 8480
rect 20530 8440 20536 8452
rect 20588 8440 20594 8492
rect 20714 8480 20720 8492
rect 20675 8452 20720 8480
rect 20714 8440 20720 8452
rect 20772 8440 20778 8492
rect 21726 8440 21732 8492
rect 21784 8480 21790 8492
rect 22649 8483 22707 8489
rect 22649 8480 22661 8483
rect 21784 8452 22661 8480
rect 21784 8440 21790 8452
rect 22649 8449 22661 8452
rect 22695 8449 22707 8483
rect 22756 8480 22784 8520
rect 23014 8508 23020 8560
rect 23072 8548 23078 8560
rect 23937 8551 23995 8557
rect 23937 8548 23949 8551
rect 23072 8520 23949 8548
rect 23072 8508 23078 8520
rect 23937 8517 23949 8520
rect 23983 8517 23995 8551
rect 23937 8511 23995 8517
rect 24153 8551 24211 8557
rect 24153 8517 24165 8551
rect 24199 8548 24211 8551
rect 25038 8548 25044 8560
rect 24199 8520 25044 8548
rect 24199 8517 24211 8520
rect 24153 8511 24211 8517
rect 25038 8508 25044 8520
rect 25096 8508 25102 8560
rect 25130 8508 25136 8560
rect 25188 8548 25194 8560
rect 25188 8520 25452 8548
rect 25188 8508 25194 8520
rect 23106 8480 23112 8492
rect 22756 8452 23112 8480
rect 22649 8443 22707 8449
rect 23106 8440 23112 8452
rect 23164 8440 23170 8492
rect 23198 8440 23204 8492
rect 23256 8480 23262 8492
rect 23293 8483 23351 8489
rect 23293 8480 23305 8483
rect 23256 8452 23305 8480
rect 23256 8440 23262 8452
rect 23293 8449 23305 8452
rect 23339 8449 23351 8483
rect 23293 8443 23351 8449
rect 24394 8440 24400 8492
rect 24452 8480 24458 8492
rect 24857 8483 24915 8489
rect 24857 8480 24869 8483
rect 24452 8452 24869 8480
rect 24452 8440 24458 8452
rect 24857 8449 24869 8452
rect 24903 8449 24915 8483
rect 25222 8480 25228 8492
rect 25183 8452 25228 8480
rect 24857 8443 24915 8449
rect 25222 8440 25228 8452
rect 25280 8440 25286 8492
rect 25424 8489 25452 8520
rect 26050 8508 26056 8560
rect 26108 8548 26114 8560
rect 27798 8548 27804 8560
rect 26108 8520 27804 8548
rect 26108 8508 26114 8520
rect 27798 8508 27804 8520
rect 27856 8548 27862 8560
rect 28629 8551 28687 8557
rect 28629 8548 28641 8551
rect 27856 8520 28641 8548
rect 27856 8508 27862 8520
rect 28629 8517 28641 8520
rect 28675 8517 28687 8551
rect 28629 8511 28687 8517
rect 25409 8483 25467 8489
rect 25409 8449 25421 8483
rect 25455 8449 25467 8483
rect 25409 8443 25467 8449
rect 25685 8483 25743 8489
rect 25685 8449 25697 8483
rect 25731 8480 25743 8483
rect 26145 8483 26203 8489
rect 26145 8480 26157 8483
rect 25731 8452 26157 8480
rect 25731 8449 25743 8452
rect 25685 8443 25743 8449
rect 26145 8449 26157 8452
rect 26191 8449 26203 8483
rect 26145 8443 26203 8449
rect 27065 8483 27123 8489
rect 27065 8449 27077 8483
rect 27111 8480 27123 8483
rect 27614 8480 27620 8492
rect 27111 8452 27620 8480
rect 27111 8449 27123 8452
rect 27065 8443 27123 8449
rect 27614 8440 27620 8452
rect 27672 8440 27678 8492
rect 27893 8483 27951 8489
rect 27893 8449 27905 8483
rect 27939 8480 27951 8483
rect 29730 8480 29736 8492
rect 27939 8452 29736 8480
rect 27939 8449 27951 8452
rect 27893 8443 27951 8449
rect 29730 8440 29736 8452
rect 29788 8440 29794 8492
rect 31018 8480 31024 8492
rect 30979 8452 31024 8480
rect 31018 8440 31024 8452
rect 31076 8440 31082 8492
rect 19444 8384 19555 8412
rect 15212 8316 16574 8344
rect 13412 8248 13952 8276
rect 16546 8276 16574 8316
rect 17954 8304 17960 8356
rect 18012 8344 18018 8356
rect 18049 8347 18107 8353
rect 18049 8344 18061 8347
rect 18012 8316 18061 8344
rect 18012 8304 18018 8316
rect 18049 8313 18061 8316
rect 18095 8344 18107 8347
rect 18506 8344 18512 8356
rect 18095 8316 18512 8344
rect 18095 8313 18107 8316
rect 18049 8307 18107 8313
rect 18506 8304 18512 8316
rect 18564 8304 18570 8356
rect 19444 8276 19472 8384
rect 19610 8304 19616 8356
rect 19668 8344 19674 8356
rect 20073 8347 20131 8353
rect 20073 8344 20085 8347
rect 19668 8316 20085 8344
rect 19668 8304 19674 8316
rect 20073 8313 20085 8316
rect 20119 8313 20131 8347
rect 20073 8307 20131 8313
rect 20548 8276 20576 8440
rect 22373 8415 22431 8421
rect 22373 8381 22385 8415
rect 22419 8412 22431 8415
rect 22554 8412 22560 8424
rect 22419 8384 22560 8412
rect 22419 8381 22431 8384
rect 22373 8375 22431 8381
rect 22554 8372 22560 8384
rect 22612 8372 22618 8424
rect 22830 8372 22836 8424
rect 22888 8412 22894 8424
rect 25774 8412 25780 8424
rect 22888 8384 22933 8412
rect 23032 8384 25780 8412
rect 22888 8372 22894 8384
rect 20622 8304 20628 8356
rect 20680 8344 20686 8356
rect 23032 8344 23060 8384
rect 25774 8372 25780 8384
rect 25832 8372 25838 8424
rect 27338 8372 27344 8424
rect 27396 8412 27402 8424
rect 28169 8415 28227 8421
rect 28169 8412 28181 8415
rect 27396 8384 28181 8412
rect 27396 8372 27402 8384
rect 28169 8381 28181 8384
rect 28215 8381 28227 8415
rect 31294 8412 31300 8424
rect 28169 8375 28227 8381
rect 28276 8384 30972 8412
rect 31255 8384 31300 8412
rect 28276 8356 28304 8384
rect 20680 8316 23060 8344
rect 23385 8347 23443 8353
rect 20680 8304 20686 8316
rect 23385 8313 23397 8347
rect 23431 8344 23443 8347
rect 23750 8344 23756 8356
rect 23431 8316 23756 8344
rect 23431 8313 23443 8316
rect 23385 8307 23443 8313
rect 23750 8304 23756 8316
rect 23808 8304 23814 8356
rect 24305 8347 24363 8353
rect 24305 8313 24317 8347
rect 24351 8344 24363 8347
rect 24578 8344 24584 8356
rect 24351 8316 24584 8344
rect 24351 8313 24363 8316
rect 24305 8307 24363 8313
rect 24578 8304 24584 8316
rect 24636 8304 24642 8356
rect 24857 8347 24915 8353
rect 24857 8313 24869 8347
rect 24903 8344 24915 8347
rect 25685 8347 25743 8353
rect 25685 8344 25697 8347
rect 24903 8316 25697 8344
rect 24903 8313 24915 8316
rect 24857 8307 24915 8313
rect 25685 8313 25697 8316
rect 25731 8313 25743 8347
rect 25685 8307 25743 8313
rect 26329 8347 26387 8353
rect 26329 8313 26341 8347
rect 26375 8344 26387 8347
rect 26602 8344 26608 8356
rect 26375 8316 26608 8344
rect 26375 8313 26387 8316
rect 26329 8307 26387 8313
rect 26602 8304 26608 8316
rect 26660 8344 26666 8356
rect 27522 8344 27528 8356
rect 26660 8316 27528 8344
rect 26660 8304 26666 8316
rect 27522 8304 27528 8316
rect 27580 8304 27586 8356
rect 28077 8347 28135 8353
rect 28077 8313 28089 8347
rect 28123 8344 28135 8347
rect 28258 8344 28264 8356
rect 28123 8316 28264 8344
rect 28123 8313 28135 8316
rect 28077 8307 28135 8313
rect 28258 8304 28264 8316
rect 28316 8304 28322 8356
rect 30190 8304 30196 8356
rect 30248 8344 30254 8356
rect 30837 8347 30895 8353
rect 30837 8344 30849 8347
rect 30248 8316 30849 8344
rect 30248 8304 30254 8316
rect 30837 8313 30849 8316
rect 30883 8313 30895 8347
rect 30944 8344 30972 8384
rect 31294 8372 31300 8384
rect 31352 8372 31358 8424
rect 31205 8347 31263 8353
rect 31205 8344 31217 8347
rect 30944 8316 31217 8344
rect 30837 8307 30895 8313
rect 31205 8313 31217 8316
rect 31251 8344 31263 8347
rect 31386 8344 31392 8356
rect 31251 8316 31392 8344
rect 31251 8313 31263 8316
rect 31205 8307 31263 8313
rect 31386 8304 31392 8316
rect 31444 8304 31450 8356
rect 16546 8248 20576 8276
rect 13412 8236 13418 8248
rect 22278 8236 22284 8288
rect 22336 8276 22342 8288
rect 23290 8276 23296 8288
rect 22336 8248 23296 8276
rect 22336 8236 22342 8248
rect 23290 8236 23296 8248
rect 23348 8236 23354 8288
rect 24121 8279 24179 8285
rect 24121 8245 24133 8279
rect 24167 8276 24179 8279
rect 24486 8276 24492 8288
rect 24167 8248 24492 8276
rect 24167 8245 24179 8248
rect 24121 8239 24179 8245
rect 24486 8236 24492 8248
rect 24544 8236 24550 8288
rect 25590 8276 25596 8288
rect 25551 8248 25596 8276
rect 25590 8236 25596 8248
rect 25648 8236 25654 8288
rect 27157 8279 27215 8285
rect 27157 8245 27169 8279
rect 27203 8276 27215 8279
rect 27246 8276 27252 8288
rect 27203 8248 27252 8276
rect 27203 8245 27215 8248
rect 27157 8239 27215 8245
rect 27246 8236 27252 8248
rect 27304 8236 27310 8288
rect 27709 8279 27767 8285
rect 27709 8245 27721 8279
rect 27755 8276 27767 8279
rect 27982 8276 27988 8288
rect 27755 8248 27988 8276
rect 27755 8245 27767 8248
rect 27709 8239 27767 8245
rect 27982 8236 27988 8248
rect 28040 8236 28046 8288
rect 29086 8236 29092 8288
rect 29144 8276 29150 8288
rect 29638 8276 29644 8288
rect 29144 8248 29644 8276
rect 29144 8236 29150 8248
rect 29638 8236 29644 8248
rect 29696 8276 29702 8288
rect 29917 8279 29975 8285
rect 29917 8276 29929 8279
rect 29696 8248 29929 8276
rect 29696 8236 29702 8248
rect 29917 8245 29929 8248
rect 29963 8245 29975 8279
rect 29917 8239 29975 8245
rect 1104 8186 32016 8208
rect 0 8140 800 8154
rect 0 8112 1072 8140
rect 1104 8134 2136 8186
rect 2188 8134 12440 8186
rect 12492 8134 22744 8186
rect 22796 8134 32016 8186
rect 1104 8112 32016 8134
rect 32125 8143 32183 8149
rect 0 8098 800 8112
rect 1044 8072 1072 8112
rect 32125 8109 32137 8143
rect 32171 8140 32183 8143
rect 32320 8140 33120 8154
rect 32171 8112 33120 8140
rect 32171 8109 32183 8112
rect 32125 8103 32183 8109
rect 32320 8098 33120 8112
rect 2682 8072 2688 8084
rect 1044 8044 2688 8072
rect 2682 8032 2688 8044
rect 2740 8032 2746 8084
rect 3789 8075 3847 8081
rect 3789 8041 3801 8075
rect 3835 8072 3847 8075
rect 6454 8072 6460 8084
rect 3835 8044 6460 8072
rect 3835 8041 3847 8044
rect 3789 8035 3847 8041
rect 6454 8032 6460 8044
rect 6512 8032 6518 8084
rect 8202 8072 8208 8084
rect 8163 8044 8208 8072
rect 8202 8032 8208 8044
rect 8260 8032 8266 8084
rect 8941 8075 8999 8081
rect 8941 8041 8953 8075
rect 8987 8072 8999 8075
rect 9214 8072 9220 8084
rect 8987 8044 9220 8072
rect 8987 8041 8999 8044
rect 8941 8035 8999 8041
rect 9214 8032 9220 8044
rect 9272 8032 9278 8084
rect 10594 8032 10600 8084
rect 10652 8072 10658 8084
rect 11149 8075 11207 8081
rect 11149 8072 11161 8075
rect 10652 8044 11161 8072
rect 10652 8032 10658 8044
rect 11149 8041 11161 8044
rect 11195 8041 11207 8075
rect 13446 8072 13452 8084
rect 13407 8044 13452 8072
rect 11149 8035 11207 8041
rect 13446 8032 13452 8044
rect 13504 8032 13510 8084
rect 15381 8075 15439 8081
rect 15381 8041 15393 8075
rect 15427 8072 15439 8075
rect 16206 8072 16212 8084
rect 15427 8044 16212 8072
rect 15427 8041 15439 8044
rect 15381 8035 15439 8041
rect 16206 8032 16212 8044
rect 16264 8032 16270 8084
rect 16850 8032 16856 8084
rect 16908 8072 16914 8084
rect 17218 8072 17224 8084
rect 16908 8044 17224 8072
rect 16908 8032 16914 8044
rect 17218 8032 17224 8044
rect 17276 8032 17282 8084
rect 18417 8075 18475 8081
rect 18417 8041 18429 8075
rect 18463 8072 18475 8075
rect 18782 8072 18788 8084
rect 18463 8044 18788 8072
rect 18463 8041 18475 8044
rect 18417 8035 18475 8041
rect 18782 8032 18788 8044
rect 18840 8032 18846 8084
rect 20714 8072 20720 8084
rect 20675 8044 20720 8072
rect 20714 8032 20720 8044
rect 20772 8072 20778 8084
rect 21634 8072 21640 8084
rect 20772 8044 21640 8072
rect 20772 8032 20778 8044
rect 21634 8032 21640 8044
rect 21692 8032 21698 8084
rect 21726 8032 21732 8084
rect 21784 8072 21790 8084
rect 21821 8075 21879 8081
rect 21821 8072 21833 8075
rect 21784 8044 21833 8072
rect 21784 8032 21790 8044
rect 21821 8041 21833 8044
rect 21867 8041 21879 8075
rect 21821 8035 21879 8041
rect 22370 8032 22376 8084
rect 22428 8072 22434 8084
rect 27065 8075 27123 8081
rect 22428 8044 24808 8072
rect 22428 8032 22434 8044
rect 6178 8004 6184 8016
rect 4264 7976 6184 8004
rect 1394 7896 1400 7948
rect 1452 7936 1458 7948
rect 2406 7936 2412 7948
rect 1452 7908 2412 7936
rect 1452 7896 1458 7908
rect 2406 7896 2412 7908
rect 2464 7936 2470 7948
rect 3050 7936 3056 7948
rect 2464 7908 3056 7936
rect 2464 7896 2470 7908
rect 1581 7871 1639 7877
rect 1581 7837 1593 7871
rect 1627 7868 1639 7871
rect 1762 7868 1768 7880
rect 1627 7840 1768 7868
rect 1627 7837 1639 7840
rect 1581 7831 1639 7837
rect 1762 7828 1768 7840
rect 1820 7828 1826 7880
rect 2222 7868 2228 7880
rect 2183 7840 2228 7868
rect 2222 7828 2228 7840
rect 2280 7828 2286 7880
rect 2498 7868 2504 7880
rect 2459 7840 2504 7868
rect 2498 7828 2504 7840
rect 2556 7828 2562 7880
rect 2700 7877 2728 7908
rect 3050 7896 3056 7908
rect 3108 7896 3114 7948
rect 4264 7945 4292 7976
rect 6178 7964 6184 7976
rect 6236 7964 6242 8016
rect 8018 8004 8024 8016
rect 7979 7976 8024 8004
rect 8018 7964 8024 7976
rect 8076 7964 8082 8016
rect 9953 8007 10011 8013
rect 9953 7973 9965 8007
rect 9999 8004 10011 8007
rect 10226 8004 10232 8016
rect 9999 7976 10232 8004
rect 9999 7973 10011 7976
rect 9953 7967 10011 7973
rect 10226 7964 10232 7976
rect 10284 8004 10290 8016
rect 11057 8007 11115 8013
rect 11057 8004 11069 8007
rect 10284 7976 11069 8004
rect 10284 7964 10290 7976
rect 11057 7973 11069 7976
rect 11103 8004 11115 8007
rect 11606 8004 11612 8016
rect 11103 7976 11612 8004
rect 11103 7973 11115 7976
rect 11057 7967 11115 7973
rect 11606 7964 11612 7976
rect 11664 7964 11670 8016
rect 12618 7964 12624 8016
rect 12676 8004 12682 8016
rect 12713 8007 12771 8013
rect 12713 8004 12725 8007
rect 12676 7976 12725 8004
rect 12676 7964 12682 7976
rect 12713 7973 12725 7976
rect 12759 8004 12771 8007
rect 16022 8004 16028 8016
rect 12759 7976 16028 8004
rect 12759 7973 12771 7976
rect 12713 7967 12771 7973
rect 16022 7964 16028 7976
rect 16080 7964 16086 8016
rect 4249 7939 4307 7945
rect 4249 7905 4261 7939
rect 4295 7905 4307 7939
rect 5074 7936 5080 7948
rect 4249 7899 4307 7905
rect 4724 7908 5080 7936
rect 2685 7871 2743 7877
rect 2685 7837 2697 7871
rect 2731 7837 2743 7871
rect 2685 7831 2743 7837
rect 3973 7871 4031 7877
rect 3973 7837 3985 7871
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 4157 7871 4215 7877
rect 4157 7837 4169 7871
rect 4203 7868 4215 7871
rect 4724 7868 4752 7908
rect 5074 7896 5080 7908
rect 5132 7896 5138 7948
rect 5258 7936 5264 7948
rect 5171 7908 5264 7936
rect 4203 7840 4752 7868
rect 4203 7837 4215 7840
rect 4157 7831 4215 7837
rect 3602 7800 3608 7812
rect 1412 7772 3608 7800
rect 1412 7741 1440 7772
rect 3602 7760 3608 7772
rect 3660 7760 3666 7812
rect 3988 7800 4016 7831
rect 4798 7828 4804 7880
rect 4856 7868 4862 7880
rect 5184 7877 5212 7908
rect 5258 7896 5264 7908
rect 5316 7936 5322 7948
rect 5442 7936 5448 7948
rect 5316 7908 5448 7936
rect 5316 7896 5322 7908
rect 5442 7896 5448 7908
rect 5500 7936 5506 7948
rect 5500 7908 6500 7936
rect 5500 7896 5506 7908
rect 4893 7871 4951 7877
rect 4893 7868 4905 7871
rect 4856 7840 4905 7868
rect 4856 7828 4862 7840
rect 4893 7837 4905 7840
rect 4939 7837 4951 7871
rect 4893 7831 4951 7837
rect 5169 7871 5227 7877
rect 5169 7837 5181 7871
rect 5215 7837 5227 7871
rect 5169 7831 5227 7837
rect 5353 7871 5411 7877
rect 5353 7837 5365 7871
rect 5399 7868 5411 7871
rect 5534 7868 5540 7880
rect 5399 7840 5540 7868
rect 5399 7837 5411 7840
rect 5353 7831 5411 7837
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 6472 7877 6500 7908
rect 6730 7896 6736 7948
rect 6788 7936 6794 7948
rect 6788 7908 7328 7936
rect 6788 7896 6794 7908
rect 6181 7871 6239 7877
rect 6181 7837 6193 7871
rect 6227 7837 6239 7871
rect 6181 7831 6239 7837
rect 6457 7871 6515 7877
rect 6457 7837 6469 7871
rect 6503 7837 6515 7871
rect 6457 7831 6515 7837
rect 6641 7871 6699 7877
rect 6641 7837 6653 7871
rect 6687 7868 6699 7871
rect 7098 7868 7104 7880
rect 6687 7840 7104 7868
rect 6687 7837 6699 7840
rect 6641 7831 6699 7837
rect 5997 7803 6055 7809
rect 5997 7800 6009 7803
rect 3988 7772 6009 7800
rect 5997 7769 6009 7772
rect 6043 7769 6055 7803
rect 6196 7800 6224 7831
rect 7098 7828 7104 7840
rect 7156 7828 7162 7880
rect 7300 7877 7328 7908
rect 7374 7896 7380 7948
rect 7432 7936 7438 7948
rect 7745 7939 7803 7945
rect 7745 7936 7757 7939
rect 7432 7908 7757 7936
rect 7432 7896 7438 7908
rect 7745 7905 7757 7908
rect 7791 7936 7803 7939
rect 9766 7936 9772 7948
rect 7791 7908 9772 7936
rect 7791 7905 7803 7908
rect 7745 7899 7803 7905
rect 9766 7896 9772 7908
rect 9824 7896 9830 7948
rect 16298 7936 16304 7948
rect 9876 7908 11652 7936
rect 7285 7871 7343 7877
rect 7285 7837 7297 7871
rect 7331 7837 7343 7871
rect 9122 7868 9128 7880
rect 9083 7840 9128 7868
rect 7285 7831 7343 7837
rect 9122 7828 9128 7840
rect 9180 7828 9186 7880
rect 9401 7871 9459 7877
rect 9401 7868 9413 7871
rect 9223 7840 9413 7868
rect 6914 7800 6920 7812
rect 6196 7772 6920 7800
rect 5997 7763 6055 7769
rect 6914 7760 6920 7772
rect 6972 7760 6978 7812
rect 9030 7760 9036 7812
rect 9088 7800 9094 7812
rect 9223 7800 9251 7840
rect 9401 7837 9413 7840
rect 9447 7837 9459 7871
rect 9401 7831 9459 7837
rect 9674 7828 9680 7880
rect 9732 7868 9738 7880
rect 9876 7868 9904 7908
rect 9732 7840 9904 7868
rect 9953 7871 10011 7877
rect 9732 7828 9738 7840
rect 9953 7837 9965 7871
rect 9999 7868 10011 7871
rect 10229 7871 10287 7877
rect 10229 7868 10241 7871
rect 9999 7840 10241 7868
rect 9999 7837 10011 7840
rect 9953 7831 10011 7837
rect 10229 7837 10241 7840
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 10410 7828 10416 7880
rect 10468 7868 10474 7880
rect 10520 7877 10548 7908
rect 10505 7871 10563 7877
rect 10505 7868 10517 7871
rect 10468 7840 10517 7868
rect 10468 7828 10474 7840
rect 10505 7837 10517 7840
rect 10551 7837 10563 7871
rect 10505 7831 10563 7837
rect 10689 7871 10747 7877
rect 10689 7837 10701 7871
rect 10735 7868 10747 7871
rect 10962 7868 10968 7880
rect 10735 7840 10968 7868
rect 10735 7837 10747 7840
rect 10689 7831 10747 7837
rect 9088 7772 9251 7800
rect 9309 7803 9367 7809
rect 9088 7760 9094 7772
rect 9309 7769 9321 7803
rect 9355 7800 9367 7803
rect 10704 7800 10732 7831
rect 10962 7828 10968 7840
rect 11020 7828 11026 7880
rect 11624 7877 11652 7908
rect 11891 7908 16304 7936
rect 11057 7871 11115 7877
rect 11057 7837 11069 7871
rect 11103 7868 11115 7871
rect 11333 7871 11391 7877
rect 11333 7868 11345 7871
rect 11103 7840 11345 7868
rect 11103 7837 11115 7840
rect 11057 7831 11115 7837
rect 11333 7837 11345 7840
rect 11379 7837 11391 7871
rect 11333 7831 11391 7837
rect 11609 7871 11667 7877
rect 11609 7837 11621 7871
rect 11655 7837 11667 7871
rect 11609 7831 11667 7837
rect 11698 7828 11704 7880
rect 11756 7868 11762 7880
rect 11793 7871 11851 7877
rect 11793 7868 11805 7871
rect 11756 7840 11805 7868
rect 11756 7828 11762 7840
rect 11793 7837 11805 7840
rect 11839 7837 11851 7871
rect 11793 7831 11851 7837
rect 9355 7772 10732 7800
rect 9355 7769 9367 7772
rect 9309 7763 9367 7769
rect 10778 7760 10784 7812
rect 10836 7800 10842 7812
rect 11891 7800 11919 7908
rect 16298 7896 16304 7908
rect 16356 7896 16362 7948
rect 21910 7896 21916 7948
rect 21968 7936 21974 7948
rect 24780 7945 24808 8044
rect 27065 8041 27077 8075
rect 27111 8072 27123 8075
rect 29270 8072 29276 8084
rect 27111 8044 29276 8072
rect 27111 8041 27123 8044
rect 27065 8035 27123 8041
rect 29270 8032 29276 8044
rect 29328 8032 29334 8084
rect 30929 8075 30987 8081
rect 30929 8072 30941 8075
rect 29564 8044 30941 8072
rect 26513 8007 26571 8013
rect 26513 7973 26525 8007
rect 26559 7973 26571 8007
rect 26513 7967 26571 7973
rect 24765 7939 24823 7945
rect 21968 7908 22508 7936
rect 21968 7896 21974 7908
rect 12526 7868 12532 7880
rect 12487 7840 12532 7868
rect 12526 7828 12532 7840
rect 12584 7828 12590 7880
rect 12802 7868 12808 7880
rect 12763 7840 12808 7868
rect 12802 7828 12808 7840
rect 12860 7828 12866 7880
rect 13357 7871 13415 7877
rect 13357 7837 13369 7871
rect 13403 7868 13415 7871
rect 14090 7868 14096 7880
rect 13403 7840 14096 7868
rect 13403 7837 13415 7840
rect 13357 7831 13415 7837
rect 14090 7828 14096 7840
rect 14148 7868 14154 7880
rect 14274 7868 14280 7880
rect 14148 7840 14280 7868
rect 14148 7828 14154 7840
rect 14274 7828 14280 7840
rect 14332 7828 14338 7880
rect 14369 7871 14427 7877
rect 14369 7837 14381 7871
rect 14415 7837 14427 7871
rect 14369 7831 14427 7837
rect 10836 7772 11919 7800
rect 14384 7800 14412 7831
rect 14734 7828 14740 7880
rect 14792 7868 14798 7880
rect 15102 7868 15108 7880
rect 14792 7840 15108 7868
rect 14792 7828 14798 7840
rect 15102 7828 15108 7840
rect 15160 7868 15166 7880
rect 15565 7871 15623 7877
rect 15565 7868 15577 7871
rect 15160 7840 15577 7868
rect 15160 7828 15166 7840
rect 15565 7837 15577 7840
rect 15611 7837 15623 7871
rect 15565 7831 15623 7837
rect 15841 7871 15899 7877
rect 15841 7837 15853 7871
rect 15887 7837 15899 7871
rect 15841 7831 15899 7837
rect 15010 7800 15016 7812
rect 14384 7772 15016 7800
rect 10836 7760 10842 7772
rect 15010 7760 15016 7772
rect 15068 7800 15074 7812
rect 15856 7800 15884 7831
rect 15930 7828 15936 7880
rect 15988 7868 15994 7880
rect 16025 7871 16083 7877
rect 16025 7868 16037 7871
rect 15988 7840 16037 7868
rect 15988 7828 15994 7840
rect 16025 7837 16037 7840
rect 16071 7837 16083 7871
rect 16025 7831 16083 7837
rect 16666 7828 16672 7880
rect 16724 7868 16730 7880
rect 17037 7871 17095 7877
rect 17037 7868 17049 7871
rect 16724 7840 17049 7868
rect 16724 7828 16730 7840
rect 17037 7837 17049 7840
rect 17083 7868 17095 7871
rect 17678 7868 17684 7880
rect 17083 7840 17684 7868
rect 17083 7837 17095 7840
rect 17037 7831 17095 7837
rect 17678 7828 17684 7840
rect 17736 7868 17742 7880
rect 19337 7871 19395 7877
rect 19337 7868 19349 7871
rect 17736 7840 19349 7868
rect 17736 7828 17742 7840
rect 19337 7837 19349 7840
rect 19383 7868 19395 7871
rect 20162 7868 20168 7880
rect 19383 7840 20168 7868
rect 19383 7837 19395 7840
rect 19337 7831 19395 7837
rect 20162 7828 20168 7840
rect 20220 7828 20226 7880
rect 21266 7868 21272 7880
rect 21227 7840 21272 7868
rect 21266 7828 21272 7840
rect 21324 7828 21330 7880
rect 22002 7828 22008 7880
rect 22060 7868 22066 7880
rect 22094 7868 22100 7880
rect 22060 7840 22100 7868
rect 22060 7828 22066 7840
rect 22094 7828 22100 7840
rect 22152 7868 22158 7880
rect 22373 7871 22431 7877
rect 22373 7868 22385 7871
rect 22152 7840 22385 7868
rect 22152 7828 22158 7840
rect 22373 7837 22385 7840
rect 22419 7837 22431 7871
rect 22480 7868 22508 7908
rect 24765 7905 24777 7939
rect 24811 7905 24823 7939
rect 24765 7899 24823 7905
rect 25133 7939 25191 7945
rect 25133 7905 25145 7939
rect 25179 7936 25191 7939
rect 26528 7936 26556 7967
rect 26970 7936 26976 7948
rect 25179 7908 26976 7936
rect 25179 7905 25191 7908
rect 25133 7899 25191 7905
rect 24118 7868 24124 7880
rect 22480 7840 24124 7868
rect 22373 7831 22431 7837
rect 24118 7828 24124 7840
rect 24176 7828 24182 7880
rect 24946 7868 24952 7880
rect 24907 7840 24952 7868
rect 24946 7828 24952 7840
rect 25004 7828 25010 7880
rect 25590 7868 25596 7880
rect 25503 7840 25596 7868
rect 25590 7828 25596 7840
rect 25648 7828 25654 7880
rect 25792 7877 25820 7908
rect 26970 7896 26976 7908
rect 27028 7936 27034 7948
rect 27801 7939 27859 7945
rect 27801 7936 27813 7939
rect 27028 7908 27813 7936
rect 27028 7896 27034 7908
rect 27801 7905 27813 7908
rect 27847 7905 27859 7939
rect 27801 7899 27859 7905
rect 28215 7939 28273 7945
rect 28215 7905 28227 7939
rect 28261 7936 28273 7939
rect 29564 7936 29592 8044
rect 30929 8041 30941 8044
rect 30975 8072 30987 8075
rect 31294 8072 31300 8084
rect 30975 8044 31300 8072
rect 30975 8041 30987 8044
rect 30929 8035 30987 8041
rect 31294 8032 31300 8044
rect 31352 8032 31358 8084
rect 28261 7908 29592 7936
rect 28261 7905 28273 7908
rect 28215 7899 28273 7905
rect 25777 7871 25835 7877
rect 25777 7837 25789 7871
rect 25823 7837 25835 7871
rect 25777 7831 25835 7837
rect 27065 7871 27123 7877
rect 27065 7837 27077 7871
rect 27111 7868 27123 7871
rect 27157 7871 27215 7877
rect 27157 7868 27169 7871
rect 27111 7840 27169 7868
rect 27111 7837 27123 7840
rect 27065 7831 27123 7837
rect 27157 7837 27169 7840
rect 27203 7837 27215 7871
rect 27338 7868 27344 7880
rect 27299 7840 27344 7868
rect 27157 7831 27215 7837
rect 27338 7828 27344 7840
rect 27396 7828 27402 7880
rect 28074 7828 28080 7880
rect 28132 7868 28138 7880
rect 28350 7868 28356 7880
rect 28132 7840 28177 7868
rect 28311 7840 28356 7868
rect 28132 7828 28138 7840
rect 28350 7828 28356 7840
rect 28408 7828 28414 7880
rect 29549 7871 29607 7877
rect 29549 7837 29561 7871
rect 29595 7868 29607 7871
rect 29638 7868 29644 7880
rect 29595 7840 29644 7868
rect 29595 7837 29607 7840
rect 29549 7831 29607 7837
rect 29638 7828 29644 7840
rect 29696 7828 29702 7880
rect 29822 7877 29828 7880
rect 29816 7868 29828 7877
rect 29783 7840 29828 7868
rect 29816 7831 29828 7840
rect 29822 7828 29828 7831
rect 29880 7828 29886 7880
rect 16942 7800 16948 7812
rect 15068 7772 16948 7800
rect 15068 7760 15074 7772
rect 16942 7760 16948 7772
rect 17000 7760 17006 7812
rect 17304 7803 17362 7809
rect 17304 7769 17316 7803
rect 17350 7800 17362 7803
rect 17494 7800 17500 7812
rect 17350 7772 17500 7800
rect 17350 7769 17362 7772
rect 17304 7763 17362 7769
rect 17494 7760 17500 7772
rect 17552 7760 17558 7812
rect 19426 7760 19432 7812
rect 19484 7800 19490 7812
rect 19582 7803 19640 7809
rect 19582 7800 19594 7803
rect 19484 7772 19594 7800
rect 19484 7760 19490 7772
rect 19582 7769 19594 7772
rect 19628 7769 19640 7803
rect 19582 7763 19640 7769
rect 21818 7760 21824 7812
rect 21876 7800 21882 7812
rect 22618 7803 22676 7809
rect 22618 7800 22630 7803
rect 21876 7772 22630 7800
rect 21876 7760 21882 7772
rect 22618 7769 22630 7772
rect 22664 7769 22676 7803
rect 25608 7800 25636 7828
rect 26142 7800 26148 7812
rect 25608 7772 26148 7800
rect 22618 7763 22676 7769
rect 26142 7760 26148 7772
rect 26200 7800 26206 7812
rect 26237 7803 26295 7809
rect 26237 7800 26249 7803
rect 26200 7772 26249 7800
rect 26200 7760 26206 7772
rect 26237 7769 26249 7772
rect 26283 7769 26295 7803
rect 26237 7763 26295 7769
rect 28828 7772 29776 7800
rect 1397 7735 1455 7741
rect 1397 7701 1409 7735
rect 1443 7701 1455 7735
rect 1397 7695 1455 7701
rect 1946 7692 1952 7744
rect 2004 7732 2010 7744
rect 2041 7735 2099 7741
rect 2041 7732 2053 7735
rect 2004 7704 2053 7732
rect 2004 7692 2010 7704
rect 2041 7701 2053 7704
rect 2087 7701 2099 7735
rect 2041 7695 2099 7701
rect 4709 7735 4767 7741
rect 4709 7701 4721 7735
rect 4755 7732 4767 7735
rect 6546 7732 6552 7744
rect 4755 7704 6552 7732
rect 4755 7701 4767 7704
rect 4709 7695 4767 7701
rect 6546 7692 6552 7704
rect 6604 7692 6610 7744
rect 7101 7735 7159 7741
rect 7101 7701 7113 7735
rect 7147 7732 7159 7735
rect 9953 7735 10011 7741
rect 9953 7732 9965 7735
rect 7147 7704 9965 7732
rect 7147 7701 7159 7704
rect 7101 7695 7159 7701
rect 9953 7701 9965 7704
rect 9999 7701 10011 7735
rect 9953 7695 10011 7701
rect 10045 7735 10103 7741
rect 10045 7701 10057 7735
rect 10091 7732 10103 7735
rect 10410 7732 10416 7744
rect 10091 7704 10416 7732
rect 10091 7701 10103 7704
rect 10045 7695 10103 7701
rect 10410 7692 10416 7704
rect 10468 7692 10474 7744
rect 12342 7732 12348 7744
rect 12303 7704 12348 7732
rect 12342 7692 12348 7704
rect 12400 7692 12406 7744
rect 13538 7692 13544 7744
rect 13596 7732 13602 7744
rect 16850 7732 16856 7744
rect 13596 7704 16856 7732
rect 13596 7692 13602 7704
rect 16850 7692 16856 7704
rect 16908 7692 16914 7744
rect 21082 7692 21088 7744
rect 21140 7732 21146 7744
rect 21646 7735 21704 7741
rect 21646 7732 21658 7735
rect 21140 7704 21658 7732
rect 21140 7692 21146 7704
rect 21646 7701 21658 7704
rect 21692 7701 21704 7735
rect 21646 7695 21704 7701
rect 23658 7692 23664 7744
rect 23716 7732 23722 7744
rect 23753 7735 23811 7741
rect 23753 7732 23765 7735
rect 23716 7704 23765 7732
rect 23716 7692 23722 7704
rect 23753 7701 23765 7704
rect 23799 7701 23811 7735
rect 23753 7695 23811 7701
rect 25685 7735 25743 7741
rect 25685 7701 25697 7735
rect 25731 7732 25743 7735
rect 25774 7732 25780 7744
rect 25731 7704 25780 7732
rect 25731 7701 25743 7704
rect 25685 7695 25743 7701
rect 25774 7692 25780 7704
rect 25832 7692 25838 7744
rect 26694 7732 26700 7744
rect 26655 7704 26700 7732
rect 26694 7692 26700 7704
rect 26752 7692 26758 7744
rect 28074 7692 28080 7744
rect 28132 7732 28138 7744
rect 28828 7732 28856 7772
rect 28994 7732 29000 7744
rect 28132 7704 28856 7732
rect 28955 7704 29000 7732
rect 28132 7692 28138 7704
rect 28994 7692 29000 7704
rect 29052 7692 29058 7744
rect 29748 7732 29776 7772
rect 31202 7732 31208 7744
rect 29748 7704 31208 7732
rect 31202 7692 31208 7704
rect 31260 7692 31266 7744
rect 1104 7642 32016 7664
rect 1104 7590 7288 7642
rect 7340 7590 17592 7642
rect 17644 7590 27896 7642
rect 27948 7590 32016 7642
rect 1104 7568 32016 7590
rect 2038 7528 2044 7540
rect 1999 7500 2044 7528
rect 2038 7488 2044 7500
rect 2096 7488 2102 7540
rect 3970 7488 3976 7540
rect 4028 7528 4034 7540
rect 5258 7528 5264 7540
rect 4028 7500 5264 7528
rect 4028 7488 4034 7500
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 5350 7488 5356 7540
rect 5408 7488 5414 7540
rect 5626 7488 5632 7540
rect 5684 7528 5690 7540
rect 5994 7528 6000 7540
rect 5684 7500 6000 7528
rect 5684 7488 5690 7500
rect 5994 7488 6000 7500
rect 6052 7528 6058 7540
rect 6181 7531 6239 7537
rect 6181 7528 6193 7531
rect 6052 7500 6193 7528
rect 6052 7488 6058 7500
rect 6181 7497 6193 7500
rect 6227 7497 6239 7531
rect 6181 7491 6239 7497
rect 6270 7488 6276 7540
rect 6328 7528 6334 7540
rect 6365 7531 6423 7537
rect 6365 7528 6377 7531
rect 6328 7500 6377 7528
rect 6328 7488 6334 7500
rect 6365 7497 6377 7500
rect 6411 7497 6423 7531
rect 8754 7528 8760 7540
rect 8715 7500 8760 7528
rect 6365 7491 6423 7497
rect 8754 7488 8760 7500
rect 8812 7488 8818 7540
rect 10042 7488 10048 7540
rect 10100 7528 10106 7540
rect 10778 7528 10784 7540
rect 10100 7500 10784 7528
rect 10100 7488 10106 7500
rect 10778 7488 10784 7500
rect 10836 7488 10842 7540
rect 10962 7528 10968 7540
rect 10923 7500 10968 7528
rect 10962 7488 10968 7500
rect 11020 7488 11026 7540
rect 12526 7488 12532 7540
rect 12584 7528 12590 7540
rect 14553 7531 14611 7537
rect 14553 7528 14565 7531
rect 12584 7500 14565 7528
rect 12584 7488 12590 7500
rect 14553 7497 14565 7500
rect 14599 7497 14611 7531
rect 15654 7528 15660 7540
rect 15615 7500 15660 7528
rect 14553 7491 14611 7497
rect 15654 7488 15660 7500
rect 15712 7488 15718 7540
rect 16574 7488 16580 7540
rect 16632 7528 16638 7540
rect 16669 7531 16727 7537
rect 16669 7528 16681 7531
rect 16632 7500 16681 7528
rect 16632 7488 16638 7500
rect 16669 7497 16681 7500
rect 16715 7497 16727 7531
rect 16669 7491 16727 7497
rect 21085 7531 21143 7537
rect 21085 7497 21097 7531
rect 21131 7528 21143 7531
rect 21818 7528 21824 7540
rect 21131 7500 21824 7528
rect 21131 7497 21143 7500
rect 21085 7491 21143 7497
rect 21818 7488 21824 7500
rect 21876 7488 21882 7540
rect 22189 7531 22247 7537
rect 22189 7528 22201 7531
rect 21928 7500 22201 7528
rect 4798 7460 4804 7472
rect 2516 7432 3372 7460
rect 2516 7404 2544 7432
rect 1581 7395 1639 7401
rect 1581 7361 1593 7395
rect 1627 7392 1639 7395
rect 1762 7392 1768 7404
rect 1627 7364 1768 7392
rect 1627 7361 1639 7364
rect 1581 7355 1639 7361
rect 1762 7352 1768 7364
rect 1820 7392 1826 7404
rect 2222 7392 2228 7404
rect 1820 7364 2084 7392
rect 2183 7364 2228 7392
rect 1820 7352 1826 7364
rect 2056 7256 2084 7364
rect 2222 7352 2228 7364
rect 2280 7352 2286 7404
rect 2498 7392 2504 7404
rect 2459 7364 2504 7392
rect 2498 7352 2504 7364
rect 2556 7352 2562 7404
rect 2682 7392 2688 7404
rect 2643 7364 2688 7392
rect 2682 7352 2688 7364
rect 2740 7352 2746 7404
rect 2314 7284 2320 7336
rect 2372 7324 2378 7336
rect 2700 7324 2728 7352
rect 2372 7296 2728 7324
rect 3344 7324 3372 7432
rect 3712 7432 4804 7460
rect 3602 7352 3608 7404
rect 3660 7392 3666 7404
rect 3712 7401 3740 7432
rect 4798 7420 4804 7432
rect 4856 7420 4862 7472
rect 5368 7460 5396 7488
rect 8110 7460 8116 7472
rect 5368 7432 6868 7460
rect 3697 7395 3755 7401
rect 3697 7392 3709 7395
rect 3660 7364 3709 7392
rect 3660 7352 3666 7364
rect 3697 7361 3709 7364
rect 3743 7361 3755 7395
rect 3697 7355 3755 7361
rect 3973 7395 4031 7401
rect 3973 7361 3985 7395
rect 4019 7361 4031 7395
rect 3973 7355 4031 7361
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7392 4215 7395
rect 4522 7392 4528 7404
rect 4203 7364 4528 7392
rect 4203 7361 4215 7364
rect 4157 7355 4215 7361
rect 3988 7324 4016 7355
rect 4522 7352 4528 7364
rect 4580 7352 4586 7404
rect 5353 7395 5411 7401
rect 5353 7361 5365 7395
rect 5399 7361 5411 7395
rect 5353 7355 5411 7361
rect 4982 7324 4988 7336
rect 3344 7296 4988 7324
rect 2372 7284 2378 7296
rect 4982 7284 4988 7296
rect 5040 7284 5046 7336
rect 5368 7324 5396 7355
rect 5442 7352 5448 7404
rect 5500 7392 5506 7404
rect 5629 7395 5687 7401
rect 5629 7392 5641 7395
rect 5500 7364 5641 7392
rect 5500 7352 5506 7364
rect 5629 7361 5641 7364
rect 5675 7361 5687 7395
rect 5810 7392 5816 7404
rect 5771 7364 5816 7392
rect 5629 7355 5687 7361
rect 5810 7352 5816 7364
rect 5868 7352 5874 7404
rect 6546 7392 6552 7404
rect 6507 7364 6552 7392
rect 6546 7352 6552 7364
rect 6604 7352 6610 7404
rect 6638 7352 6644 7404
rect 6696 7392 6702 7404
rect 6840 7401 6868 7432
rect 7392 7432 8116 7460
rect 7392 7401 7420 7432
rect 8110 7420 8116 7432
rect 8168 7420 8174 7472
rect 9950 7460 9956 7472
rect 9600 7432 9956 7460
rect 9600 7401 9628 7432
rect 9950 7420 9956 7432
rect 10008 7460 10014 7472
rect 11330 7460 11336 7472
rect 10008 7432 11336 7460
rect 10008 7420 10014 7432
rect 11330 7420 11336 7432
rect 11388 7460 11394 7472
rect 11876 7463 11934 7469
rect 11388 7432 11652 7460
rect 11388 7420 11394 7432
rect 6733 7395 6791 7401
rect 6733 7392 6745 7395
rect 6696 7364 6745 7392
rect 6696 7352 6702 7364
rect 6733 7361 6745 7364
rect 6779 7361 6791 7395
rect 6733 7355 6791 7361
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7361 6883 7395
rect 6825 7355 6883 7361
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 7644 7395 7702 7401
rect 7644 7361 7656 7395
rect 7690 7392 7702 7395
rect 9585 7395 9643 7401
rect 7690 7364 9536 7392
rect 7690 7361 7702 7364
rect 7644 7355 7702 7361
rect 6914 7324 6920 7336
rect 5368 7296 6920 7324
rect 6914 7284 6920 7296
rect 6972 7284 6978 7336
rect 5994 7256 6000 7268
rect 2056 7228 6000 7256
rect 5994 7216 6000 7228
rect 6052 7216 6058 7268
rect 6181 7259 6239 7265
rect 6181 7225 6193 7259
rect 6227 7256 6239 7259
rect 7190 7256 7196 7268
rect 6227 7228 7196 7256
rect 6227 7225 6239 7228
rect 6181 7219 6239 7225
rect 7190 7216 7196 7228
rect 7248 7256 7254 7268
rect 7392 7256 7420 7355
rect 7248 7228 7420 7256
rect 7248 7216 7254 7228
rect 1397 7191 1455 7197
rect 1397 7157 1409 7191
rect 1443 7188 1455 7191
rect 2222 7188 2228 7200
rect 1443 7160 2228 7188
rect 1443 7157 1455 7160
rect 1397 7151 1455 7157
rect 2222 7148 2228 7160
rect 2280 7148 2286 7200
rect 3513 7191 3571 7197
rect 3513 7157 3525 7191
rect 3559 7188 3571 7191
rect 3970 7188 3976 7200
rect 3559 7160 3976 7188
rect 3559 7157 3571 7160
rect 3513 7151 3571 7157
rect 3970 7148 3976 7160
rect 4028 7148 4034 7200
rect 5166 7188 5172 7200
rect 5127 7160 5172 7188
rect 5166 7148 5172 7160
rect 5224 7148 5230 7200
rect 5258 7148 5264 7200
rect 5316 7188 5322 7200
rect 6086 7188 6092 7200
rect 5316 7160 6092 7188
rect 5316 7148 5322 7160
rect 6086 7148 6092 7160
rect 6144 7188 6150 7200
rect 9398 7188 9404 7200
rect 6144 7160 9404 7188
rect 6144 7148 6150 7160
rect 9398 7148 9404 7160
rect 9456 7148 9462 7200
rect 9508 7188 9536 7364
rect 9585 7361 9597 7395
rect 9631 7361 9643 7395
rect 9585 7355 9643 7361
rect 9852 7395 9910 7401
rect 9852 7361 9864 7395
rect 9898 7392 9910 7395
rect 10226 7392 10232 7404
rect 9898 7364 10232 7392
rect 9898 7361 9910 7364
rect 9852 7355 9910 7361
rect 10226 7352 10232 7364
rect 10284 7352 10290 7404
rect 10318 7352 10324 7404
rect 10376 7392 10382 7404
rect 11514 7392 11520 7404
rect 10376 7364 11520 7392
rect 10376 7352 10382 7364
rect 11514 7352 11520 7364
rect 11572 7352 11578 7404
rect 11624 7401 11652 7432
rect 11876 7429 11888 7463
rect 11922 7460 11934 7463
rect 12342 7460 12348 7472
rect 11922 7432 12348 7460
rect 11922 7429 11934 7432
rect 11876 7423 11934 7429
rect 12342 7420 12348 7432
rect 12400 7420 12406 7472
rect 13998 7460 14004 7472
rect 13911 7432 14004 7460
rect 11609 7395 11667 7401
rect 11609 7361 11621 7395
rect 11655 7361 11667 7395
rect 11609 7355 11667 7361
rect 13633 7395 13691 7401
rect 13633 7361 13645 7395
rect 13679 7392 13691 7395
rect 13814 7392 13820 7404
rect 13679 7364 13820 7392
rect 13679 7361 13691 7364
rect 13633 7355 13691 7361
rect 13814 7352 13820 7364
rect 13872 7352 13878 7404
rect 13924 7401 13952 7432
rect 13998 7420 14004 7432
rect 14056 7460 14062 7472
rect 17954 7460 17960 7472
rect 14056 7432 15056 7460
rect 14056 7420 14062 7432
rect 15028 7404 15056 7432
rect 17328 7432 17960 7460
rect 13909 7395 13967 7401
rect 13909 7361 13921 7395
rect 13955 7361 13967 7395
rect 13909 7355 13967 7361
rect 14093 7395 14151 7401
rect 14093 7361 14105 7395
rect 14139 7392 14151 7395
rect 14274 7392 14280 7404
rect 14139 7364 14280 7392
rect 14139 7361 14151 7364
rect 14093 7355 14151 7361
rect 14274 7352 14280 7364
rect 14332 7352 14338 7404
rect 14734 7392 14740 7404
rect 14695 7364 14740 7392
rect 14734 7352 14740 7364
rect 14792 7352 14798 7404
rect 15010 7392 15016 7404
rect 14971 7364 15016 7392
rect 15010 7352 15016 7364
rect 15068 7352 15074 7404
rect 15197 7395 15255 7401
rect 15197 7361 15209 7395
rect 15243 7361 15255 7395
rect 15197 7355 15255 7361
rect 15212 7324 15240 7355
rect 15470 7352 15476 7404
rect 15528 7392 15534 7404
rect 15841 7395 15899 7401
rect 15841 7392 15853 7395
rect 15528 7364 15853 7392
rect 15528 7352 15534 7364
rect 15841 7361 15853 7364
rect 15887 7361 15899 7395
rect 16022 7392 16028 7404
rect 15983 7364 16028 7392
rect 15841 7355 15899 7361
rect 16022 7352 16028 7364
rect 16080 7352 16086 7404
rect 16853 7395 16911 7401
rect 16853 7392 16865 7395
rect 16224 7364 16865 7392
rect 15378 7324 15384 7336
rect 13004 7296 15384 7324
rect 13004 7265 13032 7296
rect 15378 7284 15384 7296
rect 15436 7324 15442 7336
rect 16117 7327 16175 7333
rect 16117 7324 16129 7327
rect 15436 7296 16129 7324
rect 15436 7284 15442 7296
rect 16117 7293 16129 7296
rect 16163 7293 16175 7327
rect 16117 7287 16175 7293
rect 12989 7259 13047 7265
rect 12989 7225 13001 7259
rect 13035 7225 13047 7259
rect 12989 7219 13047 7225
rect 13814 7216 13820 7268
rect 13872 7256 13878 7268
rect 15102 7256 15108 7268
rect 13872 7228 15108 7256
rect 13872 7216 13878 7228
rect 15102 7216 15108 7228
rect 15160 7256 15166 7268
rect 16224 7256 16252 7364
rect 16853 7361 16865 7364
rect 16899 7361 16911 7395
rect 16853 7355 16911 7361
rect 16942 7352 16948 7404
rect 17000 7392 17006 7404
rect 17328 7401 17356 7432
rect 17954 7420 17960 7432
rect 18012 7420 18018 7472
rect 18690 7420 18696 7472
rect 18748 7460 18754 7472
rect 18748 7432 21220 7460
rect 18748 7420 18754 7432
rect 17129 7395 17187 7401
rect 17129 7392 17141 7395
rect 17000 7364 17141 7392
rect 17000 7352 17006 7364
rect 17129 7361 17141 7364
rect 17175 7361 17187 7395
rect 17129 7355 17187 7361
rect 17313 7395 17371 7401
rect 17313 7361 17325 7395
rect 17359 7361 17371 7395
rect 17313 7355 17371 7361
rect 17678 7352 17684 7404
rect 17736 7392 17742 7404
rect 18049 7395 18107 7401
rect 18049 7392 18061 7395
rect 17736 7364 18061 7392
rect 17736 7352 17742 7364
rect 18049 7361 18061 7364
rect 18095 7392 18107 7395
rect 18138 7392 18144 7404
rect 18095 7364 18144 7392
rect 18095 7361 18107 7364
rect 18049 7355 18107 7361
rect 18138 7352 18144 7364
rect 18196 7352 18202 7404
rect 18322 7401 18328 7404
rect 18316 7392 18328 7401
rect 18283 7364 18328 7392
rect 18316 7355 18328 7364
rect 18322 7352 18328 7355
rect 18380 7352 18386 7404
rect 20257 7395 20315 7401
rect 20257 7361 20269 7395
rect 20303 7392 20315 7395
rect 20622 7392 20628 7404
rect 20303 7364 20628 7392
rect 20303 7361 20315 7364
rect 20257 7355 20315 7361
rect 20622 7352 20628 7364
rect 20680 7352 20686 7404
rect 19610 7284 19616 7336
rect 19668 7324 19674 7336
rect 20349 7327 20407 7333
rect 20349 7324 20361 7327
rect 19668 7296 20361 7324
rect 19668 7284 19674 7296
rect 20349 7293 20361 7296
rect 20395 7293 20407 7327
rect 20349 7287 20407 7293
rect 20533 7327 20591 7333
rect 20533 7293 20545 7327
rect 20579 7324 20591 7327
rect 20990 7324 20996 7336
rect 20579 7296 20996 7324
rect 20579 7293 20591 7296
rect 20533 7287 20591 7293
rect 15160 7228 16252 7256
rect 15160 7216 15166 7228
rect 19150 7216 19156 7268
rect 19208 7256 19214 7268
rect 20548 7256 20576 7287
rect 20990 7284 20996 7296
rect 21048 7284 21054 7336
rect 19208 7228 20576 7256
rect 21192 7256 21220 7432
rect 21358 7420 21364 7472
rect 21416 7460 21422 7472
rect 21928 7460 21956 7500
rect 22189 7497 22201 7500
rect 22235 7497 22247 7531
rect 22189 7491 22247 7497
rect 22373 7531 22431 7537
rect 22373 7497 22385 7531
rect 22419 7528 22431 7531
rect 22830 7528 22836 7540
rect 22419 7500 22836 7528
rect 22419 7497 22431 7500
rect 22373 7491 22431 7497
rect 22830 7488 22836 7500
rect 22888 7488 22894 7540
rect 26142 7488 26148 7540
rect 26200 7528 26206 7540
rect 28350 7528 28356 7540
rect 26200 7500 28356 7528
rect 26200 7488 26206 7500
rect 21416 7432 21956 7460
rect 21416 7420 21422 7432
rect 23382 7420 23388 7472
rect 23440 7460 23446 7472
rect 26970 7460 26976 7472
rect 23440 7432 25268 7460
rect 26931 7432 26976 7460
rect 23440 7420 23446 7432
rect 21269 7395 21327 7401
rect 21269 7361 21281 7395
rect 21315 7392 21327 7395
rect 22646 7392 22652 7404
rect 21315 7364 22652 7392
rect 21315 7361 21327 7364
rect 21269 7355 21327 7361
rect 22646 7352 22652 7364
rect 22704 7352 22710 7404
rect 23658 7392 23664 7404
rect 23619 7364 23664 7392
rect 23658 7352 23664 7364
rect 23716 7352 23722 7404
rect 23750 7352 23756 7404
rect 23808 7392 23814 7404
rect 24397 7395 24455 7401
rect 24397 7392 24409 7395
rect 23808 7364 23853 7392
rect 23952 7364 24409 7392
rect 23808 7352 23814 7364
rect 21634 7284 21640 7336
rect 21692 7324 21698 7336
rect 21821 7327 21879 7333
rect 21821 7324 21833 7327
rect 21692 7296 21833 7324
rect 21692 7284 21698 7296
rect 21821 7293 21833 7296
rect 21867 7293 21879 7327
rect 21821 7287 21879 7293
rect 22186 7284 22192 7336
rect 22244 7324 22250 7336
rect 22370 7324 22376 7336
rect 22244 7296 22376 7324
rect 22244 7284 22250 7296
rect 22370 7284 22376 7296
rect 22428 7284 22434 7336
rect 23290 7284 23296 7336
rect 23348 7324 23354 7336
rect 23952 7324 23980 7364
rect 24397 7361 24409 7364
rect 24443 7392 24455 7395
rect 25130 7392 25136 7404
rect 24443 7364 25136 7392
rect 24443 7361 24455 7364
rect 24397 7355 24455 7361
rect 25130 7352 25136 7364
rect 25188 7352 25194 7404
rect 24486 7324 24492 7336
rect 23348 7296 23980 7324
rect 24447 7296 24492 7324
rect 23348 7284 23354 7296
rect 24486 7284 24492 7296
rect 24544 7284 24550 7336
rect 25240 7324 25268 7432
rect 26970 7420 26976 7432
rect 27028 7420 27034 7472
rect 26050 7392 26056 7404
rect 26011 7364 26056 7392
rect 26050 7352 26056 7364
rect 26108 7352 26114 7404
rect 26145 7395 26203 7401
rect 26145 7361 26157 7395
rect 26191 7392 26203 7395
rect 26418 7392 26424 7404
rect 26191 7364 26424 7392
rect 26191 7361 26203 7364
rect 26145 7355 26203 7361
rect 26418 7352 26424 7364
rect 26476 7352 26482 7404
rect 26237 7327 26295 7333
rect 26237 7324 26249 7327
rect 25240 7296 26249 7324
rect 26237 7293 26249 7296
rect 26283 7324 26295 7327
rect 27062 7324 27068 7336
rect 26283 7296 27068 7324
rect 26283 7293 26295 7296
rect 26237 7287 26295 7293
rect 27062 7284 27068 7296
rect 27120 7284 27126 7336
rect 27430 7324 27436 7336
rect 27172 7296 27436 7324
rect 24765 7259 24823 7265
rect 24765 7256 24777 7259
rect 21192 7228 24777 7256
rect 19208 7216 19214 7228
rect 24765 7225 24777 7228
rect 24811 7256 24823 7259
rect 27172 7256 27200 7296
rect 27430 7284 27436 7296
rect 27488 7284 27494 7336
rect 24811 7228 27200 7256
rect 27341 7259 27399 7265
rect 24811 7225 24823 7228
rect 24765 7219 24823 7225
rect 27341 7225 27353 7259
rect 27387 7256 27399 7259
rect 27540 7256 27568 7500
rect 28350 7488 28356 7500
rect 28408 7488 28414 7540
rect 29270 7528 29276 7540
rect 29231 7500 29276 7528
rect 29270 7488 29276 7500
rect 29328 7528 29334 7540
rect 30282 7528 30288 7540
rect 29328 7500 30288 7528
rect 29328 7488 29334 7500
rect 30282 7488 30288 7500
rect 30340 7488 30346 7540
rect 31202 7488 31208 7540
rect 31260 7528 31266 7540
rect 31297 7531 31355 7537
rect 31297 7528 31309 7531
rect 31260 7500 31309 7528
rect 31260 7488 31266 7500
rect 31297 7497 31309 7500
rect 31343 7497 31355 7531
rect 31297 7491 31355 7497
rect 29638 7460 29644 7472
rect 27908 7432 29644 7460
rect 27908 7401 27936 7432
rect 29638 7420 29644 7432
rect 29696 7420 29702 7472
rect 30190 7469 30196 7472
rect 30184 7460 30196 7469
rect 30151 7432 30196 7460
rect 30184 7423 30196 7432
rect 30190 7420 30196 7423
rect 30248 7420 30254 7472
rect 27893 7395 27951 7401
rect 27893 7361 27905 7395
rect 27939 7361 27951 7395
rect 27893 7355 27951 7361
rect 27982 7352 27988 7404
rect 28040 7392 28046 7404
rect 28149 7395 28207 7401
rect 28149 7392 28161 7395
rect 28040 7364 28161 7392
rect 28040 7352 28046 7364
rect 28149 7361 28161 7364
rect 28195 7361 28207 7395
rect 28149 7355 28207 7361
rect 29638 7284 29644 7336
rect 29696 7324 29702 7336
rect 29914 7324 29920 7336
rect 29696 7296 29920 7324
rect 29696 7284 29702 7296
rect 29914 7284 29920 7296
rect 29972 7284 29978 7336
rect 27387 7228 27568 7256
rect 27387 7225 27399 7228
rect 27341 7219 27399 7225
rect 10318 7188 10324 7200
rect 9508 7160 10324 7188
rect 10318 7148 10324 7160
rect 10376 7148 10382 7200
rect 10594 7148 10600 7200
rect 10652 7188 10658 7200
rect 12894 7188 12900 7200
rect 10652 7160 12900 7188
rect 10652 7148 10658 7160
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 13446 7188 13452 7200
rect 13407 7160 13452 7188
rect 13446 7148 13452 7160
rect 13504 7148 13510 7200
rect 14734 7148 14740 7200
rect 14792 7188 14798 7200
rect 15930 7188 15936 7200
rect 14792 7160 15936 7188
rect 14792 7148 14798 7160
rect 15930 7148 15936 7160
rect 15988 7148 15994 7200
rect 16298 7148 16304 7200
rect 16356 7188 16362 7200
rect 19242 7188 19248 7200
rect 16356 7160 19248 7188
rect 16356 7148 16362 7160
rect 19242 7148 19248 7160
rect 19300 7148 19306 7200
rect 19429 7191 19487 7197
rect 19429 7157 19441 7191
rect 19475 7188 19487 7191
rect 19794 7188 19800 7200
rect 19475 7160 19800 7188
rect 19475 7157 19487 7160
rect 19429 7151 19487 7157
rect 19794 7148 19800 7160
rect 19852 7148 19858 7200
rect 19889 7191 19947 7197
rect 19889 7157 19901 7191
rect 19935 7188 19947 7191
rect 20898 7188 20904 7200
rect 19935 7160 20904 7188
rect 19935 7157 19947 7160
rect 19889 7151 19947 7157
rect 20898 7148 20904 7160
rect 20956 7148 20962 7200
rect 21634 7148 21640 7200
rect 21692 7188 21698 7200
rect 22189 7191 22247 7197
rect 22189 7188 22201 7191
rect 21692 7160 22201 7188
rect 21692 7148 21698 7160
rect 22189 7157 22201 7160
rect 22235 7157 22247 7191
rect 22189 7151 22247 7157
rect 25498 7148 25504 7200
rect 25556 7188 25562 7200
rect 25685 7191 25743 7197
rect 25685 7188 25697 7191
rect 25556 7160 25697 7188
rect 25556 7148 25562 7160
rect 25685 7157 25697 7160
rect 25731 7157 25743 7191
rect 25685 7151 25743 7157
rect 27433 7191 27491 7197
rect 27433 7157 27445 7191
rect 27479 7188 27491 7191
rect 27522 7188 27528 7200
rect 27479 7160 27528 7188
rect 27479 7157 27491 7160
rect 27433 7151 27491 7157
rect 27522 7148 27528 7160
rect 27580 7148 27586 7200
rect 27614 7148 27620 7200
rect 27672 7188 27678 7200
rect 28166 7188 28172 7200
rect 27672 7160 28172 7188
rect 27672 7148 27678 7160
rect 28166 7148 28172 7160
rect 28224 7148 28230 7200
rect 1104 7098 32016 7120
rect 1104 7046 2136 7098
rect 2188 7046 12440 7098
rect 12492 7046 22744 7098
rect 22796 7046 32016 7098
rect 1104 7024 32016 7046
rect 1302 6944 1308 6996
rect 1360 6984 1366 6996
rect 3602 6984 3608 6996
rect 1360 6956 3608 6984
rect 1360 6944 1366 6956
rect 3602 6944 3608 6956
rect 3660 6944 3666 6996
rect 4062 6944 4068 6996
rect 4120 6984 4126 6996
rect 5534 6984 5540 6996
rect 4120 6956 5540 6984
rect 4120 6944 4126 6956
rect 5534 6944 5540 6956
rect 5592 6944 5598 6996
rect 8110 6984 8116 6996
rect 8071 6956 8116 6984
rect 8110 6944 8116 6956
rect 8168 6944 8174 6996
rect 10226 6984 10232 6996
rect 10187 6956 10232 6984
rect 10226 6944 10232 6956
rect 10284 6944 10290 6996
rect 12894 6944 12900 6996
rect 12952 6984 12958 6996
rect 12952 6956 15976 6984
rect 12952 6944 12958 6956
rect 2406 6876 2412 6928
rect 2464 6916 2470 6928
rect 2777 6919 2835 6925
rect 2777 6916 2789 6919
rect 2464 6888 2789 6916
rect 2464 6876 2470 6888
rect 2777 6885 2789 6888
rect 2823 6916 2835 6919
rect 2823 6888 4292 6916
rect 2823 6885 2835 6888
rect 2777 6879 2835 6885
rect 4264 6857 4292 6888
rect 4614 6876 4620 6928
rect 4672 6916 4678 6928
rect 4798 6916 4804 6928
rect 4672 6888 4804 6916
rect 4672 6876 4678 6888
rect 4798 6876 4804 6888
rect 4856 6876 4862 6928
rect 10594 6916 10600 6928
rect 8312 6888 10600 6916
rect 4157 6851 4215 6857
rect 4157 6848 4169 6851
rect 3160 6820 4169 6848
rect 1394 6780 1400 6792
rect 1355 6752 1400 6780
rect 1394 6740 1400 6752
rect 1452 6740 1458 6792
rect 3160 6780 3188 6820
rect 4157 6817 4169 6820
rect 4203 6817 4215 6851
rect 4157 6811 4215 6817
rect 4249 6851 4307 6857
rect 4249 6817 4261 6851
rect 4295 6817 4307 6851
rect 4249 6811 4307 6817
rect 3970 6780 3976 6792
rect 2332 6752 3188 6780
rect 3931 6752 3976 6780
rect 2332 6724 2360 6752
rect 3970 6740 3976 6752
rect 4028 6740 4034 6792
rect 4264 6780 4292 6811
rect 4338 6808 4344 6860
rect 4396 6848 4402 6860
rect 8312 6848 8340 6888
rect 10594 6876 10600 6888
rect 10652 6876 10658 6928
rect 12713 6919 12771 6925
rect 12713 6885 12725 6919
rect 12759 6916 12771 6919
rect 12802 6916 12808 6928
rect 12759 6888 12808 6916
rect 12759 6885 12771 6888
rect 12713 6879 12771 6885
rect 12802 6876 12808 6888
rect 12860 6916 12866 6928
rect 14274 6916 14280 6928
rect 12860 6888 14280 6916
rect 12860 6876 12866 6888
rect 14274 6876 14280 6888
rect 14332 6916 14338 6928
rect 15948 6916 15976 6956
rect 17126 6944 17132 6996
rect 17184 6984 17190 6996
rect 17770 6984 17776 6996
rect 17184 6956 17776 6984
rect 17184 6944 17190 6956
rect 17770 6944 17776 6956
rect 17828 6944 17834 6996
rect 19337 6987 19395 6993
rect 19337 6953 19349 6987
rect 19383 6984 19395 6987
rect 19426 6984 19432 6996
rect 19383 6956 19432 6984
rect 19383 6953 19395 6956
rect 19337 6947 19395 6953
rect 19426 6944 19432 6956
rect 19484 6944 19490 6996
rect 21634 6984 21640 6996
rect 19536 6956 21220 6984
rect 21595 6956 21640 6984
rect 19536 6916 19564 6956
rect 14332 6888 15148 6916
rect 15948 6888 19564 6916
rect 21192 6916 21220 6956
rect 21634 6944 21640 6956
rect 21692 6944 21698 6996
rect 22278 6944 22284 6996
rect 22336 6984 22342 6996
rect 22557 6987 22615 6993
rect 22557 6984 22569 6987
rect 22336 6956 22569 6984
rect 22336 6944 22342 6956
rect 22557 6953 22569 6956
rect 22603 6953 22615 6987
rect 22557 6947 22615 6953
rect 22646 6944 22652 6996
rect 22704 6984 22710 6996
rect 22741 6987 22799 6993
rect 22741 6984 22753 6987
rect 22704 6956 22753 6984
rect 22704 6944 22710 6956
rect 22741 6953 22753 6956
rect 22787 6953 22799 6987
rect 22741 6947 22799 6953
rect 23198 6944 23204 6996
rect 23256 6984 23262 6996
rect 23569 6987 23627 6993
rect 23569 6984 23581 6987
rect 23256 6956 23581 6984
rect 23256 6944 23262 6956
rect 23569 6953 23581 6956
rect 23615 6953 23627 6987
rect 23569 6947 23627 6953
rect 23753 6987 23811 6993
rect 23753 6953 23765 6987
rect 23799 6984 23811 6987
rect 24486 6984 24492 6996
rect 23799 6956 24492 6984
rect 23799 6953 23811 6956
rect 23753 6947 23811 6953
rect 24486 6944 24492 6956
rect 24544 6944 24550 6996
rect 25958 6944 25964 6996
rect 26016 6984 26022 6996
rect 27338 6984 27344 6996
rect 26016 6956 27344 6984
rect 26016 6944 26022 6956
rect 27338 6944 27344 6956
rect 27396 6944 27402 6996
rect 32125 6919 32183 6925
rect 32125 6916 32137 6919
rect 21192 6888 32137 6916
rect 14332 6876 14338 6888
rect 4396 6820 8340 6848
rect 4396 6808 4402 6820
rect 8754 6808 8760 6860
rect 8812 6848 8818 6860
rect 8941 6851 8999 6857
rect 8941 6848 8953 6851
rect 8812 6820 8953 6848
rect 8812 6808 8818 6820
rect 8941 6817 8953 6820
rect 8987 6817 8999 6851
rect 8941 6811 8999 6817
rect 9217 6851 9275 6857
rect 9217 6817 9229 6851
rect 9263 6848 9275 6851
rect 9766 6848 9772 6860
rect 9263 6820 9772 6848
rect 9263 6817 9275 6820
rect 9217 6811 9275 6817
rect 9766 6808 9772 6820
rect 9824 6848 9830 6860
rect 10689 6851 10747 6857
rect 10689 6848 10701 6851
rect 9824 6820 10701 6848
rect 9824 6808 9830 6820
rect 10689 6817 10701 6820
rect 10735 6817 10747 6851
rect 11330 6848 11336 6860
rect 11291 6820 11336 6848
rect 10689 6811 10747 6817
rect 11330 6808 11336 6820
rect 11388 6808 11394 6860
rect 13449 6851 13507 6857
rect 13449 6848 13461 6851
rect 13280 6820 13461 6848
rect 4614 6780 4620 6792
rect 4264 6752 4620 6780
rect 4614 6740 4620 6752
rect 4672 6740 4678 6792
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6780 5135 6783
rect 5258 6780 5264 6792
rect 5123 6752 5264 6780
rect 5123 6749 5135 6752
rect 5077 6743 5135 6749
rect 5258 6740 5264 6752
rect 5316 6740 5322 6792
rect 5353 6783 5411 6789
rect 5353 6749 5365 6783
rect 5399 6780 5411 6783
rect 5442 6780 5448 6792
rect 5399 6752 5448 6780
rect 5399 6749 5411 6752
rect 5353 6743 5411 6749
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 10226 6780 10232 6792
rect 5552 6752 10232 6780
rect 1664 6715 1722 6721
rect 1664 6681 1676 6715
rect 1710 6712 1722 6715
rect 1762 6712 1768 6724
rect 1710 6684 1768 6712
rect 1710 6681 1722 6684
rect 1664 6675 1722 6681
rect 1762 6672 1768 6684
rect 1820 6672 1826 6724
rect 2314 6672 2320 6724
rect 2372 6672 2378 6724
rect 5552 6712 5580 6752
rect 10226 6740 10232 6752
rect 10284 6740 10290 6792
rect 10410 6780 10416 6792
rect 10371 6752 10416 6780
rect 10410 6740 10416 6752
rect 10468 6740 10474 6792
rect 10594 6780 10600 6792
rect 10555 6752 10600 6780
rect 10594 6740 10600 6752
rect 10652 6740 10658 6792
rect 11974 6740 11980 6792
rect 12032 6780 12038 6792
rect 13078 6780 13084 6792
rect 12032 6752 13084 6780
rect 12032 6740 12038 6752
rect 13078 6740 13084 6752
rect 13136 6740 13142 6792
rect 13280 6780 13308 6820
rect 13449 6817 13461 6820
rect 13495 6848 13507 6851
rect 14458 6848 14464 6860
rect 13495 6820 14464 6848
rect 13495 6817 13507 6820
rect 13449 6811 13507 6817
rect 14458 6808 14464 6820
rect 14516 6808 14522 6860
rect 14553 6851 14611 6857
rect 14553 6817 14565 6851
rect 14599 6848 14611 6851
rect 14734 6848 14740 6860
rect 14599 6820 14740 6848
rect 14599 6817 14611 6820
rect 14553 6811 14611 6817
rect 14734 6808 14740 6820
rect 14792 6808 14798 6860
rect 15010 6848 15016 6860
rect 14971 6820 15016 6848
rect 15010 6808 15016 6820
rect 15068 6808 15074 6860
rect 15120 6848 15148 6888
rect 32125 6885 32137 6888
rect 32171 6885 32183 6919
rect 32125 6879 32183 6885
rect 15289 6851 15347 6857
rect 15289 6848 15301 6851
rect 15120 6820 15301 6848
rect 15289 6817 15301 6820
rect 15335 6817 15347 6851
rect 15289 6811 15347 6817
rect 15378 6808 15384 6860
rect 15436 6857 15442 6860
rect 15436 6851 15464 6857
rect 15452 6817 15464 6851
rect 15436 6811 15464 6817
rect 15565 6851 15623 6857
rect 15565 6817 15577 6851
rect 15611 6848 15623 6851
rect 15746 6848 15752 6860
rect 15611 6820 15752 6848
rect 15611 6817 15623 6820
rect 15565 6811 15623 6817
rect 15436 6808 15442 6811
rect 15746 6808 15752 6820
rect 15804 6808 15810 6860
rect 16761 6851 16819 6857
rect 16761 6817 16773 6851
rect 16807 6848 16819 6851
rect 18049 6851 18107 6857
rect 18049 6848 18061 6851
rect 16807 6820 18061 6848
rect 16807 6817 16819 6820
rect 16761 6811 16819 6817
rect 18049 6817 18061 6820
rect 18095 6817 18107 6851
rect 19702 6848 19708 6860
rect 19663 6820 19708 6848
rect 18049 6811 18107 6817
rect 19702 6808 19708 6820
rect 19760 6808 19766 6860
rect 22922 6808 22928 6860
rect 22980 6848 22986 6860
rect 25498 6848 25504 6860
rect 22980 6820 24716 6848
rect 25459 6820 25504 6848
rect 22980 6808 22986 6820
rect 14366 6780 14372 6792
rect 13188 6752 13308 6780
rect 14327 6752 14372 6780
rect 6638 6712 6644 6724
rect 4172 6684 5580 6712
rect 6599 6684 6644 6712
rect 3050 6604 3056 6656
rect 3108 6644 3114 6656
rect 3789 6647 3847 6653
rect 3789 6644 3801 6647
rect 3108 6616 3801 6644
rect 3108 6604 3114 6616
rect 3789 6613 3801 6616
rect 3835 6613 3847 6647
rect 3789 6607 3847 6613
rect 3878 6604 3884 6656
rect 3936 6644 3942 6656
rect 4172 6644 4200 6684
rect 6638 6672 6644 6684
rect 6696 6712 6702 6724
rect 11600 6715 11658 6721
rect 6696 6684 9674 6712
rect 6696 6672 6702 6684
rect 3936 6616 4200 6644
rect 3936 6604 3942 6616
rect 4246 6604 4252 6656
rect 4304 6644 4310 6656
rect 7374 6644 7380 6656
rect 4304 6616 7380 6644
rect 4304 6604 4310 6616
rect 7374 6604 7380 6616
rect 7432 6604 7438 6656
rect 9646 6644 9674 6684
rect 11600 6681 11612 6715
rect 11646 6712 11658 6715
rect 12250 6712 12256 6724
rect 11646 6684 12256 6712
rect 11646 6681 11658 6684
rect 11600 6675 11658 6681
rect 12250 6672 12256 6684
rect 12308 6672 12314 6724
rect 11882 6644 11888 6656
rect 9646 6616 11888 6644
rect 11882 6604 11888 6616
rect 11940 6644 11946 6656
rect 13188 6644 13216 6752
rect 14366 6740 14372 6752
rect 14424 6740 14430 6792
rect 16209 6783 16267 6789
rect 16209 6749 16221 6783
rect 16255 6780 16267 6783
rect 16482 6780 16488 6792
rect 16255 6752 16488 6780
rect 16255 6749 16267 6752
rect 16209 6743 16267 6749
rect 16482 6740 16488 6752
rect 16540 6740 16546 6792
rect 16942 6780 16948 6792
rect 16903 6752 16948 6780
rect 16942 6740 16948 6752
rect 17000 6740 17006 6792
rect 17126 6780 17132 6792
rect 17087 6752 17132 6780
rect 17126 6740 17132 6752
rect 17184 6740 17190 6792
rect 17221 6783 17279 6789
rect 17221 6749 17233 6783
rect 17267 6780 17279 6783
rect 17310 6780 17316 6792
rect 17267 6752 17316 6780
rect 17267 6749 17279 6752
rect 17221 6743 17279 6749
rect 13265 6715 13323 6721
rect 13265 6681 13277 6715
rect 13311 6681 13323 6715
rect 13265 6675 13323 6681
rect 16040 6684 16528 6712
rect 11940 6616 13216 6644
rect 13280 6644 13308 6675
rect 16040 6656 16068 6684
rect 15838 6644 15844 6656
rect 13280 6616 15844 6644
rect 11940 6604 11946 6616
rect 15838 6604 15844 6616
rect 15896 6604 15902 6656
rect 16022 6604 16028 6656
rect 16080 6604 16086 6656
rect 16500 6644 16528 6684
rect 16574 6672 16580 6724
rect 16632 6712 16638 6724
rect 17236 6712 17264 6743
rect 17310 6740 17316 6752
rect 17368 6780 17374 6792
rect 17678 6780 17684 6792
rect 17368 6752 17684 6780
rect 17368 6740 17374 6752
rect 17678 6740 17684 6752
rect 17736 6740 17742 6792
rect 17862 6780 17868 6792
rect 17823 6752 17868 6780
rect 17862 6740 17868 6752
rect 17920 6740 17926 6792
rect 17954 6740 17960 6792
rect 18012 6780 18018 6792
rect 18141 6783 18199 6789
rect 18141 6780 18153 6783
rect 18012 6752 18153 6780
rect 18012 6740 18018 6752
rect 18141 6749 18153 6752
rect 18187 6749 18199 6783
rect 19518 6780 19524 6792
rect 19479 6752 19524 6780
rect 18141 6743 18199 6749
rect 19518 6740 19524 6752
rect 19576 6740 19582 6792
rect 19794 6780 19800 6792
rect 19755 6752 19800 6780
rect 19794 6740 19800 6752
rect 19852 6740 19858 6792
rect 20257 6783 20315 6789
rect 20257 6749 20269 6783
rect 20303 6780 20315 6783
rect 22094 6780 22100 6792
rect 20303 6752 22100 6780
rect 20303 6749 20315 6752
rect 20257 6743 20315 6749
rect 22094 6740 22100 6752
rect 22152 6740 22158 6792
rect 23201 6783 23259 6789
rect 23201 6749 23213 6783
rect 23247 6780 23259 6783
rect 23290 6780 23296 6792
rect 23247 6752 23296 6780
rect 23247 6749 23259 6752
rect 23201 6743 23259 6749
rect 23290 6740 23296 6752
rect 23348 6740 23354 6792
rect 24578 6780 24584 6792
rect 24539 6752 24584 6780
rect 24578 6740 24584 6752
rect 24636 6740 24642 6792
rect 24688 6780 24716 6820
rect 25498 6808 25504 6820
rect 25556 6808 25562 6860
rect 25593 6851 25651 6857
rect 25593 6817 25605 6851
rect 25639 6817 25651 6851
rect 25593 6811 25651 6817
rect 25608 6780 25636 6811
rect 27062 6808 27068 6860
rect 27120 6848 27126 6860
rect 27157 6851 27215 6857
rect 27157 6848 27169 6851
rect 27120 6820 27169 6848
rect 27120 6808 27126 6820
rect 27157 6817 27169 6820
rect 27203 6817 27215 6851
rect 27157 6811 27215 6817
rect 28258 6808 28264 6860
rect 28316 6848 28322 6860
rect 28353 6851 28411 6857
rect 28353 6848 28365 6851
rect 28316 6820 28365 6848
rect 28316 6808 28322 6820
rect 28353 6817 28365 6820
rect 28399 6817 28411 6851
rect 29730 6848 29736 6860
rect 29691 6820 29736 6848
rect 28353 6811 28411 6817
rect 29730 6808 29736 6820
rect 29788 6808 29794 6860
rect 30742 6848 30748 6860
rect 30208 6820 30748 6848
rect 24688 6752 25636 6780
rect 27246 6740 27252 6792
rect 27304 6780 27310 6792
rect 27982 6780 27988 6792
rect 27304 6752 27988 6780
rect 27304 6740 27310 6752
rect 27982 6740 27988 6752
rect 28040 6780 28046 6792
rect 30208 6789 30236 6820
rect 30742 6808 30748 6820
rect 30800 6808 30806 6860
rect 31110 6808 31116 6860
rect 31168 6848 31174 6860
rect 31297 6851 31355 6857
rect 31297 6848 31309 6851
rect 31168 6820 31309 6848
rect 31168 6808 31174 6820
rect 31297 6817 31309 6820
rect 31343 6817 31355 6851
rect 31297 6811 31355 6817
rect 28077 6783 28135 6789
rect 28077 6780 28089 6783
rect 28040 6752 28089 6780
rect 28040 6740 28046 6752
rect 28077 6749 28089 6752
rect 28123 6749 28135 6783
rect 28077 6743 28135 6749
rect 29917 6783 29975 6789
rect 29917 6749 29929 6783
rect 29963 6749 29975 6783
rect 29917 6743 29975 6749
rect 30193 6783 30251 6789
rect 30193 6749 30205 6783
rect 30239 6749 30251 6783
rect 30193 6743 30251 6749
rect 19886 6712 19892 6724
rect 16632 6684 17264 6712
rect 17328 6684 19892 6712
rect 16632 6672 16638 6684
rect 17328 6644 17356 6684
rect 19886 6672 19892 6684
rect 19944 6672 19950 6724
rect 20524 6715 20582 6721
rect 20524 6681 20536 6715
rect 20570 6712 20582 6715
rect 21818 6712 21824 6724
rect 20570 6684 21824 6712
rect 20570 6681 20582 6684
rect 20524 6675 20582 6681
rect 21818 6672 21824 6684
rect 21876 6672 21882 6724
rect 22373 6715 22431 6721
rect 22373 6681 22385 6715
rect 22419 6681 22431 6715
rect 22373 6675 22431 6681
rect 22589 6715 22647 6721
rect 22589 6681 22601 6715
rect 22635 6712 22647 6715
rect 25409 6715 25467 6721
rect 22635 6684 23152 6712
rect 22635 6681 22647 6684
rect 22589 6675 22647 6681
rect 16500 6616 17356 6644
rect 17681 6647 17739 6653
rect 17681 6613 17693 6647
rect 17727 6644 17739 6647
rect 21082 6644 21088 6656
rect 17727 6616 21088 6644
rect 17727 6613 17739 6616
rect 17681 6607 17739 6613
rect 21082 6604 21088 6616
rect 21140 6604 21146 6656
rect 22388 6644 22416 6675
rect 22830 6644 22836 6656
rect 22388 6616 22836 6644
rect 22830 6604 22836 6616
rect 22888 6604 22894 6656
rect 23124 6644 23152 6684
rect 25409 6681 25421 6715
rect 25455 6712 25467 6715
rect 26973 6715 27031 6721
rect 25455 6684 26648 6712
rect 25455 6681 25467 6684
rect 25409 6675 25467 6681
rect 23578 6647 23636 6653
rect 23578 6644 23590 6647
rect 23124 6616 23590 6644
rect 23578 6613 23590 6616
rect 23624 6644 23636 6647
rect 24397 6647 24455 6653
rect 24397 6644 24409 6647
rect 23624 6616 24409 6644
rect 23624 6613 23636 6616
rect 23578 6607 23636 6613
rect 24397 6613 24409 6616
rect 24443 6613 24455 6647
rect 25038 6644 25044 6656
rect 24999 6616 25044 6644
rect 24397 6607 24455 6613
rect 25038 6604 25044 6616
rect 25096 6604 25102 6656
rect 26620 6653 26648 6684
rect 26973 6681 26985 6715
rect 27019 6712 27031 6715
rect 28994 6712 29000 6724
rect 27019 6684 29000 6712
rect 27019 6681 27031 6684
rect 26973 6675 27031 6681
rect 28994 6672 29000 6684
rect 29052 6672 29058 6724
rect 29932 6712 29960 6743
rect 30282 6740 30288 6792
rect 30340 6780 30346 6792
rect 30377 6783 30435 6789
rect 30377 6780 30389 6783
rect 30340 6752 30389 6780
rect 30340 6740 30346 6752
rect 30377 6749 30389 6752
rect 30423 6749 30435 6783
rect 30377 6743 30435 6749
rect 30558 6740 30564 6792
rect 30616 6780 30622 6792
rect 31021 6783 31079 6789
rect 31021 6780 31033 6783
rect 30616 6752 31033 6780
rect 30616 6740 30622 6752
rect 31021 6749 31033 6752
rect 31067 6749 31079 6783
rect 31021 6743 31079 6749
rect 31205 6783 31263 6789
rect 31205 6749 31217 6783
rect 31251 6780 31263 6783
rect 31386 6780 31392 6792
rect 31251 6752 31392 6780
rect 31251 6749 31263 6752
rect 31205 6743 31263 6749
rect 31386 6740 31392 6752
rect 31444 6740 31450 6792
rect 30466 6712 30472 6724
rect 29932 6684 30472 6712
rect 30466 6672 30472 6684
rect 30524 6672 30530 6724
rect 26605 6647 26663 6653
rect 26605 6613 26617 6647
rect 26651 6613 26663 6647
rect 26605 6607 26663 6613
rect 27065 6647 27123 6653
rect 27065 6613 27077 6647
rect 27111 6644 27123 6647
rect 27706 6644 27712 6656
rect 27111 6616 27712 6644
rect 27111 6613 27123 6616
rect 27065 6607 27123 6613
rect 27706 6604 27712 6616
rect 27764 6604 27770 6656
rect 30190 6604 30196 6656
rect 30248 6644 30254 6656
rect 30837 6647 30895 6653
rect 30837 6644 30849 6647
rect 30248 6616 30849 6644
rect 30248 6604 30254 6616
rect 30837 6613 30849 6616
rect 30883 6613 30895 6647
rect 30837 6607 30895 6613
rect 1104 6554 32016 6576
rect 1104 6502 7288 6554
rect 7340 6502 17592 6554
rect 17644 6502 27896 6554
rect 27948 6502 32016 6554
rect 1104 6480 32016 6502
rect 1762 6440 1768 6452
rect 1723 6412 1768 6440
rect 1762 6400 1768 6412
rect 1820 6400 1826 6452
rect 2406 6400 2412 6452
rect 2464 6440 2470 6452
rect 2866 6440 2872 6452
rect 2464 6412 2872 6440
rect 2464 6400 2470 6412
rect 2866 6400 2872 6412
rect 2924 6400 2930 6452
rect 4154 6400 4160 6452
rect 4212 6440 4218 6452
rect 4525 6443 4583 6449
rect 4525 6440 4537 6443
rect 4212 6412 4537 6440
rect 4212 6400 4218 6412
rect 4525 6409 4537 6412
rect 4571 6409 4583 6443
rect 4525 6403 4583 6409
rect 4614 6400 4620 6452
rect 4672 6440 4678 6452
rect 5629 6443 5687 6449
rect 5629 6440 5641 6443
rect 4672 6412 5641 6440
rect 4672 6400 4678 6412
rect 5629 6409 5641 6412
rect 5675 6409 5687 6443
rect 10318 6440 10324 6452
rect 10279 6412 10324 6440
rect 5629 6403 5687 6409
rect 10318 6400 10324 6412
rect 10376 6400 10382 6452
rect 10410 6400 10416 6452
rect 10468 6440 10474 6452
rect 12250 6440 12256 6452
rect 10468 6412 11744 6440
rect 12211 6412 12256 6440
rect 10468 6400 10474 6412
rect 0 6372 800 6386
rect 2498 6372 2504 6384
rect 0 6344 2504 6372
rect 0 6330 800 6344
rect 2498 6332 2504 6344
rect 2556 6332 2562 6384
rect 3237 6375 3295 6381
rect 3237 6341 3249 6375
rect 3283 6372 3295 6375
rect 6638 6372 6644 6384
rect 3283 6344 6644 6372
rect 3283 6341 3295 6344
rect 3237 6335 3295 6341
rect 6638 6332 6644 6344
rect 6696 6332 6702 6384
rect 9217 6375 9275 6381
rect 9217 6341 9229 6375
rect 9263 6372 9275 6375
rect 9263 6344 10548 6372
rect 9263 6341 9275 6344
rect 9217 6335 9275 6341
rect 1210 6264 1216 6316
rect 1268 6304 1274 6316
rect 1762 6304 1768 6316
rect 1268 6276 1768 6304
rect 1268 6264 1274 6276
rect 1762 6264 1768 6276
rect 1820 6264 1826 6316
rect 1946 6304 1952 6316
rect 1907 6276 1952 6304
rect 1946 6264 1952 6276
rect 2004 6264 2010 6316
rect 2225 6307 2283 6313
rect 2225 6273 2237 6307
rect 2271 6304 2283 6307
rect 2682 6304 2688 6316
rect 2271 6276 2688 6304
rect 2271 6273 2283 6276
rect 2225 6267 2283 6273
rect 2682 6264 2688 6276
rect 2740 6264 2746 6316
rect 4430 6264 4436 6316
rect 4488 6304 4494 6316
rect 5445 6307 5503 6313
rect 5445 6304 5457 6307
rect 4488 6276 5457 6304
rect 4488 6264 4494 6276
rect 5445 6273 5457 6276
rect 5491 6273 5503 6307
rect 5445 6267 5503 6273
rect 5721 6307 5779 6313
rect 5721 6273 5733 6307
rect 5767 6273 5779 6307
rect 5721 6267 5779 6273
rect 1486 6196 1492 6248
rect 1544 6236 1550 6248
rect 2133 6239 2191 6245
rect 2133 6236 2145 6239
rect 1544 6208 2145 6236
rect 1544 6196 1550 6208
rect 2133 6205 2145 6208
rect 2179 6236 2191 6239
rect 2314 6236 2320 6248
rect 2179 6208 2320 6236
rect 2179 6205 2191 6208
rect 2133 6199 2191 6205
rect 2314 6196 2320 6208
rect 2372 6196 2378 6248
rect 2590 6196 2596 6248
rect 2648 6236 2654 6248
rect 5736 6236 5764 6267
rect 5994 6264 6000 6316
rect 6052 6304 6058 6316
rect 7929 6307 7987 6313
rect 7929 6304 7941 6307
rect 6052 6276 7941 6304
rect 6052 6264 6058 6276
rect 6656 6245 6684 6276
rect 7929 6273 7941 6276
rect 7975 6273 7987 6307
rect 7929 6267 7987 6273
rect 8205 6307 8263 6313
rect 8205 6273 8217 6307
rect 8251 6304 8263 6307
rect 9306 6304 9312 6316
rect 8251 6276 9312 6304
rect 8251 6273 8263 6276
rect 8205 6267 8263 6273
rect 9306 6264 9312 6276
rect 9364 6304 9370 6316
rect 9401 6307 9459 6313
rect 9401 6304 9413 6307
rect 9364 6276 9413 6304
rect 9364 6264 9370 6276
rect 9401 6273 9413 6276
rect 9447 6273 9459 6307
rect 9674 6304 9680 6316
rect 9635 6276 9680 6304
rect 9401 6267 9459 6273
rect 9674 6264 9680 6276
rect 9732 6264 9738 6316
rect 9766 6264 9772 6316
rect 9824 6304 9830 6316
rect 10520 6313 10548 6344
rect 9861 6307 9919 6313
rect 9861 6304 9873 6307
rect 9824 6276 9873 6304
rect 9824 6264 9830 6276
rect 9861 6273 9873 6276
rect 9907 6273 9919 6307
rect 9861 6267 9919 6273
rect 10505 6307 10563 6313
rect 10505 6273 10517 6307
rect 10551 6273 10563 6307
rect 10505 6267 10563 6273
rect 10781 6307 10839 6313
rect 10781 6273 10793 6307
rect 10827 6304 10839 6307
rect 11514 6304 11520 6316
rect 10827 6276 11520 6304
rect 10827 6273 10839 6276
rect 10781 6267 10839 6273
rect 11514 6264 11520 6276
rect 11572 6264 11578 6316
rect 11609 6307 11667 6313
rect 11609 6273 11621 6307
rect 11655 6273 11667 6307
rect 11609 6267 11667 6273
rect 2648 6208 5764 6236
rect 6641 6239 6699 6245
rect 2648 6196 2654 6208
rect 6641 6205 6653 6239
rect 6687 6205 6699 6239
rect 6914 6236 6920 6248
rect 6875 6208 6920 6236
rect 6641 6199 6699 6205
rect 6914 6196 6920 6208
rect 6972 6196 6978 6248
rect 9692 6236 9720 6264
rect 10410 6236 10416 6248
rect 9692 6208 10416 6236
rect 10410 6196 10416 6208
rect 10468 6196 10474 6248
rect 8938 6128 8944 6180
rect 8996 6168 9002 6180
rect 11624 6168 11652 6267
rect 11716 6236 11744 6412
rect 12250 6400 12256 6412
rect 12308 6400 12314 6452
rect 13078 6400 13084 6452
rect 13136 6440 13142 6452
rect 14182 6440 14188 6452
rect 13136 6412 14188 6440
rect 13136 6400 13142 6412
rect 14182 6400 14188 6412
rect 14240 6400 14246 6452
rect 14918 6440 14924 6452
rect 14879 6412 14924 6440
rect 14918 6400 14924 6412
rect 14976 6400 14982 6452
rect 15010 6400 15016 6452
rect 15068 6440 15074 6452
rect 15378 6440 15384 6452
rect 15068 6412 15384 6440
rect 15068 6400 15074 6412
rect 15378 6400 15384 6412
rect 15436 6400 15442 6452
rect 16669 6443 16727 6449
rect 15580 6412 16436 6440
rect 12437 6307 12495 6313
rect 12437 6273 12449 6307
rect 12483 6304 12495 6307
rect 13446 6304 13452 6316
rect 12483 6276 13452 6304
rect 12483 6273 12495 6276
rect 12437 6267 12495 6273
rect 13446 6264 13452 6276
rect 13504 6264 13510 6316
rect 13814 6304 13820 6316
rect 13775 6276 13820 6304
rect 13814 6264 13820 6276
rect 13872 6264 13878 6316
rect 13998 6264 14004 6316
rect 14056 6304 14062 6316
rect 14093 6307 14151 6313
rect 14093 6304 14105 6307
rect 14056 6276 14105 6304
rect 14056 6264 14062 6276
rect 14093 6273 14105 6276
rect 14139 6273 14151 6307
rect 14093 6267 14151 6273
rect 14277 6307 14335 6313
rect 14277 6273 14289 6307
rect 14323 6304 14335 6307
rect 14366 6304 14372 6316
rect 14323 6276 14372 6304
rect 14323 6273 14335 6276
rect 14277 6267 14335 6273
rect 14366 6264 14372 6276
rect 14424 6264 14430 6316
rect 14734 6304 14740 6316
rect 14695 6276 14740 6304
rect 14734 6264 14740 6276
rect 14792 6264 14798 6316
rect 15580 6313 15608 6412
rect 15841 6375 15899 6381
rect 15841 6341 15853 6375
rect 15887 6372 15899 6375
rect 16114 6372 16120 6384
rect 15887 6344 16120 6372
rect 15887 6341 15899 6344
rect 15841 6335 15899 6341
rect 16114 6332 16120 6344
rect 16172 6332 16178 6384
rect 15565 6307 15623 6313
rect 15565 6273 15577 6307
rect 15611 6273 15623 6307
rect 15565 6267 15623 6273
rect 15749 6307 15807 6313
rect 15749 6273 15761 6307
rect 15795 6273 15807 6307
rect 15749 6267 15807 6273
rect 15933 6307 15991 6313
rect 15933 6273 15945 6307
rect 15979 6304 15991 6307
rect 16298 6304 16304 6316
rect 15979 6276 16304 6304
rect 15979 6273 15991 6276
rect 15933 6267 15991 6273
rect 12618 6236 12624 6248
rect 11716 6208 12434 6236
rect 12579 6208 12624 6236
rect 8996 6140 11652 6168
rect 12406 6168 12434 6208
rect 12618 6196 12624 6208
rect 12676 6196 12682 6248
rect 12713 6239 12771 6245
rect 12713 6205 12725 6239
rect 12759 6236 12771 6239
rect 12805 6239 12863 6245
rect 12805 6236 12817 6239
rect 12759 6208 12817 6236
rect 12759 6205 12771 6208
rect 12713 6199 12771 6205
rect 12805 6205 12817 6208
rect 12851 6205 12863 6239
rect 12805 6199 12863 6205
rect 13633 6239 13691 6245
rect 13633 6205 13645 6239
rect 13679 6236 13691 6239
rect 15470 6236 15476 6248
rect 13679 6208 15476 6236
rect 13679 6205 13691 6208
rect 13633 6199 13691 6205
rect 15470 6196 15476 6208
rect 15528 6196 15534 6248
rect 15764 6236 15792 6267
rect 16298 6264 16304 6276
rect 16356 6264 16362 6316
rect 16408 6304 16436 6412
rect 16669 6409 16681 6443
rect 16715 6440 16727 6443
rect 17954 6440 17960 6452
rect 16715 6412 17960 6440
rect 16715 6409 16727 6412
rect 16669 6403 16727 6409
rect 17954 6400 17960 6412
rect 18012 6400 18018 6452
rect 18138 6400 18144 6452
rect 18196 6440 18202 6452
rect 19705 6443 19763 6449
rect 19705 6440 19717 6443
rect 18196 6412 19717 6440
rect 18196 6400 18202 6412
rect 19705 6409 19717 6412
rect 19751 6409 19763 6443
rect 19705 6403 19763 6409
rect 19886 6400 19892 6452
rect 19944 6440 19950 6452
rect 22186 6440 22192 6452
rect 19944 6412 22192 6440
rect 19944 6400 19950 6412
rect 22186 6400 22192 6412
rect 22244 6400 22250 6452
rect 27062 6440 27068 6452
rect 22287 6412 27068 6440
rect 16482 6332 16488 6384
rect 16540 6372 16546 6384
rect 17218 6372 17224 6384
rect 16540 6344 17080 6372
rect 16540 6332 16546 6344
rect 16758 6304 16764 6316
rect 16408 6276 16764 6304
rect 16758 6264 16764 6276
rect 16816 6264 16822 6316
rect 17052 6313 17080 6344
rect 17144 6344 17224 6372
rect 17144 6313 17172 6344
rect 17218 6332 17224 6344
rect 17276 6332 17282 6384
rect 16945 6307 17003 6313
rect 16945 6273 16957 6307
rect 16991 6273 17003 6307
rect 16945 6267 17003 6273
rect 17037 6307 17095 6313
rect 17037 6273 17049 6307
rect 17083 6273 17095 6307
rect 17037 6267 17095 6273
rect 17129 6307 17187 6313
rect 17129 6273 17141 6307
rect 17175 6273 17187 6307
rect 17310 6304 17316 6316
rect 17271 6276 17316 6304
rect 17129 6267 17187 6273
rect 16022 6236 16028 6248
rect 15764 6208 16028 6236
rect 16022 6196 16028 6208
rect 16080 6196 16086 6248
rect 16960 6236 16988 6267
rect 17310 6264 17316 6276
rect 17368 6264 17374 6316
rect 17678 6264 17684 6316
rect 17736 6304 17742 6316
rect 17773 6307 17831 6313
rect 17773 6304 17785 6307
rect 17736 6276 17785 6304
rect 17736 6264 17742 6276
rect 17773 6273 17785 6276
rect 17819 6273 17831 6307
rect 17773 6267 17831 6273
rect 18417 6307 18475 6313
rect 18417 6273 18429 6307
rect 18463 6304 18475 6307
rect 21726 6304 21732 6316
rect 18463 6276 21732 6304
rect 18463 6273 18475 6276
rect 18417 6267 18475 6273
rect 21726 6264 21732 6276
rect 21784 6264 21790 6316
rect 17862 6236 17868 6248
rect 16960 6208 17868 6236
rect 17862 6196 17868 6208
rect 17920 6196 17926 6248
rect 17954 6196 17960 6248
rect 18012 6236 18018 6248
rect 20625 6239 20683 6245
rect 20625 6236 20637 6239
rect 18012 6208 20637 6236
rect 18012 6196 18018 6208
rect 20625 6205 20637 6208
rect 20671 6205 20683 6239
rect 22287 6236 22315 6412
rect 27062 6400 27068 6412
rect 27120 6400 27126 6452
rect 27430 6400 27436 6452
rect 27488 6400 27494 6452
rect 27709 6443 27767 6449
rect 27709 6409 27721 6443
rect 27755 6440 27767 6443
rect 29270 6440 29276 6452
rect 27755 6412 29276 6440
rect 27755 6409 27767 6412
rect 27709 6403 27767 6409
rect 29270 6400 29276 6412
rect 29328 6400 29334 6452
rect 30374 6400 30380 6452
rect 30432 6440 30438 6452
rect 30469 6443 30527 6449
rect 30469 6440 30481 6443
rect 30432 6412 30481 6440
rect 30432 6400 30438 6412
rect 30469 6409 30481 6412
rect 30515 6409 30527 6443
rect 30469 6403 30527 6409
rect 26694 6332 26700 6384
rect 26752 6372 26758 6384
rect 27448 6372 27476 6400
rect 32320 6372 33120 6386
rect 26752 6344 27200 6372
rect 27448 6344 33120 6372
rect 26752 6332 26758 6344
rect 22462 6304 22468 6316
rect 22423 6276 22468 6304
rect 22462 6264 22468 6276
rect 22520 6264 22526 6316
rect 23661 6307 23719 6313
rect 23661 6273 23673 6307
rect 23707 6304 23719 6307
rect 24397 6307 24455 6313
rect 24397 6304 24409 6307
rect 23707 6276 24409 6304
rect 23707 6273 23719 6276
rect 23661 6267 23719 6273
rect 24397 6273 24409 6276
rect 24443 6273 24455 6307
rect 24397 6267 24455 6273
rect 24486 6264 24492 6316
rect 24544 6304 24550 6316
rect 24581 6307 24639 6313
rect 24581 6304 24593 6307
rect 24544 6276 24593 6304
rect 24544 6264 24550 6276
rect 24581 6273 24593 6276
rect 24627 6273 24639 6307
rect 24854 6304 24860 6316
rect 24815 6276 24860 6304
rect 24581 6267 24639 6273
rect 24854 6264 24860 6276
rect 24912 6264 24918 6316
rect 24946 6264 24952 6316
rect 25004 6304 25010 6316
rect 25041 6307 25099 6313
rect 25041 6304 25053 6307
rect 25004 6276 25053 6304
rect 25004 6264 25010 6276
rect 25041 6273 25053 6276
rect 25087 6273 25099 6307
rect 25590 6304 25596 6316
rect 25551 6276 25596 6304
rect 25041 6267 25099 6273
rect 25590 6264 25596 6276
rect 25648 6264 25654 6316
rect 25774 6304 25780 6316
rect 25735 6276 25780 6304
rect 25774 6264 25780 6276
rect 25832 6264 25838 6316
rect 25869 6307 25927 6313
rect 25869 6273 25881 6307
rect 25915 6273 25927 6307
rect 25869 6267 25927 6273
rect 20625 6199 20683 6205
rect 20732 6208 22315 6236
rect 22741 6239 22799 6245
rect 20732 6168 20760 6208
rect 22741 6205 22753 6239
rect 22787 6236 22799 6239
rect 22830 6236 22836 6248
rect 22787 6208 22836 6236
rect 22787 6205 22799 6208
rect 22741 6199 22799 6205
rect 22830 6196 22836 6208
rect 22888 6196 22894 6248
rect 23937 6239 23995 6245
rect 23937 6205 23949 6239
rect 23983 6236 23995 6239
rect 25682 6236 25688 6248
rect 23983 6208 25688 6236
rect 23983 6205 23995 6208
rect 23937 6199 23995 6205
rect 25682 6196 25688 6208
rect 25740 6196 25746 6248
rect 20898 6168 20904 6180
rect 12406 6140 20760 6168
rect 20859 6140 20904 6168
rect 8996 6128 9002 6140
rect 20898 6128 20904 6140
rect 20956 6128 20962 6180
rect 24578 6128 24584 6180
rect 24636 6168 24642 6180
rect 25884 6168 25912 6267
rect 25958 6264 25964 6316
rect 26016 6304 26022 6316
rect 26510 6304 26516 6316
rect 26016 6276 26516 6304
rect 26016 6264 26022 6276
rect 26510 6264 26516 6276
rect 26568 6264 26574 6316
rect 27172 6313 27200 6344
rect 32320 6330 33120 6344
rect 26973 6307 27031 6313
rect 26973 6273 26985 6307
rect 27019 6273 27031 6307
rect 26973 6267 27031 6273
rect 27157 6307 27215 6313
rect 27157 6273 27169 6307
rect 27203 6273 27215 6307
rect 27157 6267 27215 6273
rect 27249 6307 27307 6313
rect 27249 6273 27261 6307
rect 27295 6273 27307 6307
rect 27249 6267 27307 6273
rect 26988 6236 27016 6267
rect 27264 6236 27292 6267
rect 27338 6264 27344 6316
rect 27396 6313 27402 6316
rect 27396 6307 27445 6313
rect 27396 6273 27399 6307
rect 27433 6304 27445 6307
rect 27433 6273 27476 6304
rect 27396 6266 27476 6273
rect 27396 6264 27402 6266
rect 27982 6264 27988 6316
rect 28040 6304 28046 6316
rect 28169 6307 28227 6313
rect 28169 6304 28181 6307
rect 28040 6276 28181 6304
rect 28040 6264 28046 6276
rect 28169 6273 28181 6276
rect 28215 6273 28227 6307
rect 29178 6304 29184 6316
rect 29139 6276 29184 6304
rect 28169 6267 28227 6273
rect 29178 6264 29184 6276
rect 29236 6264 29242 6316
rect 30466 6264 30472 6316
rect 30524 6304 30530 6316
rect 30653 6307 30711 6313
rect 30653 6304 30665 6307
rect 30524 6276 30665 6304
rect 30524 6264 30530 6276
rect 30653 6273 30665 6276
rect 30699 6273 30711 6307
rect 30653 6267 30711 6273
rect 30742 6264 30748 6316
rect 30800 6304 30806 6316
rect 30929 6307 30987 6313
rect 30929 6304 30941 6307
rect 30800 6276 30941 6304
rect 30800 6264 30806 6276
rect 30929 6273 30941 6276
rect 30975 6273 30987 6307
rect 30929 6267 30987 6273
rect 31113 6307 31171 6313
rect 31113 6273 31125 6307
rect 31159 6304 31171 6307
rect 31294 6304 31300 6316
rect 31159 6276 31300 6304
rect 31159 6273 31171 6276
rect 31113 6267 31171 6273
rect 31294 6264 31300 6276
rect 31352 6264 31358 6316
rect 27614 6236 27620 6248
rect 26988 6208 27108 6236
rect 27264 6208 27620 6236
rect 24636 6140 25912 6168
rect 27080 6168 27108 6208
rect 27614 6196 27620 6208
rect 27672 6196 27678 6248
rect 29457 6239 29515 6245
rect 29457 6205 29469 6239
rect 29503 6236 29515 6239
rect 30760 6236 30788 6264
rect 29503 6208 30788 6236
rect 29503 6205 29515 6208
rect 29457 6199 29515 6205
rect 27709 6171 27767 6177
rect 27709 6168 27721 6171
rect 27080 6140 27721 6168
rect 24636 6128 24642 6140
rect 27709 6137 27721 6140
rect 27755 6137 27767 6171
rect 27709 6131 27767 6137
rect 28353 6171 28411 6177
rect 28353 6137 28365 6171
rect 28399 6168 28411 6171
rect 29730 6168 29736 6180
rect 28399 6140 29736 6168
rect 28399 6137 28411 6140
rect 28353 6131 28411 6137
rect 29730 6128 29736 6140
rect 29788 6128 29794 6180
rect 1486 6060 1492 6112
rect 1544 6100 1550 6112
rect 4338 6100 4344 6112
rect 1544 6072 4344 6100
rect 1544 6060 1550 6072
rect 4338 6060 4344 6072
rect 4396 6060 4402 6112
rect 4706 6060 4712 6112
rect 4764 6100 4770 6112
rect 5445 6103 5503 6109
rect 5445 6100 5457 6103
rect 4764 6072 5457 6100
rect 4764 6060 4770 6072
rect 5445 6069 5457 6072
rect 5491 6069 5503 6103
rect 5445 6063 5503 6069
rect 10594 6060 10600 6112
rect 10652 6100 10658 6112
rect 10689 6103 10747 6109
rect 10689 6100 10701 6103
rect 10652 6072 10701 6100
rect 10652 6060 10658 6072
rect 10689 6069 10701 6072
rect 10735 6100 10747 6103
rect 11701 6103 11759 6109
rect 11701 6100 11713 6103
rect 10735 6072 11713 6100
rect 10735 6069 10747 6072
rect 10689 6063 10747 6069
rect 11701 6069 11713 6072
rect 11747 6069 11759 6103
rect 11701 6063 11759 6069
rect 12805 6103 12863 6109
rect 12805 6069 12817 6103
rect 12851 6100 12863 6103
rect 13814 6100 13820 6112
rect 12851 6072 13820 6100
rect 12851 6069 12863 6072
rect 12805 6063 12863 6069
rect 13814 6060 13820 6072
rect 13872 6060 13878 6112
rect 15010 6060 15016 6112
rect 15068 6100 15074 6112
rect 15930 6100 15936 6112
rect 15068 6072 15936 6100
rect 15068 6060 15074 6072
rect 15930 6060 15936 6072
rect 15988 6060 15994 6112
rect 16117 6103 16175 6109
rect 16117 6069 16129 6103
rect 16163 6100 16175 6103
rect 16574 6100 16580 6112
rect 16163 6072 16580 6100
rect 16163 6069 16175 6072
rect 16117 6063 16175 6069
rect 16574 6060 16580 6072
rect 16632 6060 16638 6112
rect 16850 6060 16856 6112
rect 16908 6100 16914 6112
rect 17954 6100 17960 6112
rect 16908 6072 17960 6100
rect 16908 6060 16914 6072
rect 17954 6060 17960 6072
rect 18012 6060 18018 6112
rect 20714 6060 20720 6112
rect 20772 6100 20778 6112
rect 21085 6103 21143 6109
rect 21085 6100 21097 6103
rect 20772 6072 21097 6100
rect 20772 6060 20778 6072
rect 21085 6069 21097 6072
rect 21131 6069 21143 6103
rect 21085 6063 21143 6069
rect 22094 6060 22100 6112
rect 22152 6100 22158 6112
rect 22281 6103 22339 6109
rect 22281 6100 22293 6103
rect 22152 6072 22293 6100
rect 22152 6060 22158 6072
rect 22281 6069 22293 6072
rect 22327 6069 22339 6103
rect 22646 6100 22652 6112
rect 22607 6072 22652 6100
rect 22281 6063 22339 6069
rect 22646 6060 22652 6072
rect 22704 6060 22710 6112
rect 23474 6100 23480 6112
rect 23435 6072 23480 6100
rect 23474 6060 23480 6072
rect 23532 6060 23538 6112
rect 23750 6060 23756 6112
rect 23808 6100 23814 6112
rect 23845 6103 23903 6109
rect 23845 6100 23857 6103
rect 23808 6072 23857 6100
rect 23808 6060 23814 6072
rect 23845 6069 23857 6072
rect 23891 6069 23903 6103
rect 23845 6063 23903 6069
rect 25774 6060 25780 6112
rect 25832 6100 25838 6112
rect 26145 6103 26203 6109
rect 26145 6100 26157 6103
rect 25832 6072 26157 6100
rect 25832 6060 25838 6072
rect 26145 6069 26157 6072
rect 26191 6069 26203 6103
rect 26145 6063 26203 6069
rect 27062 6060 27068 6112
rect 27120 6100 27126 6112
rect 27525 6103 27583 6109
rect 27525 6100 27537 6103
rect 27120 6072 27537 6100
rect 27120 6060 27126 6072
rect 27525 6069 27537 6072
rect 27571 6069 27583 6103
rect 27525 6063 27583 6069
rect 28626 6060 28632 6112
rect 28684 6100 28690 6112
rect 30650 6100 30656 6112
rect 28684 6072 30656 6100
rect 28684 6060 28690 6072
rect 30650 6060 30656 6072
rect 30708 6060 30714 6112
rect 1104 6010 32016 6032
rect 1104 5958 2136 6010
rect 2188 5958 12440 6010
rect 12492 5958 22744 6010
rect 22796 5958 32016 6010
rect 1104 5936 32016 5958
rect 1486 5856 1492 5908
rect 1544 5896 1550 5908
rect 1581 5899 1639 5905
rect 1581 5896 1593 5899
rect 1544 5868 1593 5896
rect 1544 5856 1550 5868
rect 1581 5865 1593 5868
rect 1627 5865 1639 5899
rect 1581 5859 1639 5865
rect 1949 5899 2007 5905
rect 1949 5865 1961 5899
rect 1995 5896 2007 5899
rect 1995 5868 24164 5896
rect 1995 5865 2007 5868
rect 1949 5859 2007 5865
rect 1397 5695 1455 5701
rect 1397 5661 1409 5695
rect 1443 5692 1455 5695
rect 1964 5692 1992 5859
rect 2317 5831 2375 5837
rect 2317 5797 2329 5831
rect 2363 5828 2375 5831
rect 2406 5828 2412 5840
rect 2363 5800 2412 5828
rect 2363 5797 2375 5800
rect 2317 5791 2375 5797
rect 2406 5788 2412 5800
rect 2464 5788 2470 5840
rect 3145 5831 3203 5837
rect 2884 5800 3087 5828
rect 2777 5763 2835 5769
rect 2777 5729 2789 5763
rect 2823 5760 2835 5763
rect 2884 5760 2912 5800
rect 2823 5732 2912 5760
rect 3059 5760 3087 5800
rect 3145 5797 3157 5831
rect 3191 5828 3203 5831
rect 3602 5828 3608 5840
rect 3191 5800 3608 5828
rect 3191 5797 3203 5800
rect 3145 5791 3203 5797
rect 3602 5788 3608 5800
rect 3660 5828 3666 5840
rect 3878 5828 3884 5840
rect 3660 5800 3884 5828
rect 3660 5788 3666 5800
rect 3878 5788 3884 5800
rect 3936 5788 3942 5840
rect 4709 5831 4767 5837
rect 4709 5797 4721 5831
rect 4755 5828 4767 5831
rect 5074 5828 5080 5840
rect 4755 5800 5080 5828
rect 4755 5797 4767 5800
rect 4709 5791 4767 5797
rect 5074 5788 5080 5800
rect 5132 5788 5138 5840
rect 6362 5788 6368 5840
rect 6420 5828 6426 5840
rect 6457 5831 6515 5837
rect 6457 5828 6469 5831
rect 6420 5800 6469 5828
rect 6420 5788 6426 5800
rect 6457 5797 6469 5800
rect 6503 5797 6515 5831
rect 8389 5831 8447 5837
rect 8389 5828 8401 5831
rect 6457 5791 6515 5797
rect 6564 5800 8401 5828
rect 4338 5760 4344 5772
rect 3059 5732 3188 5760
rect 2823 5729 2835 5732
rect 2777 5723 2835 5729
rect 1443 5664 1992 5692
rect 3160 5692 3188 5732
rect 3436 5732 4344 5760
rect 3436 5692 3464 5732
rect 4338 5720 4344 5732
rect 4396 5720 4402 5772
rect 6086 5720 6092 5772
rect 6144 5760 6150 5772
rect 6564 5760 6592 5800
rect 8389 5797 8401 5800
rect 8435 5797 8447 5831
rect 8389 5791 8447 5797
rect 11517 5831 11575 5837
rect 11517 5797 11529 5831
rect 11563 5828 11575 5831
rect 11698 5828 11704 5840
rect 11563 5800 11704 5828
rect 11563 5797 11575 5800
rect 11517 5791 11575 5797
rect 11698 5788 11704 5800
rect 11756 5788 11762 5840
rect 12618 5788 12624 5840
rect 12676 5828 12682 5840
rect 12894 5828 12900 5840
rect 12676 5800 12900 5828
rect 12676 5788 12682 5800
rect 12894 5788 12900 5800
rect 12952 5828 12958 5840
rect 12989 5831 13047 5837
rect 12989 5828 13001 5831
rect 12952 5800 13001 5828
rect 12952 5788 12958 5800
rect 12989 5797 13001 5800
rect 13035 5797 13047 5831
rect 12989 5791 13047 5797
rect 14645 5831 14703 5837
rect 14645 5797 14657 5831
rect 14691 5828 14703 5831
rect 16577 5831 16635 5837
rect 14691 5800 16068 5828
rect 14691 5797 14703 5800
rect 14645 5791 14703 5797
rect 7466 5760 7472 5772
rect 6144 5732 6592 5760
rect 7427 5732 7472 5760
rect 6144 5720 6150 5732
rect 7466 5720 7472 5732
rect 7524 5720 7530 5772
rect 9490 5760 9496 5772
rect 9451 5732 9496 5760
rect 9490 5720 9496 5732
rect 9548 5720 9554 5772
rect 9950 5720 9956 5772
rect 10008 5760 10014 5772
rect 10137 5763 10195 5769
rect 10137 5760 10149 5763
rect 10008 5732 10149 5760
rect 10008 5720 10014 5732
rect 10137 5729 10149 5732
rect 10183 5729 10195 5763
rect 13538 5760 13544 5772
rect 10137 5723 10195 5729
rect 12406 5732 13544 5760
rect 3160 5664 3464 5692
rect 4157 5695 4215 5701
rect 1443 5661 1455 5664
rect 1397 5655 1455 5661
rect 4157 5661 4169 5695
rect 4203 5661 4215 5695
rect 4157 5655 4215 5661
rect 2133 5627 2191 5633
rect 2133 5593 2145 5627
rect 2179 5624 2191 5627
rect 2682 5624 2688 5636
rect 2179 5596 2688 5624
rect 2179 5593 2191 5596
rect 2133 5587 2191 5593
rect 2682 5584 2688 5596
rect 2740 5584 2746 5636
rect 4172 5624 4200 5655
rect 4246 5652 4252 5704
rect 4304 5692 4310 5704
rect 5077 5695 5135 5701
rect 5077 5692 5089 5695
rect 4304 5664 5089 5692
rect 4304 5652 4310 5664
rect 5077 5661 5089 5664
rect 5123 5692 5135 5695
rect 5626 5692 5632 5704
rect 5123 5664 5632 5692
rect 5123 5661 5135 5664
rect 5077 5655 5135 5661
rect 5626 5652 5632 5664
rect 5684 5652 5690 5704
rect 8205 5695 8263 5701
rect 8205 5661 8217 5695
rect 8251 5692 8263 5695
rect 8938 5692 8944 5704
rect 8251 5664 8944 5692
rect 8251 5661 8263 5664
rect 8205 5655 8263 5661
rect 8938 5652 8944 5664
rect 8996 5652 9002 5704
rect 9398 5692 9404 5704
rect 9359 5664 9404 5692
rect 9398 5652 9404 5664
rect 9456 5652 9462 5704
rect 10404 5695 10462 5701
rect 10404 5661 10416 5695
rect 10450 5661 10462 5695
rect 11974 5692 11980 5704
rect 11935 5664 11980 5692
rect 10404 5655 10462 5661
rect 5350 5633 5356 5636
rect 4709 5627 4767 5633
rect 4709 5624 4721 5627
rect 4172 5596 4721 5624
rect 4709 5593 4721 5596
rect 4755 5593 4767 5627
rect 4709 5587 4767 5593
rect 5344 5587 5356 5633
rect 5408 5624 5414 5636
rect 5408 5596 5444 5624
rect 5350 5584 5356 5587
rect 5408 5584 5414 5596
rect 5534 5584 5540 5636
rect 5592 5624 5598 5636
rect 7285 5627 7343 5633
rect 7285 5624 7297 5627
rect 5592 5596 7297 5624
rect 5592 5584 5598 5596
rect 7285 5593 7297 5596
rect 7331 5593 7343 5627
rect 7285 5587 7343 5593
rect 7374 5584 7380 5636
rect 7432 5624 7438 5636
rect 7432 5596 7477 5624
rect 7432 5584 7438 5596
rect 8662 5584 8668 5636
rect 8720 5624 8726 5636
rect 9309 5627 9367 5633
rect 9309 5624 9321 5627
rect 8720 5596 9321 5624
rect 8720 5584 8726 5596
rect 9309 5593 9321 5596
rect 9355 5593 9367 5627
rect 10428 5624 10456 5655
rect 11974 5652 11980 5664
rect 12032 5652 12038 5704
rect 12161 5695 12219 5701
rect 12161 5661 12173 5695
rect 12207 5692 12219 5695
rect 12406 5692 12434 5732
rect 13538 5720 13544 5732
rect 13596 5760 13602 5772
rect 15010 5760 15016 5772
rect 13596 5732 15016 5760
rect 13596 5720 13602 5732
rect 15010 5720 15016 5732
rect 15068 5720 15074 5772
rect 15930 5760 15936 5772
rect 15120 5732 15936 5760
rect 12802 5692 12808 5704
rect 12207 5664 12434 5692
rect 12763 5664 12808 5692
rect 12207 5661 12219 5664
rect 12161 5655 12219 5661
rect 12802 5652 12808 5664
rect 12860 5652 12866 5704
rect 13078 5692 13084 5704
rect 13039 5664 13084 5692
rect 13078 5652 13084 5664
rect 13136 5652 13142 5704
rect 14829 5695 14887 5701
rect 14829 5661 14841 5695
rect 14875 5661 14887 5695
rect 14829 5655 14887 5661
rect 10502 5624 10508 5636
rect 10428 5596 10508 5624
rect 9309 5587 9367 5593
rect 10502 5584 10508 5596
rect 10560 5584 10566 5636
rect 12069 5627 12127 5633
rect 12069 5593 12081 5627
rect 12115 5624 12127 5627
rect 13170 5624 13176 5636
rect 12115 5596 13176 5624
rect 12115 5593 12127 5596
rect 12069 5587 12127 5593
rect 13170 5584 13176 5596
rect 13228 5584 13234 5636
rect 14844 5624 14872 5655
rect 14918 5652 14924 5704
rect 14976 5692 14982 5704
rect 15120 5701 15148 5732
rect 15930 5720 15936 5732
rect 15988 5720 15994 5772
rect 16040 5760 16068 5800
rect 16577 5797 16589 5831
rect 16623 5828 16635 5831
rect 16942 5828 16948 5840
rect 16623 5800 16948 5828
rect 16623 5797 16635 5800
rect 16577 5791 16635 5797
rect 16942 5788 16948 5800
rect 17000 5788 17006 5840
rect 18233 5831 18291 5837
rect 18233 5797 18245 5831
rect 18279 5828 18291 5831
rect 19150 5828 19156 5840
rect 18279 5800 19156 5828
rect 18279 5797 18291 5800
rect 18233 5791 18291 5797
rect 19150 5788 19156 5800
rect 19208 5788 19214 5840
rect 20622 5828 20628 5840
rect 20583 5800 20628 5828
rect 20622 5788 20628 5800
rect 20680 5788 20686 5840
rect 17310 5760 17316 5772
rect 16040 5732 17316 5760
rect 17310 5720 17316 5732
rect 17368 5720 17374 5772
rect 17865 5763 17923 5769
rect 17865 5729 17877 5763
rect 17911 5760 17923 5763
rect 17954 5760 17960 5772
rect 17911 5732 17960 5760
rect 17911 5729 17923 5732
rect 17865 5723 17923 5729
rect 17954 5720 17960 5732
rect 18012 5720 18018 5772
rect 24136 5760 24164 5868
rect 24486 5856 24492 5908
rect 24544 5896 24550 5908
rect 24544 5868 25544 5896
rect 24544 5856 24550 5868
rect 25516 5828 25544 5868
rect 25682 5856 25688 5908
rect 25740 5896 25746 5908
rect 25961 5899 26019 5905
rect 25961 5896 25973 5899
rect 25740 5868 25973 5896
rect 25740 5856 25746 5868
rect 25961 5865 25973 5868
rect 26007 5865 26019 5899
rect 27706 5896 27712 5908
rect 27667 5868 27712 5896
rect 25961 5859 26019 5865
rect 27706 5856 27712 5868
rect 27764 5856 27770 5908
rect 28074 5856 28080 5908
rect 28132 5896 28138 5908
rect 29917 5899 29975 5905
rect 29917 5896 29929 5899
rect 28132 5868 29929 5896
rect 28132 5856 28138 5868
rect 29917 5865 29929 5868
rect 29963 5865 29975 5899
rect 29917 5859 29975 5865
rect 30469 5899 30527 5905
rect 30469 5865 30481 5899
rect 30515 5896 30527 5899
rect 31018 5896 31024 5908
rect 30515 5868 31024 5896
rect 30515 5865 30527 5868
rect 30469 5859 30527 5865
rect 31018 5856 31024 5868
rect 31076 5856 31082 5908
rect 26326 5828 26332 5840
rect 25516 5800 26332 5828
rect 26326 5788 26332 5800
rect 26384 5828 26390 5840
rect 26421 5831 26479 5837
rect 26421 5828 26433 5831
rect 26384 5800 26433 5828
rect 26384 5788 26390 5800
rect 26421 5797 26433 5800
rect 26467 5797 26479 5831
rect 29822 5828 29828 5840
rect 26421 5791 26479 5797
rect 27264 5800 29828 5828
rect 24136 5732 24716 5760
rect 15105 5695 15163 5701
rect 14976 5664 15021 5692
rect 14976 5652 14982 5664
rect 15105 5661 15117 5695
rect 15151 5661 15163 5695
rect 15105 5655 15163 5661
rect 15197 5695 15255 5701
rect 15197 5661 15209 5695
rect 15243 5692 15255 5695
rect 15289 5695 15347 5701
rect 15289 5692 15301 5695
rect 15243 5664 15301 5692
rect 15243 5661 15255 5664
rect 15197 5655 15255 5661
rect 15289 5661 15301 5664
rect 15335 5661 15347 5695
rect 15654 5692 15660 5704
rect 15615 5664 15660 5692
rect 15289 5655 15347 5661
rect 15654 5652 15660 5664
rect 15712 5652 15718 5704
rect 15746 5652 15752 5704
rect 15804 5692 15810 5704
rect 15841 5695 15899 5701
rect 15841 5692 15853 5695
rect 15804 5664 15853 5692
rect 15804 5652 15810 5664
rect 15841 5661 15853 5664
rect 15887 5661 15899 5695
rect 15841 5655 15899 5661
rect 16761 5695 16819 5701
rect 16761 5661 16773 5695
rect 16807 5661 16819 5695
rect 17034 5692 17040 5704
rect 16995 5664 17040 5692
rect 16761 5655 16819 5661
rect 16298 5624 16304 5636
rect 14844 5596 16304 5624
rect 16298 5584 16304 5596
rect 16356 5584 16362 5636
rect 16776 5624 16804 5655
rect 17034 5652 17040 5664
rect 17092 5652 17098 5704
rect 17221 5695 17279 5701
rect 17221 5661 17233 5695
rect 17267 5692 17279 5695
rect 19245 5695 19303 5701
rect 17267 5664 17908 5692
rect 17267 5661 17279 5664
rect 17221 5655 17279 5661
rect 17880 5636 17908 5664
rect 19245 5661 19257 5695
rect 19291 5692 19303 5695
rect 21821 5695 21879 5701
rect 21821 5692 21833 5695
rect 19291 5664 21833 5692
rect 19291 5661 19303 5664
rect 19245 5655 19303 5661
rect 21821 5661 21833 5664
rect 21867 5692 21879 5695
rect 21910 5692 21916 5704
rect 21867 5664 21916 5692
rect 21867 5661 21879 5664
rect 21821 5655 21879 5661
rect 21910 5652 21916 5664
rect 21968 5652 21974 5704
rect 22094 5701 22100 5704
rect 22088 5655 22100 5701
rect 22152 5692 22158 5704
rect 22152 5664 22188 5692
rect 22094 5652 22100 5655
rect 22152 5652 22158 5664
rect 24026 5652 24032 5704
rect 24084 5692 24090 5704
rect 24581 5695 24639 5701
rect 24581 5692 24593 5695
rect 24084 5664 24593 5692
rect 24084 5652 24090 5664
rect 24581 5661 24593 5664
rect 24627 5661 24639 5695
rect 24688 5692 24716 5732
rect 25406 5692 25412 5704
rect 24688 5664 25412 5692
rect 24581 5655 24639 5661
rect 25406 5652 25412 5664
rect 25464 5652 25470 5704
rect 26602 5692 26608 5704
rect 26515 5664 26608 5692
rect 26602 5652 26608 5664
rect 26660 5692 26666 5704
rect 26697 5695 26755 5701
rect 26697 5692 26709 5695
rect 26660 5664 26709 5692
rect 26660 5652 26666 5664
rect 26697 5661 26709 5664
rect 26743 5661 26755 5695
rect 27062 5692 27068 5704
rect 27120 5701 27126 5704
rect 27264 5701 27292 5800
rect 29822 5788 29828 5800
rect 29880 5788 29886 5840
rect 28718 5760 28724 5772
rect 28460 5732 28724 5760
rect 27030 5664 27068 5692
rect 26697 5655 26755 5661
rect 27062 5652 27068 5664
rect 27120 5655 27130 5701
rect 27213 5695 27292 5701
rect 27213 5661 27225 5695
rect 27259 5661 27292 5695
rect 27213 5660 27292 5661
rect 27213 5655 27271 5660
rect 27120 5652 27126 5655
rect 27522 5652 27528 5704
rect 27580 5701 27586 5704
rect 27580 5692 27588 5701
rect 27580 5664 27625 5692
rect 27580 5655 27588 5664
rect 27580 5652 27586 5655
rect 17310 5624 17316 5636
rect 16776 5596 17316 5624
rect 17310 5584 17316 5596
rect 17368 5584 17374 5636
rect 17862 5584 17868 5636
rect 17920 5584 17926 5636
rect 19512 5627 19570 5633
rect 19512 5593 19524 5627
rect 19558 5624 19570 5627
rect 19702 5624 19708 5636
rect 19558 5596 19708 5624
rect 19558 5593 19570 5596
rect 19512 5587 19570 5593
rect 19702 5584 19708 5596
rect 19760 5584 19766 5636
rect 21177 5627 21235 5633
rect 21177 5593 21189 5627
rect 21223 5624 21235 5627
rect 22554 5624 22560 5636
rect 21223 5596 22560 5624
rect 21223 5593 21235 5596
rect 21177 5587 21235 5593
rect 22554 5584 22560 5596
rect 22612 5584 22618 5636
rect 23658 5584 23664 5636
rect 23716 5624 23722 5636
rect 24826 5627 24884 5633
rect 24826 5624 24838 5627
rect 23716 5596 24838 5624
rect 23716 5584 23722 5596
rect 24826 5593 24838 5596
rect 24872 5593 24884 5627
rect 24826 5587 24884 5593
rect 25866 5584 25872 5636
rect 25924 5624 25930 5636
rect 26142 5624 26148 5636
rect 25924 5596 26148 5624
rect 25924 5584 25930 5596
rect 26142 5584 26148 5596
rect 26200 5624 26206 5636
rect 27341 5627 27399 5633
rect 27341 5624 27353 5627
rect 26200 5596 27353 5624
rect 26200 5584 26206 5596
rect 27341 5593 27353 5596
rect 27387 5593 27399 5627
rect 27341 5587 27399 5593
rect 27433 5627 27491 5633
rect 27433 5593 27445 5627
rect 27479 5624 27491 5627
rect 28460 5624 28488 5732
rect 28718 5720 28724 5732
rect 28776 5720 28782 5772
rect 28828 5732 30788 5760
rect 28828 5701 28856 5732
rect 30760 5704 30788 5732
rect 28537 5695 28595 5701
rect 28537 5661 28549 5695
rect 28583 5661 28595 5695
rect 28537 5655 28595 5661
rect 28813 5695 28871 5701
rect 28813 5661 28825 5695
rect 28859 5661 28871 5695
rect 28813 5655 28871 5661
rect 28997 5695 29055 5701
rect 28997 5661 29009 5695
rect 29043 5692 29055 5695
rect 29270 5692 29276 5704
rect 29043 5664 29276 5692
rect 29043 5661 29055 5664
rect 28997 5655 29055 5661
rect 27479 5596 28488 5624
rect 28552 5624 28580 5655
rect 29270 5652 29276 5664
rect 29328 5692 29334 5704
rect 29733 5695 29791 5701
rect 29328 5664 29684 5692
rect 29328 5652 29334 5664
rect 29656 5624 29684 5664
rect 29733 5661 29745 5695
rect 29779 5692 29791 5695
rect 29917 5695 29975 5701
rect 29917 5692 29929 5695
rect 29779 5664 29929 5692
rect 29779 5661 29791 5664
rect 29733 5655 29791 5661
rect 29917 5661 29929 5664
rect 29963 5661 29975 5695
rect 29917 5655 29975 5661
rect 30466 5652 30472 5704
rect 30524 5692 30530 5704
rect 30653 5695 30711 5701
rect 30653 5692 30665 5695
rect 30524 5664 30665 5692
rect 30524 5652 30530 5664
rect 30653 5661 30665 5664
rect 30699 5661 30711 5695
rect 30653 5655 30711 5661
rect 30742 5652 30748 5704
rect 30800 5692 30806 5704
rect 30929 5695 30987 5701
rect 30929 5692 30941 5695
rect 30800 5664 30941 5692
rect 30800 5652 30806 5664
rect 30929 5661 30941 5664
rect 30975 5661 30987 5695
rect 31110 5692 31116 5704
rect 31071 5664 31116 5692
rect 30929 5655 30987 5661
rect 31110 5652 31116 5664
rect 31168 5652 31174 5704
rect 30006 5624 30012 5636
rect 28552 5596 29592 5624
rect 29656 5596 30012 5624
rect 27479 5593 27491 5596
rect 27433 5587 27491 5593
rect 3234 5556 3240 5568
rect 3195 5528 3240 5556
rect 3234 5516 3240 5528
rect 3292 5516 3298 5568
rect 3786 5556 3792 5568
rect 3747 5528 3792 5556
rect 3786 5516 3792 5528
rect 3844 5516 3850 5568
rect 4249 5559 4307 5565
rect 4249 5525 4261 5559
rect 4295 5556 4307 5559
rect 4430 5556 4436 5568
rect 4295 5528 4436 5556
rect 4295 5525 4307 5528
rect 4249 5519 4307 5525
rect 4430 5516 4436 5528
rect 4488 5516 4494 5568
rect 6914 5556 6920 5568
rect 6875 5528 6920 5556
rect 6914 5516 6920 5528
rect 6972 5516 6978 5568
rect 8478 5516 8484 5568
rect 8536 5556 8542 5568
rect 8941 5559 8999 5565
rect 8941 5556 8953 5559
rect 8536 5528 8953 5556
rect 8536 5516 8542 5528
rect 8941 5525 8953 5528
rect 8987 5525 8999 5559
rect 8941 5519 8999 5525
rect 12158 5516 12164 5568
rect 12216 5556 12222 5568
rect 12621 5559 12679 5565
rect 12621 5556 12633 5559
rect 12216 5528 12633 5556
rect 12216 5516 12222 5528
rect 12621 5525 12633 5528
rect 12667 5525 12679 5559
rect 12621 5519 12679 5525
rect 15102 5516 15108 5568
rect 15160 5556 15166 5568
rect 15289 5559 15347 5565
rect 15289 5556 15301 5559
rect 15160 5528 15301 5556
rect 15160 5516 15166 5528
rect 15289 5525 15301 5528
rect 15335 5525 15347 5559
rect 15289 5519 15347 5525
rect 15378 5516 15384 5568
rect 15436 5556 15442 5568
rect 15746 5556 15752 5568
rect 15436 5528 15752 5556
rect 15436 5516 15442 5528
rect 15746 5516 15752 5528
rect 15804 5516 15810 5568
rect 16022 5556 16028 5568
rect 15935 5528 16028 5556
rect 16022 5516 16028 5528
rect 16080 5556 16086 5568
rect 17218 5556 17224 5568
rect 16080 5528 17224 5556
rect 16080 5516 16086 5528
rect 17218 5516 17224 5528
rect 17276 5516 17282 5568
rect 17954 5516 17960 5568
rect 18012 5556 18018 5568
rect 18325 5559 18383 5565
rect 18325 5556 18337 5559
rect 18012 5528 18337 5556
rect 18012 5516 18018 5528
rect 18325 5525 18337 5528
rect 18371 5525 18383 5559
rect 18325 5519 18383 5525
rect 20254 5516 20260 5568
rect 20312 5556 20318 5568
rect 21269 5559 21327 5565
rect 21269 5556 21281 5559
rect 20312 5528 21281 5556
rect 20312 5516 20318 5528
rect 21269 5525 21281 5528
rect 21315 5525 21327 5559
rect 23198 5556 23204 5568
rect 23159 5528 23204 5556
rect 21269 5519 21327 5525
rect 23198 5516 23204 5528
rect 23256 5516 23262 5568
rect 26697 5559 26755 5565
rect 26697 5525 26709 5559
rect 26743 5556 26755 5559
rect 28074 5556 28080 5568
rect 26743 5528 28080 5556
rect 26743 5525 26755 5528
rect 26697 5519 26755 5525
rect 28074 5516 28080 5528
rect 28132 5516 28138 5568
rect 28353 5559 28411 5565
rect 28353 5525 28365 5559
rect 28399 5556 28411 5559
rect 29454 5556 29460 5568
rect 28399 5528 29460 5556
rect 28399 5525 28411 5528
rect 28353 5519 28411 5525
rect 29454 5516 29460 5528
rect 29512 5516 29518 5568
rect 29564 5565 29592 5596
rect 30006 5584 30012 5596
rect 30064 5584 30070 5636
rect 29549 5559 29607 5565
rect 29549 5525 29561 5559
rect 29595 5556 29607 5559
rect 30466 5556 30472 5568
rect 29595 5528 30472 5556
rect 29595 5525 29607 5528
rect 29549 5519 29607 5525
rect 30466 5516 30472 5528
rect 30524 5516 30530 5568
rect 1104 5466 32016 5488
rect 1104 5414 7288 5466
rect 7340 5414 17592 5466
rect 17644 5414 27896 5466
rect 27948 5414 32016 5466
rect 1104 5392 32016 5414
rect 2682 5312 2688 5364
rect 2740 5352 2746 5364
rect 5350 5352 5356 5364
rect 2740 5324 5120 5352
rect 5311 5324 5356 5352
rect 2740 5312 2746 5324
rect 2314 5284 2320 5296
rect 2240 5256 2320 5284
rect 2038 5216 2044 5228
rect 1999 5188 2044 5216
rect 2038 5176 2044 5188
rect 2096 5176 2102 5228
rect 2240 5225 2268 5256
rect 2314 5244 2320 5256
rect 2372 5244 2378 5296
rect 4154 5284 4160 5296
rect 2792 5256 4160 5284
rect 2792 5225 2820 5256
rect 4154 5244 4160 5256
rect 4212 5244 4218 5296
rect 4724 5293 4752 5324
rect 4709 5287 4767 5293
rect 4709 5253 4721 5287
rect 4755 5253 4767 5287
rect 4709 5247 4767 5253
rect 4893 5287 4951 5293
rect 4893 5253 4905 5287
rect 4939 5284 4951 5287
rect 4982 5284 4988 5296
rect 4939 5256 4988 5284
rect 4939 5253 4951 5256
rect 4893 5247 4951 5253
rect 4982 5244 4988 5256
rect 5040 5244 5046 5296
rect 5092 5284 5120 5324
rect 5350 5312 5356 5324
rect 5408 5312 5414 5364
rect 6914 5312 6920 5364
rect 6972 5352 6978 5364
rect 7745 5355 7803 5361
rect 7745 5352 7757 5355
rect 6972 5324 7757 5352
rect 6972 5312 6978 5324
rect 7745 5321 7757 5324
rect 7791 5321 7803 5355
rect 7745 5315 7803 5321
rect 9033 5355 9091 5361
rect 9033 5321 9045 5355
rect 9079 5352 9091 5355
rect 9079 5324 16344 5352
rect 9079 5321 9091 5324
rect 9033 5315 9091 5321
rect 5258 5284 5264 5296
rect 5092 5256 5264 5284
rect 5258 5244 5264 5256
rect 5316 5244 5322 5296
rect 5442 5244 5448 5296
rect 5500 5284 5506 5296
rect 5500 5256 6868 5284
rect 5500 5244 5506 5256
rect 3050 5225 3056 5228
rect 2225 5219 2283 5225
rect 2225 5185 2237 5219
rect 2271 5185 2283 5219
rect 2225 5179 2283 5185
rect 2777 5219 2835 5225
rect 2777 5185 2789 5219
rect 2823 5185 2835 5219
rect 3044 5216 3056 5225
rect 3011 5188 3056 5216
rect 2777 5179 2835 5185
rect 3044 5179 3056 5188
rect 2317 5151 2375 5157
rect 2317 5117 2329 5151
rect 2363 5148 2375 5151
rect 2590 5148 2596 5160
rect 2363 5120 2596 5148
rect 2363 5117 2375 5120
rect 2317 5111 2375 5117
rect 2590 5108 2596 5120
rect 2648 5108 2654 5160
rect 1394 5040 1400 5092
rect 1452 5080 1458 5092
rect 2792 5080 2820 5179
rect 3050 5176 3056 5179
rect 3108 5176 3114 5228
rect 5537 5219 5595 5225
rect 5537 5185 5549 5219
rect 5583 5216 5595 5219
rect 6365 5219 6423 5225
rect 6365 5216 6377 5219
rect 5583 5188 6377 5216
rect 5583 5185 5595 5188
rect 5537 5179 5595 5185
rect 6365 5185 6377 5188
rect 6411 5185 6423 5219
rect 6546 5216 6552 5228
rect 6507 5188 6552 5216
rect 6365 5179 6423 5185
rect 6546 5176 6552 5188
rect 6604 5176 6610 5228
rect 6840 5225 6868 5256
rect 7834 5244 7840 5296
rect 7892 5284 7898 5296
rect 8113 5287 8171 5293
rect 8113 5284 8125 5287
rect 7892 5256 8125 5284
rect 7892 5244 7898 5256
rect 8113 5253 8125 5256
rect 8159 5253 8171 5287
rect 8478 5284 8484 5296
rect 8439 5256 8484 5284
rect 8113 5247 8171 5253
rect 8478 5244 8484 5256
rect 8536 5244 8542 5296
rect 8849 5287 8907 5293
rect 8849 5253 8861 5287
rect 8895 5284 8907 5287
rect 9398 5284 9404 5296
rect 8895 5256 9404 5284
rect 8895 5253 8907 5256
rect 8849 5247 8907 5253
rect 9398 5244 9404 5256
rect 9456 5244 9462 5296
rect 16316 5284 16344 5324
rect 16390 5312 16396 5364
rect 16448 5352 16454 5364
rect 27157 5355 27215 5361
rect 27157 5352 27169 5355
rect 16448 5324 27169 5352
rect 16448 5312 16454 5324
rect 27157 5321 27169 5324
rect 27203 5321 27215 5355
rect 27157 5315 27215 5321
rect 17037 5287 17095 5293
rect 16316 5256 16620 5284
rect 6825 5219 6883 5225
rect 6825 5185 6837 5219
rect 6871 5185 6883 5219
rect 6825 5179 6883 5185
rect 7009 5219 7067 5225
rect 7009 5185 7021 5219
rect 7055 5185 7067 5219
rect 7009 5179 7067 5185
rect 5813 5151 5871 5157
rect 5813 5117 5825 5151
rect 5859 5148 5871 5151
rect 6181 5151 6239 5157
rect 6181 5148 6193 5151
rect 5859 5120 6193 5148
rect 5859 5117 5871 5120
rect 5813 5111 5871 5117
rect 6181 5117 6193 5120
rect 6227 5117 6239 5151
rect 6181 5111 6239 5117
rect 6454 5108 6460 5160
rect 6512 5148 6518 5160
rect 7024 5148 7052 5179
rect 7926 5176 7932 5228
rect 7984 5216 7990 5228
rect 8021 5219 8079 5225
rect 8021 5216 8033 5219
rect 7984 5188 8033 5216
rect 7984 5176 7990 5188
rect 8021 5185 8033 5188
rect 8067 5185 8079 5219
rect 8021 5179 8079 5185
rect 8570 5176 8576 5228
rect 8628 5216 8634 5228
rect 10134 5216 10140 5228
rect 8628 5188 10140 5216
rect 8628 5176 8634 5188
rect 10134 5176 10140 5188
rect 10192 5216 10198 5228
rect 10502 5216 10508 5228
rect 10192 5188 10508 5216
rect 10192 5176 10198 5188
rect 10502 5176 10508 5188
rect 10560 5176 10566 5228
rect 11977 5219 12035 5225
rect 11977 5185 11989 5219
rect 12023 5216 12035 5219
rect 14001 5219 14059 5225
rect 14001 5216 14013 5219
rect 12023 5188 14013 5216
rect 12023 5185 12035 5188
rect 11977 5179 12035 5185
rect 14001 5185 14013 5188
rect 14047 5185 14059 5219
rect 14001 5179 14059 5185
rect 14185 5219 14243 5225
rect 14185 5185 14197 5219
rect 14231 5216 14243 5219
rect 14274 5216 14280 5228
rect 14231 5188 14280 5216
rect 14231 5185 14243 5188
rect 14185 5179 14243 5185
rect 14274 5176 14280 5188
rect 14332 5176 14338 5228
rect 14366 5176 14372 5228
rect 14424 5216 14430 5228
rect 14461 5219 14519 5225
rect 14461 5216 14473 5219
rect 14424 5188 14473 5216
rect 14424 5176 14430 5188
rect 14461 5185 14473 5188
rect 14507 5185 14519 5219
rect 14461 5179 14519 5185
rect 14645 5219 14703 5225
rect 14645 5185 14657 5219
rect 14691 5185 14703 5219
rect 14645 5179 14703 5185
rect 6512 5120 7052 5148
rect 8786 5120 9444 5148
rect 6512 5108 6518 5120
rect 1452 5052 2820 5080
rect 1452 5040 1458 5052
rect 3878 5040 3884 5092
rect 3936 5080 3942 5092
rect 7650 5080 7656 5092
rect 3936 5052 7656 5080
rect 3936 5040 3942 5052
rect 7650 5040 7656 5052
rect 7708 5040 7714 5092
rect 9416 5080 9444 5120
rect 9490 5108 9496 5160
rect 9548 5148 9554 5160
rect 9585 5151 9643 5157
rect 9585 5148 9597 5151
rect 9548 5120 9597 5148
rect 9548 5108 9554 5120
rect 9585 5117 9597 5120
rect 9631 5117 9643 5151
rect 9585 5111 9643 5117
rect 9861 5151 9919 5157
rect 9861 5117 9873 5151
rect 9907 5148 9919 5151
rect 9950 5148 9956 5160
rect 9907 5120 9956 5148
rect 9907 5117 9919 5120
rect 9861 5111 9919 5117
rect 9950 5108 9956 5120
rect 10008 5108 10014 5160
rect 12253 5151 12311 5157
rect 12253 5117 12265 5151
rect 12299 5148 12311 5151
rect 12618 5148 12624 5160
rect 12299 5120 12624 5148
rect 12299 5117 12311 5120
rect 12253 5111 12311 5117
rect 12618 5108 12624 5120
rect 12676 5108 12682 5160
rect 12713 5151 12771 5157
rect 12713 5117 12725 5151
rect 12759 5117 12771 5151
rect 12713 5111 12771 5117
rect 9766 5080 9772 5092
rect 9416 5052 9772 5080
rect 9766 5040 9772 5052
rect 9824 5040 9830 5092
rect 12161 5083 12219 5089
rect 12161 5049 12173 5083
rect 12207 5080 12219 5083
rect 12526 5080 12532 5092
rect 12207 5052 12532 5080
rect 12207 5049 12219 5052
rect 12161 5043 12219 5049
rect 12526 5040 12532 5052
rect 12584 5040 12590 5092
rect 1670 4972 1676 5024
rect 1728 5012 1734 5024
rect 1857 5015 1915 5021
rect 1857 5012 1869 5015
rect 1728 4984 1869 5012
rect 1728 4972 1734 4984
rect 1857 4981 1869 4984
rect 1903 4981 1915 5015
rect 1857 4975 1915 4981
rect 4062 4972 4068 5024
rect 4120 5012 4126 5024
rect 4157 5015 4215 5021
rect 4157 5012 4169 5015
rect 4120 4984 4169 5012
rect 4120 4972 4126 4984
rect 4157 4981 4169 4984
rect 4203 5012 4215 5015
rect 4522 5012 4528 5024
rect 4203 4984 4528 5012
rect 4203 4981 4215 4984
rect 4157 4975 4215 4981
rect 4522 4972 4528 4984
rect 4580 4972 4586 5024
rect 5721 5015 5779 5021
rect 5721 4981 5733 5015
rect 5767 5012 5779 5015
rect 6086 5012 6092 5024
rect 5767 4984 6092 5012
rect 5767 4981 5779 4984
rect 5721 4975 5779 4981
rect 6086 4972 6092 4984
rect 6144 4972 6150 5024
rect 6181 5015 6239 5021
rect 6181 4981 6193 5015
rect 6227 5012 6239 5015
rect 7098 5012 7104 5024
rect 6227 4984 7104 5012
rect 6227 4981 6239 4984
rect 6181 4975 6239 4981
rect 7098 4972 7104 4984
rect 7156 4972 7162 5024
rect 11790 5012 11796 5024
rect 11751 4984 11796 5012
rect 11790 4972 11796 4984
rect 11848 4972 11854 5024
rect 12728 5012 12756 5111
rect 12894 5108 12900 5160
rect 12952 5148 12958 5160
rect 12989 5151 13047 5157
rect 12989 5148 13001 5151
rect 12952 5120 13001 5148
rect 12952 5108 12958 5120
rect 12989 5117 13001 5120
rect 13035 5117 13047 5151
rect 12989 5111 13047 5117
rect 13814 5108 13820 5160
rect 13872 5148 13878 5160
rect 14660 5148 14688 5179
rect 14826 5176 14832 5228
rect 14884 5216 14890 5228
rect 15473 5219 15531 5225
rect 15473 5216 15485 5219
rect 14884 5188 15485 5216
rect 14884 5176 14890 5188
rect 15473 5185 15485 5188
rect 15519 5185 15531 5219
rect 15473 5179 15531 5185
rect 15565 5219 15623 5225
rect 15565 5185 15577 5219
rect 15611 5216 15623 5219
rect 16482 5216 16488 5228
rect 15611 5188 16488 5216
rect 15611 5185 15623 5188
rect 15565 5179 15623 5185
rect 16482 5176 16488 5188
rect 16540 5176 16546 5228
rect 14918 5148 14924 5160
rect 13872 5120 14924 5148
rect 13872 5108 13878 5120
rect 14918 5108 14924 5120
rect 14976 5108 14982 5160
rect 15102 5148 15108 5160
rect 15063 5120 15108 5148
rect 15102 5108 15108 5120
rect 15160 5108 15166 5160
rect 15289 5151 15347 5157
rect 15289 5117 15301 5151
rect 15335 5117 15347 5151
rect 15289 5111 15347 5117
rect 13998 5040 14004 5092
rect 14056 5080 14062 5092
rect 15010 5080 15016 5092
rect 14056 5052 15016 5080
rect 14056 5040 14062 5052
rect 15010 5040 15016 5052
rect 15068 5040 15074 5092
rect 15304 5080 15332 5111
rect 15378 5108 15384 5160
rect 15436 5148 15442 5160
rect 15654 5148 15660 5160
rect 15436 5120 15660 5148
rect 15436 5108 15442 5120
rect 15654 5108 15660 5120
rect 15712 5148 15718 5160
rect 16390 5148 16396 5160
rect 15712 5120 16396 5148
rect 15712 5108 15718 5120
rect 16390 5108 16396 5120
rect 16448 5108 16454 5160
rect 16592 5148 16620 5256
rect 17037 5253 17049 5287
rect 17083 5284 17095 5287
rect 18230 5284 18236 5296
rect 17083 5256 18236 5284
rect 17083 5253 17095 5256
rect 17037 5247 17095 5253
rect 18230 5244 18236 5256
rect 18288 5244 18294 5296
rect 18414 5293 18420 5296
rect 18408 5247 18420 5293
rect 18472 5284 18478 5296
rect 18472 5256 18508 5284
rect 18414 5244 18420 5247
rect 18472 5244 18478 5256
rect 19794 5244 19800 5296
rect 19852 5284 19858 5296
rect 20901 5287 20959 5293
rect 20901 5284 20913 5287
rect 19852 5256 20913 5284
rect 19852 5244 19858 5256
rect 20901 5253 20913 5256
rect 20947 5253 20959 5287
rect 20901 5247 20959 5253
rect 21082 5244 21088 5296
rect 21140 5293 21146 5296
rect 21140 5287 21159 5293
rect 21147 5253 21159 5287
rect 22370 5284 22376 5296
rect 21140 5247 21159 5253
rect 21560 5256 22376 5284
rect 21140 5244 21146 5247
rect 16669 5219 16727 5225
rect 16669 5185 16681 5219
rect 16715 5216 16727 5219
rect 16761 5219 16819 5225
rect 16761 5216 16773 5219
rect 16715 5188 16773 5216
rect 16715 5185 16727 5188
rect 16669 5179 16727 5185
rect 16761 5185 16773 5188
rect 16807 5185 16819 5219
rect 16761 5179 16819 5185
rect 16850 5176 16856 5228
rect 16908 5216 16914 5228
rect 16945 5219 17003 5225
rect 16945 5216 16957 5219
rect 16908 5188 16957 5216
rect 16908 5176 16914 5188
rect 16945 5185 16957 5188
rect 16991 5185 17003 5219
rect 16945 5179 17003 5185
rect 17129 5219 17187 5225
rect 17129 5185 17141 5219
rect 17175 5216 17187 5219
rect 17310 5216 17316 5228
rect 17175 5188 17316 5216
rect 17175 5185 17187 5188
rect 17129 5179 17187 5185
rect 17310 5176 17316 5188
rect 17368 5176 17374 5228
rect 19334 5216 19340 5228
rect 17972 5188 19340 5216
rect 17972 5148 18000 5188
rect 19334 5176 19340 5188
rect 19392 5176 19398 5228
rect 19886 5176 19892 5228
rect 19944 5216 19950 5228
rect 20165 5219 20223 5225
rect 20165 5216 20177 5219
rect 19944 5188 20177 5216
rect 19944 5176 19950 5188
rect 20165 5185 20177 5188
rect 20211 5185 20223 5219
rect 21560 5216 21588 5256
rect 22370 5244 22376 5256
rect 22428 5244 22434 5296
rect 23474 5244 23480 5296
rect 23532 5284 23538 5296
rect 24182 5287 24240 5293
rect 24182 5284 24194 5287
rect 23532 5256 24194 5284
rect 23532 5244 23538 5256
rect 24182 5253 24194 5256
rect 24228 5253 24240 5287
rect 24182 5247 24240 5253
rect 25682 5244 25688 5296
rect 25740 5284 25746 5296
rect 26145 5287 26203 5293
rect 26145 5284 26157 5287
rect 25740 5256 26157 5284
rect 25740 5244 25746 5256
rect 26145 5253 26157 5256
rect 26191 5253 26203 5287
rect 30374 5284 30380 5296
rect 26145 5247 26203 5253
rect 26988 5256 30380 5284
rect 22261 5219 22319 5225
rect 22261 5216 22273 5219
rect 20165 5179 20223 5185
rect 21100 5188 21588 5216
rect 21621 5188 22273 5216
rect 18138 5148 18144 5160
rect 16592 5120 18000 5148
rect 18099 5120 18144 5148
rect 18138 5108 18144 5120
rect 18196 5108 18202 5160
rect 20438 5148 20444 5160
rect 20399 5120 20444 5148
rect 20438 5108 20444 5120
rect 20496 5108 20502 5160
rect 15746 5080 15752 5092
rect 15304 5052 15752 5080
rect 15746 5040 15752 5052
rect 15804 5040 15810 5092
rect 16669 5083 16727 5089
rect 16669 5049 16681 5083
rect 16715 5080 16727 5083
rect 16715 5052 18196 5080
rect 16715 5049 16727 5052
rect 16669 5043 16727 5049
rect 15562 5012 15568 5024
rect 12728 4984 15568 5012
rect 15562 4972 15568 4984
rect 15620 4972 15626 5024
rect 16942 4972 16948 5024
rect 17000 5012 17006 5024
rect 17313 5015 17371 5021
rect 17313 5012 17325 5015
rect 17000 4984 17325 5012
rect 17000 4972 17006 4984
rect 17313 4981 17325 4984
rect 17359 4981 17371 5015
rect 18168 5012 18196 5052
rect 18782 5012 18788 5024
rect 18168 4984 18788 5012
rect 17313 4975 17371 4981
rect 18782 4972 18788 4984
rect 18840 5012 18846 5024
rect 19521 5015 19579 5021
rect 19521 5012 19533 5015
rect 18840 4984 19533 5012
rect 18840 4972 18846 4984
rect 19521 4981 19533 4984
rect 19567 4981 19579 5015
rect 19978 5012 19984 5024
rect 19939 4984 19984 5012
rect 19521 4975 19579 4981
rect 19978 4972 19984 4984
rect 20036 4972 20042 5024
rect 20254 4972 20260 5024
rect 20312 5012 20318 5024
rect 21100 5021 21128 5188
rect 21266 5108 21272 5160
rect 21324 5148 21330 5160
rect 21621 5148 21649 5188
rect 22261 5185 22273 5188
rect 22307 5185 22319 5219
rect 22261 5179 22319 5185
rect 23937 5219 23995 5225
rect 23937 5185 23949 5219
rect 23983 5216 23995 5219
rect 24026 5216 24032 5228
rect 23983 5188 24032 5216
rect 23983 5185 23995 5188
rect 23937 5179 23995 5185
rect 24026 5176 24032 5188
rect 24084 5176 24090 5228
rect 25774 5216 25780 5228
rect 25735 5188 25780 5216
rect 25774 5176 25780 5188
rect 25832 5176 25838 5228
rect 25870 5219 25928 5225
rect 25870 5185 25882 5219
rect 25916 5185 25928 5219
rect 25870 5179 25928 5185
rect 26053 5219 26111 5225
rect 26053 5185 26065 5219
rect 26099 5185 26111 5219
rect 26053 5179 26111 5185
rect 26283 5219 26341 5225
rect 26283 5185 26295 5219
rect 26329 5216 26341 5219
rect 26694 5216 26700 5228
rect 26329 5188 26700 5216
rect 26329 5185 26341 5188
rect 26283 5179 26341 5185
rect 22002 5148 22008 5160
rect 21324 5120 21649 5148
rect 21963 5120 22008 5148
rect 21324 5108 21330 5120
rect 22002 5108 22008 5120
rect 22060 5108 22066 5160
rect 25884 5148 25912 5179
rect 25332 5120 25912 5148
rect 26068 5148 26096 5179
rect 26694 5176 26700 5188
rect 26752 5176 26758 5228
rect 26988 5225 27016 5256
rect 30374 5244 30380 5256
rect 30432 5244 30438 5296
rect 30190 5225 30196 5228
rect 26973 5219 27031 5225
rect 26973 5185 26985 5219
rect 27019 5185 27031 5219
rect 26973 5179 27031 5185
rect 27976 5219 28034 5225
rect 27976 5185 27988 5219
rect 28022 5216 28034 5219
rect 30184 5216 30196 5225
rect 28022 5188 29500 5216
rect 30151 5188 30196 5216
rect 28022 5185 28034 5188
rect 27976 5179 28034 5185
rect 26068 5120 26556 5148
rect 23290 5040 23296 5092
rect 23348 5080 23354 5092
rect 23385 5083 23443 5089
rect 23385 5080 23397 5083
rect 23348 5052 23397 5080
rect 23348 5040 23354 5052
rect 23385 5049 23397 5052
rect 23431 5049 23443 5083
rect 23385 5043 23443 5049
rect 20349 5015 20407 5021
rect 20349 5012 20361 5015
rect 20312 4984 20361 5012
rect 20312 4972 20318 4984
rect 20349 4981 20361 4984
rect 20395 4981 20407 5015
rect 20349 4975 20407 4981
rect 21085 5015 21143 5021
rect 21085 4981 21097 5015
rect 21131 4981 21143 5015
rect 21085 4975 21143 4981
rect 21269 5015 21327 5021
rect 21269 4981 21281 5015
rect 21315 5012 21327 5015
rect 22002 5012 22008 5024
rect 21315 4984 22008 5012
rect 21315 4981 21327 4984
rect 21269 4975 21327 4981
rect 22002 4972 22008 4984
rect 22060 4972 22066 5024
rect 22186 4972 22192 5024
rect 22244 5012 22250 5024
rect 23308 5012 23336 5040
rect 22244 4984 23336 5012
rect 22244 4972 22250 4984
rect 24946 4972 24952 5024
rect 25004 5012 25010 5024
rect 25332 5021 25360 5120
rect 26418 5080 26424 5092
rect 26379 5052 26424 5080
rect 26418 5040 26424 5052
rect 26476 5040 26482 5092
rect 26528 5080 26556 5120
rect 27614 5108 27620 5160
rect 27672 5148 27678 5160
rect 27709 5151 27767 5157
rect 27709 5148 27721 5151
rect 27672 5120 27721 5148
rect 27672 5108 27678 5120
rect 27709 5117 27721 5120
rect 27755 5117 27767 5151
rect 27709 5111 27767 5117
rect 27246 5080 27252 5092
rect 26528 5052 27252 5080
rect 27246 5040 27252 5052
rect 27304 5040 27310 5092
rect 25317 5015 25375 5021
rect 25317 5012 25329 5015
rect 25004 4984 25329 5012
rect 25004 4972 25010 4984
rect 25317 4981 25329 4984
rect 25363 4981 25375 5015
rect 25317 4975 25375 4981
rect 25406 4972 25412 5024
rect 25464 5012 25470 5024
rect 28626 5012 28632 5024
rect 25464 4984 28632 5012
rect 25464 4972 25470 4984
rect 28626 4972 28632 4984
rect 28684 4972 28690 5024
rect 29086 5012 29092 5024
rect 29047 4984 29092 5012
rect 29086 4972 29092 4984
rect 29144 4972 29150 5024
rect 29472 5012 29500 5188
rect 30184 5179 30196 5188
rect 30190 5176 30196 5179
rect 30248 5176 30254 5228
rect 29546 5108 29552 5160
rect 29604 5148 29610 5160
rect 29914 5148 29920 5160
rect 29604 5120 29920 5148
rect 29604 5108 29610 5120
rect 29914 5108 29920 5120
rect 29972 5108 29978 5160
rect 30650 5012 30656 5024
rect 29472 4984 30656 5012
rect 30650 4972 30656 4984
rect 30708 4972 30714 5024
rect 31294 5012 31300 5024
rect 31255 4984 31300 5012
rect 31294 4972 31300 4984
rect 31352 4972 31358 5024
rect 1104 4922 32016 4944
rect 1104 4870 2136 4922
rect 2188 4870 12440 4922
rect 12492 4870 22744 4922
rect 22796 4870 32016 4922
rect 1104 4848 32016 4870
rect 1578 4768 1584 4820
rect 1636 4808 1642 4820
rect 2777 4811 2835 4817
rect 2777 4808 2789 4811
rect 1636 4780 2789 4808
rect 1636 4768 1642 4780
rect 1394 4672 1400 4684
rect 1355 4644 1400 4672
rect 1394 4632 1400 4644
rect 1452 4632 1458 4684
rect 1670 4613 1676 4616
rect 1664 4604 1676 4613
rect 1631 4576 1676 4604
rect 1664 4567 1676 4576
rect 1670 4564 1676 4567
rect 1728 4564 1734 4616
rect 2516 4604 2544 4780
rect 2777 4777 2789 4780
rect 2823 4777 2835 4811
rect 2777 4771 2835 4777
rect 5258 4768 5264 4820
rect 5316 4808 5322 4820
rect 7558 4808 7564 4820
rect 5316 4780 7564 4808
rect 5316 4768 5322 4780
rect 7558 4768 7564 4780
rect 7616 4768 7622 4820
rect 7926 4808 7932 4820
rect 7887 4780 7932 4808
rect 7926 4768 7932 4780
rect 7984 4768 7990 4820
rect 9674 4768 9680 4820
rect 9732 4808 9738 4820
rect 14734 4808 14740 4820
rect 9732 4780 14740 4808
rect 9732 4768 9738 4780
rect 14734 4768 14740 4780
rect 14792 4768 14798 4820
rect 15010 4768 15016 4820
rect 15068 4808 15074 4820
rect 18046 4808 18052 4820
rect 15068 4780 18052 4808
rect 15068 4768 15074 4780
rect 18046 4768 18052 4780
rect 18104 4768 18110 4820
rect 18141 4811 18199 4817
rect 18141 4777 18153 4811
rect 18187 4808 18199 4811
rect 19521 4811 19579 4817
rect 19521 4808 19533 4811
rect 18187 4780 19533 4808
rect 18187 4777 18199 4780
rect 18141 4771 18199 4777
rect 19521 4777 19533 4780
rect 19567 4777 19579 4811
rect 19521 4771 19579 4777
rect 20809 4811 20867 4817
rect 20809 4777 20821 4811
rect 20855 4808 20867 4811
rect 21266 4808 21272 4820
rect 20855 4780 21272 4808
rect 20855 4777 20867 4780
rect 20809 4771 20867 4777
rect 21266 4768 21272 4780
rect 21324 4768 21330 4820
rect 24596 4780 28212 4808
rect 6178 4700 6184 4752
rect 6236 4740 6242 4752
rect 6638 4740 6644 4752
rect 6236 4712 6644 4740
rect 6236 4700 6242 4712
rect 6638 4700 6644 4712
rect 6696 4700 6702 4752
rect 7650 4700 7656 4752
rect 7708 4740 7714 4752
rect 7745 4743 7803 4749
rect 7745 4740 7757 4743
rect 7708 4712 7757 4740
rect 7708 4700 7714 4712
rect 7745 4709 7757 4712
rect 7791 4740 7803 4743
rect 8018 4740 8024 4752
rect 7791 4712 8024 4740
rect 7791 4709 7803 4712
rect 7745 4703 7803 4709
rect 8018 4700 8024 4712
rect 8076 4700 8082 4752
rect 12618 4700 12624 4752
rect 12676 4740 12682 4752
rect 12897 4743 12955 4749
rect 12897 4740 12909 4743
rect 12676 4712 12909 4740
rect 12676 4700 12682 4712
rect 12897 4709 12909 4712
rect 12943 4740 12955 4743
rect 15838 4740 15844 4752
rect 12943 4712 15844 4740
rect 12943 4709 12955 4712
rect 12897 4703 12955 4709
rect 2590 4632 2596 4684
rect 2648 4672 2654 4684
rect 9306 4672 9312 4684
rect 2648 4644 3818 4672
rect 6196 4644 9312 4672
rect 2648 4632 2654 4644
rect 2682 4604 2688 4616
rect 2516 4576 2688 4604
rect 2682 4564 2688 4576
rect 2740 4604 2746 4616
rect 6196 4613 6224 4644
rect 9306 4632 9312 4644
rect 9364 4632 9370 4684
rect 11330 4632 11336 4684
rect 11388 4672 11394 4684
rect 11517 4675 11575 4681
rect 11517 4672 11529 4675
rect 11388 4644 11529 4672
rect 11388 4632 11394 4644
rect 11517 4641 11529 4644
rect 11563 4641 11575 4675
rect 11517 4635 11575 4641
rect 13449 4675 13507 4681
rect 13449 4641 13461 4675
rect 13495 4672 13507 4675
rect 13633 4675 13691 4681
rect 13633 4672 13645 4675
rect 13495 4644 13645 4672
rect 13495 4641 13507 4644
rect 13449 4635 13507 4641
rect 13633 4641 13645 4644
rect 13679 4641 13691 4675
rect 14366 4672 14372 4684
rect 14327 4644 14372 4672
rect 13633 4635 13691 4641
rect 14366 4632 14372 4644
rect 14424 4632 14430 4684
rect 15102 4672 15108 4684
rect 14568 4644 15108 4672
rect 4341 4607 4399 4613
rect 4341 4604 4353 4607
rect 2740 4576 4353 4604
rect 2740 4564 2746 4576
rect 4341 4573 4353 4576
rect 4387 4573 4399 4607
rect 4341 4567 4399 4573
rect 6181 4607 6239 4613
rect 6181 4573 6193 4607
rect 6227 4573 6239 4607
rect 6181 4567 6239 4573
rect 6457 4607 6515 4613
rect 6457 4573 6469 4607
rect 6503 4573 6515 4607
rect 6638 4604 6644 4616
rect 6599 4576 6644 4604
rect 6457 4567 6515 4573
rect 0 4536 800 4550
rect 937 4539 995 4545
rect 937 4536 949 4539
rect 0 4508 949 4536
rect 0 4494 800 4508
rect 937 4505 949 4508
rect 983 4505 995 4539
rect 937 4499 995 4505
rect 3786 4496 3792 4548
rect 3844 4536 3850 4548
rect 3973 4539 4031 4545
rect 3973 4536 3985 4539
rect 3844 4508 3985 4536
rect 3844 4496 3850 4508
rect 3973 4505 3985 4508
rect 4019 4505 4031 4539
rect 3973 4499 4031 4505
rect 4249 4539 4307 4545
rect 4249 4505 4261 4539
rect 4295 4505 4307 4539
rect 4706 4536 4712 4548
rect 4667 4508 4712 4536
rect 4249 4499 4307 4505
rect 3234 4428 3240 4480
rect 3292 4468 3298 4480
rect 4264 4468 4292 4499
rect 4706 4496 4712 4508
rect 4764 4496 4770 4548
rect 6472 4536 6500 4567
rect 6638 4564 6644 4576
rect 6696 4564 6702 4616
rect 9493 4607 9551 4613
rect 9493 4573 9505 4607
rect 9539 4604 9551 4607
rect 9582 4604 9588 4616
rect 9539 4576 9588 4604
rect 9539 4573 9551 4576
rect 9493 4567 9551 4573
rect 9582 4564 9588 4576
rect 9640 4604 9646 4616
rect 11348 4604 11376 4632
rect 9640 4576 11376 4604
rect 11784 4607 11842 4613
rect 9640 4564 9646 4576
rect 11784 4573 11796 4607
rect 11830 4604 11842 4607
rect 12158 4604 12164 4616
rect 11830 4576 12164 4604
rect 11830 4573 11842 4576
rect 11784 4567 11842 4573
rect 12158 4564 12164 4576
rect 12216 4564 12222 4616
rect 13357 4607 13415 4613
rect 13357 4573 13369 4607
rect 13403 4573 13415 4607
rect 13538 4604 13544 4616
rect 13499 4576 13544 4604
rect 13357 4567 13415 4573
rect 6730 4536 6736 4548
rect 6472 4508 6736 4536
rect 6730 4496 6736 4508
rect 6788 4496 6794 4548
rect 7466 4536 7472 4548
rect 7427 4508 7472 4536
rect 7466 4496 7472 4508
rect 7524 4496 7530 4548
rect 9760 4539 9818 4545
rect 9760 4505 9772 4539
rect 9806 4536 9818 4539
rect 10318 4536 10324 4548
rect 9806 4508 10324 4536
rect 9806 4505 9818 4508
rect 9760 4499 9818 4505
rect 10318 4496 10324 4508
rect 10376 4496 10382 4548
rect 13372 4536 13400 4567
rect 13538 4564 13544 4576
rect 13596 4564 13602 4616
rect 14090 4604 14096 4616
rect 14003 4576 14096 4604
rect 14090 4564 14096 4576
rect 14148 4604 14154 4616
rect 14568 4604 14596 4644
rect 15102 4632 15108 4644
rect 15160 4632 15166 4684
rect 14148 4576 14596 4604
rect 14148 4564 14154 4576
rect 15010 4564 15016 4616
rect 15068 4604 15074 4616
rect 15672 4613 15700 4712
rect 15838 4700 15844 4712
rect 15896 4700 15902 4752
rect 15933 4743 15991 4749
rect 15933 4709 15945 4743
rect 15979 4740 15991 4743
rect 16022 4740 16028 4752
rect 15979 4712 16028 4740
rect 15979 4709 15991 4712
rect 15933 4703 15991 4709
rect 16022 4700 16028 4712
rect 16080 4700 16086 4752
rect 16298 4700 16304 4752
rect 16356 4740 16362 4752
rect 17310 4740 17316 4752
rect 16356 4712 17316 4740
rect 16356 4700 16362 4712
rect 17310 4700 17316 4712
rect 17368 4740 17374 4752
rect 19245 4743 19303 4749
rect 19245 4740 19257 4743
rect 17368 4712 19257 4740
rect 17368 4700 17374 4712
rect 19245 4709 19257 4712
rect 19291 4709 19303 4743
rect 19245 4703 19303 4709
rect 22094 4700 22100 4752
rect 22152 4740 22158 4752
rect 23106 4740 23112 4752
rect 22152 4712 23112 4740
rect 22152 4700 22158 4712
rect 23106 4700 23112 4712
rect 23164 4740 23170 4752
rect 23164 4712 23520 4740
rect 23164 4700 23170 4712
rect 16390 4632 16396 4684
rect 16448 4672 16454 4684
rect 18141 4675 18199 4681
rect 18141 4672 18153 4675
rect 16448 4644 18153 4672
rect 16448 4632 16454 4644
rect 18141 4641 18153 4644
rect 18187 4641 18199 4675
rect 18141 4635 18199 4641
rect 18233 4675 18291 4681
rect 18233 4641 18245 4675
rect 18279 4672 18291 4675
rect 18322 4672 18328 4684
rect 18279 4644 18328 4672
rect 18279 4641 18291 4644
rect 18233 4635 18291 4641
rect 18322 4632 18328 4644
rect 18380 4632 18386 4684
rect 18598 4672 18604 4684
rect 18559 4644 18604 4672
rect 18598 4632 18604 4644
rect 18656 4672 18662 4684
rect 20254 4672 20260 4684
rect 18656 4644 20260 4672
rect 18656 4632 18662 4644
rect 20254 4632 20260 4644
rect 20312 4632 20318 4684
rect 20349 4675 20407 4681
rect 20349 4641 20361 4675
rect 20395 4672 20407 4675
rect 20622 4672 20628 4684
rect 20395 4644 20628 4672
rect 20395 4641 20407 4644
rect 20349 4635 20407 4641
rect 20622 4632 20628 4644
rect 20680 4632 20686 4684
rect 21269 4675 21327 4681
rect 21269 4641 21281 4675
rect 21315 4672 21327 4675
rect 23198 4672 23204 4684
rect 21315 4644 23204 4672
rect 21315 4641 21327 4644
rect 21269 4635 21327 4641
rect 23198 4632 23204 4644
rect 23256 4632 23262 4684
rect 23492 4681 23520 4712
rect 23477 4675 23535 4681
rect 23477 4641 23489 4675
rect 23523 4672 23535 4675
rect 23566 4672 23572 4684
rect 23523 4644 23572 4672
rect 23523 4641 23535 4644
rect 23477 4635 23535 4641
rect 23566 4632 23572 4644
rect 23624 4632 23630 4684
rect 23842 4632 23848 4684
rect 23900 4672 23906 4684
rect 24596 4681 24624 4780
rect 26234 4700 26240 4752
rect 26292 4740 26298 4752
rect 26292 4712 26556 4740
rect 26292 4700 26298 4712
rect 24581 4675 24639 4681
rect 24581 4672 24593 4675
rect 23900 4644 24593 4672
rect 23900 4632 23906 4644
rect 24581 4641 24593 4644
rect 24627 4641 24639 4675
rect 24854 4672 24860 4684
rect 24815 4644 24860 4672
rect 24581 4635 24639 4641
rect 24854 4632 24860 4644
rect 24912 4632 24918 4684
rect 26528 4681 26556 4712
rect 26513 4675 26571 4681
rect 26513 4641 26525 4675
rect 26559 4641 26571 4675
rect 27982 4672 27988 4684
rect 26513 4635 26571 4641
rect 27632 4644 27988 4672
rect 15401 4607 15459 4613
rect 15401 4604 15413 4607
rect 15068 4576 15413 4604
rect 15068 4564 15074 4576
rect 15401 4573 15413 4576
rect 15447 4573 15459 4607
rect 15401 4567 15459 4573
rect 15657 4607 15715 4613
rect 15657 4573 15669 4607
rect 15703 4573 15715 4607
rect 15657 4567 15715 4573
rect 15795 4607 15853 4613
rect 15795 4573 15807 4607
rect 15841 4604 15853 4607
rect 16850 4604 16856 4616
rect 15841 4576 16856 4604
rect 15841 4573 15853 4576
rect 15795 4567 15853 4573
rect 16850 4564 16856 4576
rect 16908 4564 16914 4616
rect 16945 4607 17003 4613
rect 16945 4573 16957 4607
rect 16991 4573 17003 4607
rect 16945 4567 17003 4573
rect 17221 4607 17279 4613
rect 17221 4573 17233 4607
rect 17267 4604 17279 4607
rect 17310 4604 17316 4616
rect 17267 4576 17316 4604
rect 17267 4573 17279 4576
rect 17221 4567 17279 4573
rect 15194 4536 15200 4548
rect 13372 4508 15200 4536
rect 13556 4480 13584 4508
rect 15194 4496 15200 4508
rect 15252 4496 15258 4548
rect 15562 4536 15568 4548
rect 15523 4508 15568 4536
rect 15562 4496 15568 4508
rect 15620 4496 15626 4548
rect 15930 4496 15936 4548
rect 15988 4536 15994 4548
rect 16960 4536 16988 4567
rect 17310 4564 17316 4576
rect 17368 4564 17374 4616
rect 18477 4607 18535 4613
rect 18477 4573 18489 4607
rect 18523 4604 18535 4607
rect 18689 4607 18747 4613
rect 18523 4573 18552 4604
rect 18477 4567 18552 4573
rect 18689 4573 18701 4607
rect 18735 4573 18747 4607
rect 18689 4567 18747 4573
rect 18877 4607 18935 4613
rect 18877 4573 18889 4607
rect 18923 4604 18935 4607
rect 19245 4607 19303 4613
rect 19245 4604 19257 4607
rect 18923 4576 19257 4604
rect 18923 4573 18935 4576
rect 18877 4567 18935 4573
rect 19245 4573 19257 4576
rect 19291 4573 19303 4607
rect 19245 4567 19303 4573
rect 19429 4607 19487 4613
rect 19429 4573 19441 4607
rect 19475 4604 19487 4607
rect 19521 4607 19579 4613
rect 19521 4604 19533 4607
rect 19475 4576 19533 4604
rect 19475 4573 19487 4576
rect 19429 4567 19487 4573
rect 19521 4573 19533 4576
rect 19567 4573 19579 4607
rect 20070 4604 20076 4616
rect 20031 4576 20076 4604
rect 19521 4567 19579 4573
rect 15988 4508 16988 4536
rect 15988 4496 15994 4508
rect 17126 4496 17132 4548
rect 17184 4536 17190 4548
rect 17678 4536 17684 4548
rect 17184 4508 17684 4536
rect 17184 4496 17190 4508
rect 17678 4496 17684 4508
rect 17736 4496 17742 4548
rect 18322 4496 18328 4548
rect 18380 4536 18386 4548
rect 18524 4536 18552 4567
rect 18380 4508 18552 4536
rect 18708 4536 18736 4567
rect 20070 4564 20076 4576
rect 20128 4564 20134 4616
rect 20990 4604 20996 4616
rect 20951 4576 20996 4604
rect 20990 4564 20996 4576
rect 21048 4564 21054 4616
rect 21174 4604 21180 4616
rect 21135 4576 21180 4604
rect 21174 4564 21180 4576
rect 21232 4564 21238 4616
rect 21726 4604 21732 4616
rect 21687 4576 21732 4604
rect 21726 4564 21732 4576
rect 21784 4604 21790 4616
rect 21784 4576 22094 4604
rect 21784 4564 21790 4576
rect 19150 4536 19156 4548
rect 18708 4508 19156 4536
rect 18380 4496 18386 4508
rect 19150 4496 19156 4508
rect 19208 4536 19214 4548
rect 20622 4536 20628 4548
rect 19208 4508 20628 4536
rect 19208 4496 19214 4508
rect 20622 4496 20628 4508
rect 20680 4496 20686 4548
rect 22066 4536 22094 4576
rect 22554 4564 22560 4616
rect 22612 4604 22618 4616
rect 26237 4607 26295 4613
rect 26237 4604 26249 4607
rect 22612 4576 26249 4604
rect 22612 4564 22618 4576
rect 26237 4573 26249 4576
rect 26283 4604 26295 4607
rect 27632 4604 27660 4644
rect 27982 4632 27988 4644
rect 28040 4632 28046 4684
rect 28184 4681 28212 4780
rect 28169 4675 28227 4681
rect 28169 4641 28181 4675
rect 28215 4672 28227 4675
rect 29178 4672 29184 4684
rect 28215 4644 29184 4672
rect 28215 4641 28227 4644
rect 28169 4635 28227 4641
rect 29178 4632 29184 4644
rect 29236 4632 29242 4684
rect 29546 4672 29552 4684
rect 29507 4644 29552 4672
rect 29546 4632 29552 4644
rect 29604 4632 29610 4684
rect 26283 4576 27660 4604
rect 27709 4607 27767 4613
rect 26283 4573 26295 4576
rect 26237 4567 26295 4573
rect 27709 4573 27721 4607
rect 27755 4604 27767 4607
rect 28074 4604 28080 4616
rect 27755 4576 28080 4604
rect 27755 4573 27767 4576
rect 27709 4567 27767 4573
rect 28074 4564 28080 4576
rect 28132 4564 28138 4616
rect 28445 4607 28503 4613
rect 28445 4573 28457 4607
rect 28491 4604 28503 4607
rect 28534 4604 28540 4616
rect 28491 4576 28540 4604
rect 28491 4573 28503 4576
rect 28445 4567 28503 4573
rect 28534 4564 28540 4576
rect 28592 4564 28598 4616
rect 26970 4536 26976 4548
rect 22066 4508 26976 4536
rect 26970 4496 26976 4508
rect 27028 4536 27034 4548
rect 27798 4536 27804 4548
rect 27028 4508 27804 4536
rect 27028 4496 27034 4508
rect 27798 4496 27804 4508
rect 27856 4496 27862 4548
rect 29362 4496 29368 4548
rect 29420 4536 29426 4548
rect 29794 4539 29852 4545
rect 29794 4536 29806 4539
rect 29420 4508 29806 4536
rect 29420 4496 29426 4508
rect 29794 4505 29806 4508
rect 29840 4505 29852 4539
rect 32320 4536 33120 4550
rect 29794 4499 29852 4505
rect 29932 4508 33120 4536
rect 5074 4468 5080 4480
rect 3292 4440 4292 4468
rect 5035 4440 5080 4468
rect 3292 4428 3298 4440
rect 5074 4428 5080 4440
rect 5132 4428 5138 4480
rect 5258 4468 5264 4480
rect 5219 4440 5264 4468
rect 5258 4428 5264 4440
rect 5316 4428 5322 4480
rect 5997 4471 6055 4477
rect 5997 4437 6009 4471
rect 6043 4468 6055 4471
rect 6362 4468 6368 4480
rect 6043 4440 6368 4468
rect 6043 4437 6055 4440
rect 5997 4431 6055 4437
rect 6362 4428 6368 4440
rect 6420 4428 6426 4480
rect 9490 4428 9496 4480
rect 9548 4468 9554 4480
rect 10873 4471 10931 4477
rect 10873 4468 10885 4471
rect 9548 4440 10885 4468
rect 9548 4428 9554 4440
rect 10873 4437 10885 4440
rect 10919 4437 10931 4471
rect 10873 4431 10931 4437
rect 13538 4428 13544 4480
rect 13596 4428 13602 4480
rect 13633 4471 13691 4477
rect 13633 4437 13645 4471
rect 13679 4468 13691 4471
rect 15746 4468 15752 4480
rect 13679 4440 15752 4468
rect 13679 4437 13691 4440
rect 13633 4431 13691 4437
rect 15746 4428 15752 4440
rect 15804 4468 15810 4480
rect 18877 4471 18935 4477
rect 18877 4468 18889 4471
rect 15804 4440 18889 4468
rect 15804 4428 15810 4440
rect 18877 4437 18889 4440
rect 18923 4437 18935 4471
rect 18877 4431 18935 4437
rect 19889 4471 19947 4477
rect 19889 4437 19901 4471
rect 19935 4468 19947 4471
rect 20162 4468 20168 4480
rect 19935 4440 20168 4468
rect 19935 4437 19947 4440
rect 19889 4431 19947 4437
rect 20162 4428 20168 4440
rect 20220 4428 20226 4480
rect 27525 4471 27583 4477
rect 27525 4437 27537 4471
rect 27571 4468 27583 4471
rect 28258 4468 28264 4480
rect 27571 4440 28264 4468
rect 27571 4437 27583 4440
rect 27525 4431 27583 4437
rect 28258 4428 28264 4440
rect 28316 4428 28322 4480
rect 28350 4428 28356 4480
rect 28408 4468 28414 4480
rect 29932 4468 29960 4508
rect 32320 4494 33120 4508
rect 28408 4440 29960 4468
rect 28408 4428 28414 4440
rect 30006 4428 30012 4480
rect 30064 4468 30070 4480
rect 30929 4471 30987 4477
rect 30929 4468 30941 4471
rect 30064 4440 30941 4468
rect 30064 4428 30070 4440
rect 30929 4437 30941 4440
rect 30975 4468 30987 4471
rect 31110 4468 31116 4480
rect 30975 4440 31116 4468
rect 30975 4437 30987 4440
rect 30929 4431 30987 4437
rect 31110 4428 31116 4440
rect 31168 4428 31174 4480
rect 1104 4378 32016 4400
rect 1104 4326 7288 4378
rect 7340 4326 17592 4378
rect 17644 4326 27896 4378
rect 27948 4326 32016 4378
rect 1104 4304 32016 4326
rect 1949 4267 2007 4273
rect 1949 4233 1961 4267
rect 1995 4264 2007 4267
rect 2038 4264 2044 4276
rect 1995 4236 2044 4264
rect 1995 4233 2007 4236
rect 1949 4227 2007 4233
rect 2038 4224 2044 4236
rect 2096 4224 2102 4276
rect 3053 4267 3111 4273
rect 3053 4233 3065 4267
rect 3099 4264 3111 4267
rect 4706 4264 4712 4276
rect 3099 4236 4712 4264
rect 3099 4233 3111 4236
rect 3053 4227 3111 4233
rect 4706 4224 4712 4236
rect 4764 4224 4770 4276
rect 4982 4224 4988 4276
rect 5040 4264 5046 4276
rect 6733 4267 6791 4273
rect 6733 4264 6745 4267
rect 5040 4236 6745 4264
rect 5040 4224 5046 4236
rect 6733 4233 6745 4236
rect 6779 4233 6791 4267
rect 6733 4227 6791 4233
rect 7466 4224 7472 4276
rect 7524 4264 7530 4276
rect 9950 4264 9956 4276
rect 7524 4236 9956 4264
rect 7524 4224 7530 4236
rect 9950 4224 9956 4236
rect 10008 4224 10014 4276
rect 10318 4264 10324 4276
rect 10279 4236 10324 4264
rect 10318 4224 10324 4236
rect 10376 4224 10382 4276
rect 13998 4264 14004 4276
rect 10428 4236 14004 4264
rect 3970 4196 3976 4208
rect 3436 4168 3976 4196
rect 2133 4131 2191 4137
rect 2133 4097 2145 4131
rect 2179 4128 2191 4131
rect 2222 4128 2228 4140
rect 2179 4100 2228 4128
rect 2179 4097 2191 4100
rect 2133 4091 2191 4097
rect 2222 4088 2228 4100
rect 2280 4088 2286 4140
rect 2406 4128 2412 4140
rect 2367 4100 2412 4128
rect 2406 4088 2412 4100
rect 2464 4088 2470 4140
rect 2593 4131 2651 4137
rect 2593 4097 2605 4131
rect 2639 4128 2651 4131
rect 2682 4128 2688 4140
rect 2639 4100 2688 4128
rect 2639 4097 2651 4100
rect 2593 4091 2651 4097
rect 2682 4088 2688 4100
rect 2740 4088 2746 4140
rect 2866 4088 2872 4140
rect 2924 4128 2930 4140
rect 3436 4137 3464 4168
rect 3970 4156 3976 4168
rect 4028 4156 4034 4208
rect 5258 4156 5264 4208
rect 5316 4196 5322 4208
rect 10428 4196 10456 4236
rect 13998 4224 14004 4236
rect 14056 4224 14062 4276
rect 14274 4224 14280 4276
rect 14332 4264 14338 4276
rect 15105 4267 15163 4273
rect 15105 4264 15117 4267
rect 14332 4236 15117 4264
rect 14332 4224 14338 4236
rect 15105 4233 15117 4236
rect 15151 4233 15163 4267
rect 15105 4227 15163 4233
rect 15194 4224 15200 4276
rect 15252 4264 15258 4276
rect 15930 4264 15936 4276
rect 15252 4236 15936 4264
rect 15252 4224 15258 4236
rect 15930 4224 15936 4236
rect 15988 4224 15994 4276
rect 16482 4224 16488 4276
rect 16540 4264 16546 4276
rect 17589 4267 17647 4273
rect 16540 4236 17453 4264
rect 16540 4224 16546 4236
rect 11882 4196 11888 4208
rect 5316 4168 10456 4196
rect 11843 4168 11888 4196
rect 5316 4156 5322 4168
rect 11882 4156 11888 4168
rect 11940 4156 11946 4208
rect 13078 4156 13084 4208
rect 13136 4196 13142 4208
rect 15010 4196 15016 4208
rect 13136 4168 15016 4196
rect 13136 4156 13142 4168
rect 3421 4131 3479 4137
rect 3421 4128 3433 4131
rect 2924 4100 3433 4128
rect 2924 4088 2930 4100
rect 3421 4097 3433 4100
rect 3467 4097 3479 4131
rect 3421 4091 3479 4097
rect 3513 4131 3571 4137
rect 3513 4097 3525 4131
rect 3559 4128 3571 4131
rect 3786 4128 3792 4140
rect 3559 4100 3792 4128
rect 3559 4097 3571 4100
rect 3513 4091 3571 4097
rect 3786 4088 3792 4100
rect 3844 4088 3850 4140
rect 4246 4128 4252 4140
rect 4207 4100 4252 4128
rect 4246 4088 4252 4100
rect 4304 4088 4310 4140
rect 4516 4131 4574 4137
rect 4516 4097 4528 4131
rect 4562 4128 4574 4131
rect 5442 4128 5448 4140
rect 4562 4100 5448 4128
rect 4562 4097 4574 4100
rect 4516 4091 4574 4097
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 6825 4131 6883 4137
rect 6825 4097 6837 4131
rect 6871 4128 6883 4131
rect 7374 4128 7380 4140
rect 6871 4100 7380 4128
rect 6871 4097 6883 4100
rect 6825 4091 6883 4097
rect 7374 4088 7380 4100
rect 7432 4088 7438 4140
rect 7650 4088 7656 4140
rect 7708 4128 7714 4140
rect 8570 4128 8576 4140
rect 7708 4100 8576 4128
rect 7708 4088 7714 4100
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 9306 4088 9312 4140
rect 9364 4128 9370 4140
rect 9401 4131 9459 4137
rect 9401 4128 9413 4131
rect 9364 4100 9413 4128
rect 9364 4088 9370 4100
rect 9401 4097 9413 4100
rect 9447 4097 9459 4131
rect 9401 4091 9459 4097
rect 9677 4131 9735 4137
rect 9677 4097 9689 4131
rect 9723 4097 9735 4131
rect 9677 4091 9735 4097
rect 9861 4131 9919 4137
rect 9861 4097 9873 4131
rect 9907 4128 9919 4131
rect 9950 4128 9956 4140
rect 9907 4100 9956 4128
rect 9907 4097 9919 4100
rect 9861 4091 9919 4097
rect 3694 4020 3700 4072
rect 3752 4060 3758 4072
rect 7009 4063 7067 4069
rect 3752 4032 3797 4060
rect 3752 4020 3758 4032
rect 7009 4029 7021 4063
rect 7055 4060 7067 4063
rect 7098 4060 7104 4072
rect 7055 4032 7104 4060
rect 7055 4029 7067 4032
rect 7009 4023 7067 4029
rect 7098 4020 7104 4032
rect 7156 4060 7162 4072
rect 7561 4063 7619 4069
rect 7561 4060 7573 4063
rect 7156 4032 7573 4060
rect 7156 4020 7162 4032
rect 7561 4029 7573 4032
rect 7607 4029 7619 4063
rect 8757 4063 8815 4069
rect 8757 4060 8769 4063
rect 7561 4023 7619 4029
rect 7760 4032 8769 4060
rect 2406 3952 2412 4004
rect 2464 3992 2470 4004
rect 3510 3992 3516 4004
rect 2464 3964 3516 3992
rect 2464 3952 2470 3964
rect 3510 3952 3516 3964
rect 3568 3952 3574 4004
rect 5629 3995 5687 4001
rect 5629 3961 5641 3995
rect 5675 3992 5687 3995
rect 5810 3992 5816 4004
rect 5675 3964 5816 3992
rect 5675 3961 5687 3964
rect 5629 3955 5687 3961
rect 5810 3952 5816 3964
rect 5868 3952 5874 4004
rect 6730 3952 6736 4004
rect 6788 3992 6794 4004
rect 7760 3992 7788 4032
rect 8757 4029 8769 4032
rect 8803 4060 8815 4063
rect 9490 4060 9496 4072
rect 8803 4032 9496 4060
rect 8803 4029 8815 4032
rect 8757 4023 8815 4029
rect 9490 4020 9496 4032
rect 9548 4060 9554 4072
rect 9692 4060 9720 4091
rect 9950 4088 9956 4100
rect 10008 4088 10014 4140
rect 10505 4131 10563 4137
rect 10505 4097 10517 4131
rect 10551 4097 10563 4131
rect 10505 4091 10563 4097
rect 10781 4131 10839 4137
rect 10781 4097 10793 4131
rect 10827 4128 10839 4131
rect 11698 4128 11704 4140
rect 10827 4100 11704 4128
rect 10827 4097 10839 4100
rect 10781 4091 10839 4097
rect 10520 4060 10548 4091
rect 11698 4088 11704 4100
rect 11756 4088 11762 4140
rect 14274 4128 14280 4140
rect 14235 4100 14280 4128
rect 14274 4088 14280 4100
rect 14332 4088 14338 4140
rect 14366 4088 14372 4140
rect 14424 4128 14430 4140
rect 14752 4137 14780 4168
rect 15010 4156 15016 4168
rect 15068 4156 15074 4208
rect 17218 4196 17224 4208
rect 17179 4168 17224 4196
rect 17218 4156 17224 4168
rect 17276 4156 17282 4208
rect 14553 4131 14611 4137
rect 14553 4128 14565 4131
rect 14424 4100 14565 4128
rect 14424 4088 14430 4100
rect 9548 4032 9720 4060
rect 9968 4032 10548 4060
rect 14476 4060 14504 4100
rect 14553 4097 14565 4100
rect 14599 4097 14611 4131
rect 14553 4091 14611 4097
rect 14737 4131 14795 4137
rect 14737 4097 14749 4131
rect 14783 4097 14795 4131
rect 14737 4091 14795 4097
rect 15105 4131 15163 4137
rect 15105 4097 15117 4131
rect 15151 4128 15163 4131
rect 15381 4131 15439 4137
rect 15381 4128 15393 4131
rect 15151 4100 15393 4128
rect 15151 4097 15163 4100
rect 15105 4091 15163 4097
rect 15381 4097 15393 4100
rect 15427 4097 15439 4131
rect 15381 4091 15439 4097
rect 15657 4131 15715 4137
rect 15657 4097 15669 4131
rect 15703 4097 15715 4131
rect 15838 4128 15844 4140
rect 15799 4100 15844 4128
rect 15657 4091 15715 4097
rect 15672 4060 15700 4091
rect 15838 4088 15844 4100
rect 15896 4088 15902 4140
rect 16942 4128 16948 4140
rect 17000 4137 17006 4140
rect 17425 4137 17453 4236
rect 17589 4233 17601 4267
rect 17635 4264 17647 4267
rect 17678 4264 17684 4276
rect 17635 4236 17684 4264
rect 17635 4233 17647 4236
rect 17589 4227 17647 4233
rect 17678 4224 17684 4236
rect 17736 4224 17742 4276
rect 18141 4267 18199 4273
rect 18141 4233 18153 4267
rect 18187 4264 18199 4267
rect 18322 4264 18328 4276
rect 18187 4236 18328 4264
rect 18187 4233 18199 4236
rect 18141 4227 18199 4233
rect 18322 4224 18328 4236
rect 18380 4224 18386 4276
rect 20438 4264 20444 4276
rect 19996 4236 20444 4264
rect 18966 4156 18972 4208
rect 19024 4196 19030 4208
rect 19996 4196 20024 4236
rect 20438 4224 20444 4236
rect 20496 4264 20502 4276
rect 21269 4267 21327 4273
rect 21269 4264 21281 4267
rect 20496 4236 21281 4264
rect 20496 4224 20502 4236
rect 21269 4233 21281 4236
rect 21315 4233 21327 4267
rect 29362 4264 29368 4276
rect 29323 4236 29368 4264
rect 21269 4227 21327 4233
rect 29362 4224 29368 4236
rect 29420 4224 29426 4276
rect 22094 4196 22100 4208
rect 19024 4168 20024 4196
rect 20088 4168 22100 4196
rect 19024 4156 19030 4168
rect 16910 4100 16948 4128
rect 16942 4088 16948 4100
rect 17000 4091 17010 4137
rect 17093 4131 17151 4137
rect 17093 4097 17105 4131
rect 17139 4128 17151 4131
rect 17313 4131 17371 4137
rect 17139 4097 17172 4128
rect 17093 4091 17172 4097
rect 17313 4097 17325 4131
rect 17359 4097 17371 4131
rect 17313 4091 17371 4097
rect 17410 4131 17468 4137
rect 17410 4097 17422 4131
rect 17456 4097 17468 4131
rect 17410 4091 17468 4097
rect 17000 4088 17006 4091
rect 14476 4032 15700 4060
rect 9548 4020 9554 4032
rect 7926 3992 7932 4004
rect 6788 3964 7788 3992
rect 7887 3964 7932 3992
rect 6788 3952 6794 3964
rect 7926 3952 7932 3964
rect 7984 3952 7990 4004
rect 3142 3884 3148 3936
rect 3200 3924 3206 3936
rect 5718 3924 5724 3936
rect 3200 3896 5724 3924
rect 3200 3884 3206 3896
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 6365 3927 6423 3933
rect 6365 3893 6377 3927
rect 6411 3924 6423 3927
rect 6638 3924 6644 3936
rect 6411 3896 6644 3924
rect 6411 3893 6423 3896
rect 6365 3887 6423 3893
rect 6638 3884 6644 3896
rect 6696 3884 6702 3936
rect 6914 3884 6920 3936
rect 6972 3924 6978 3936
rect 8021 3927 8079 3933
rect 8021 3924 8033 3927
rect 6972 3896 8033 3924
rect 6972 3884 6978 3896
rect 8021 3893 8033 3896
rect 8067 3893 8079 3927
rect 8021 3887 8079 3893
rect 9217 3927 9275 3933
rect 9217 3893 9229 3927
rect 9263 3924 9275 3927
rect 9968 3924 9996 4032
rect 12802 3952 12808 4004
rect 12860 3992 12866 4004
rect 15197 3995 15255 4001
rect 15197 3992 15209 3995
rect 12860 3964 15209 3992
rect 12860 3952 12866 3964
rect 15197 3961 15209 3964
rect 15243 3961 15255 3995
rect 15197 3955 15255 3961
rect 16942 3952 16948 4004
rect 17000 3992 17006 4004
rect 17144 3992 17172 4091
rect 17000 3964 17172 3992
rect 17319 3992 17347 4091
rect 17862 4088 17868 4140
rect 17920 4128 17926 4140
rect 18325 4131 18383 4137
rect 18325 4128 18337 4131
rect 17920 4100 18337 4128
rect 17920 4088 17926 4100
rect 18325 4097 18337 4100
rect 18371 4097 18383 4131
rect 18598 4128 18604 4140
rect 18559 4100 18604 4128
rect 18325 4091 18383 4097
rect 18598 4088 18604 4100
rect 18656 4088 18662 4140
rect 18782 4128 18788 4140
rect 18743 4100 18788 4128
rect 18782 4088 18788 4100
rect 18840 4088 18846 4140
rect 19334 4088 19340 4140
rect 19392 4128 19398 4140
rect 19429 4131 19487 4137
rect 19429 4128 19441 4131
rect 19392 4100 19441 4128
rect 19392 4088 19398 4100
rect 19429 4097 19441 4100
rect 19475 4097 19487 4131
rect 19429 4091 19487 4097
rect 19889 4131 19947 4137
rect 19889 4097 19901 4131
rect 19935 4128 19947 4131
rect 20088 4128 20116 4168
rect 22094 4156 22100 4168
rect 22152 4156 22158 4208
rect 24854 4156 24860 4208
rect 24912 4196 24918 4208
rect 25222 4196 25228 4208
rect 24912 4168 25228 4196
rect 24912 4156 24918 4168
rect 25222 4156 25228 4168
rect 25280 4196 25286 4208
rect 25280 4168 25636 4196
rect 25280 4156 25286 4168
rect 20162 4137 20168 4140
rect 19935 4100 20116 4128
rect 19935 4097 19947 4100
rect 19889 4091 19947 4097
rect 20156 4091 20168 4137
rect 20220 4128 20226 4140
rect 22002 4128 22008 4140
rect 20220 4100 20256 4128
rect 21963 4100 22008 4128
rect 20162 4088 20168 4091
rect 20220 4088 20226 4100
rect 22002 4088 22008 4100
rect 22060 4088 22066 4140
rect 22554 4128 22560 4140
rect 22515 4100 22560 4128
rect 22554 4088 22560 4100
rect 22612 4088 22618 4140
rect 23842 4128 23848 4140
rect 23803 4100 23848 4128
rect 23842 4088 23848 4100
rect 23900 4088 23906 4140
rect 25608 4137 25636 4168
rect 27338 4156 27344 4208
rect 27396 4196 27402 4208
rect 31294 4196 31300 4208
rect 27396 4168 27441 4196
rect 30300 4168 31300 4196
rect 27396 4156 27402 4168
rect 25317 4131 25375 4137
rect 25317 4097 25329 4131
rect 25363 4097 25375 4131
rect 25317 4091 25375 4097
rect 25593 4131 25651 4137
rect 25593 4097 25605 4131
rect 25639 4097 25651 4131
rect 25593 4091 25651 4097
rect 19150 4060 19156 4072
rect 17512 4032 19156 4060
rect 17512 3992 17540 4032
rect 19150 4020 19156 4032
rect 19208 4020 19214 4072
rect 19242 4020 19248 4072
rect 19300 4060 19306 4072
rect 19300 4032 19380 4060
rect 19300 4020 19306 4032
rect 17319 3964 17540 3992
rect 17000 3952 17006 3964
rect 9263 3896 9996 3924
rect 9263 3893 9275 3896
rect 9217 3887 9275 3893
rect 10594 3884 10600 3936
rect 10652 3924 10658 3936
rect 10689 3927 10747 3933
rect 10689 3924 10701 3927
rect 10652 3896 10701 3924
rect 10652 3884 10658 3896
rect 10689 3893 10701 3896
rect 10735 3893 10747 3927
rect 10689 3887 10747 3893
rect 12894 3884 12900 3936
rect 12952 3924 12958 3936
rect 13173 3927 13231 3933
rect 13173 3924 13185 3927
rect 12952 3896 13185 3924
rect 12952 3884 12958 3896
rect 13173 3893 13185 3896
rect 13219 3893 13231 3927
rect 13173 3887 13231 3893
rect 13262 3884 13268 3936
rect 13320 3924 13326 3936
rect 14093 3927 14151 3933
rect 14093 3924 14105 3927
rect 13320 3896 14105 3924
rect 13320 3884 13326 3896
rect 14093 3893 14105 3896
rect 14139 3893 14151 3927
rect 14093 3887 14151 3893
rect 16758 3884 16764 3936
rect 16816 3924 16822 3936
rect 17678 3924 17684 3936
rect 16816 3896 17684 3924
rect 16816 3884 16822 3896
rect 17678 3884 17684 3896
rect 17736 3884 17742 3936
rect 19242 3924 19248 3936
rect 19203 3896 19248 3924
rect 19242 3884 19248 3896
rect 19300 3884 19306 3936
rect 19352 3924 19380 4032
rect 21174 4020 21180 4072
rect 21232 4060 21238 4072
rect 22646 4060 22652 4072
rect 21232 4032 22652 4060
rect 21232 4020 21238 4032
rect 22646 4020 22652 4032
rect 22704 4060 22710 4072
rect 22833 4063 22891 4069
rect 22833 4060 22845 4063
rect 22704 4032 22845 4060
rect 22704 4020 22710 4032
rect 22833 4029 22845 4032
rect 22879 4060 22891 4063
rect 23198 4060 23204 4072
rect 22879 4032 23204 4060
rect 22879 4029 22891 4032
rect 22833 4023 22891 4029
rect 23198 4020 23204 4032
rect 23256 4020 23262 4072
rect 24118 4060 24124 4072
rect 24079 4032 24124 4060
rect 24118 4020 24124 4032
rect 24176 4020 24182 4072
rect 25038 4020 25044 4072
rect 25096 4060 25102 4072
rect 25332 4060 25360 4091
rect 25682 4088 25688 4140
rect 25740 4128 25746 4140
rect 25777 4131 25835 4137
rect 25777 4128 25789 4131
rect 25740 4100 25789 4128
rect 25740 4088 25746 4100
rect 25777 4097 25789 4100
rect 25823 4097 25835 4131
rect 26418 4128 26424 4140
rect 26379 4100 26424 4128
rect 25777 4091 25835 4097
rect 26418 4088 26424 4100
rect 26476 4088 26482 4140
rect 26602 4088 26608 4140
rect 26660 4128 26666 4140
rect 26973 4131 27031 4137
rect 26973 4128 26985 4131
rect 26660 4100 26985 4128
rect 26660 4088 26666 4100
rect 26973 4097 26985 4100
rect 27019 4097 27031 4131
rect 26973 4091 27031 4097
rect 27062 4088 27068 4140
rect 27120 4128 27126 4140
rect 27246 4128 27252 4140
rect 27120 4100 27165 4128
rect 27207 4100 27252 4128
rect 27120 4088 27126 4100
rect 27246 4088 27252 4100
rect 27304 4088 27310 4140
rect 27438 4131 27496 4137
rect 27438 4097 27450 4131
rect 27484 4097 27496 4131
rect 28258 4128 28264 4140
rect 28219 4100 28264 4128
rect 27438 4091 27496 4097
rect 26326 4060 26332 4072
rect 25096 4032 26332 4060
rect 25096 4020 25102 4032
rect 26326 4020 26332 4032
rect 26384 4020 26390 4072
rect 26694 4020 26700 4072
rect 26752 4060 26758 4072
rect 27453 4060 27481 4091
rect 28258 4088 28264 4100
rect 28316 4088 28322 4140
rect 28534 4128 28540 4140
rect 28495 4100 28540 4128
rect 28534 4088 28540 4100
rect 28592 4088 28598 4140
rect 28721 4131 28779 4137
rect 28721 4097 28733 4131
rect 28767 4097 28779 4131
rect 28721 4091 28779 4097
rect 26752 4032 27481 4060
rect 28736 4060 28764 4091
rect 29454 4088 29460 4140
rect 29512 4128 29518 4140
rect 29549 4131 29607 4137
rect 29549 4128 29561 4131
rect 29512 4100 29561 4128
rect 29512 4088 29518 4100
rect 29549 4097 29561 4100
rect 29595 4097 29607 4131
rect 29822 4128 29828 4140
rect 29783 4100 29828 4128
rect 29549 4091 29607 4097
rect 29822 4088 29828 4100
rect 29880 4128 29886 4140
rect 30300 4128 30328 4168
rect 30466 4128 30472 4140
rect 29880 4100 30328 4128
rect 30427 4100 30472 4128
rect 29880 4088 29886 4100
rect 30466 4088 30472 4100
rect 30524 4088 30530 4140
rect 30742 4128 30748 4140
rect 30703 4100 30748 4128
rect 30742 4088 30748 4100
rect 30800 4088 30806 4140
rect 30944 4137 30972 4168
rect 31294 4156 31300 4168
rect 31352 4156 31358 4208
rect 30929 4131 30987 4137
rect 30929 4097 30941 4131
rect 30975 4097 30987 4131
rect 30929 4091 30987 4097
rect 29086 4060 29092 4072
rect 28736 4032 29092 4060
rect 26752 4020 26758 4032
rect 29086 4020 29092 4032
rect 29144 4060 29150 4072
rect 30098 4060 30104 4072
rect 29144 4032 30104 4060
rect 29144 4020 29150 4032
rect 30098 4020 30104 4032
rect 30156 4020 30162 4072
rect 30285 4063 30343 4069
rect 30285 4029 30297 4063
rect 30331 4060 30343 4063
rect 30558 4060 30564 4072
rect 30331 4032 30564 4060
rect 30331 4029 30343 4032
rect 30285 4023 30343 4029
rect 30558 4020 30564 4032
rect 30616 4020 30622 4072
rect 26237 3995 26295 4001
rect 26237 3992 26249 3995
rect 20824 3964 26249 3992
rect 20824 3924 20852 3964
rect 26237 3961 26249 3964
rect 26283 3961 26295 3995
rect 29730 3992 29736 4004
rect 29691 3964 29736 3992
rect 26237 3955 26295 3961
rect 29730 3952 29736 3964
rect 29788 3952 29794 4004
rect 21818 3924 21824 3936
rect 19352 3896 20852 3924
rect 21779 3896 21824 3924
rect 21818 3884 21824 3896
rect 21876 3884 21882 3936
rect 23566 3884 23572 3936
rect 23624 3924 23630 3936
rect 25133 3927 25191 3933
rect 25133 3924 25145 3927
rect 23624 3896 25145 3924
rect 23624 3884 23630 3896
rect 25133 3893 25145 3896
rect 25179 3893 25191 3927
rect 25133 3887 25191 3893
rect 26050 3884 26056 3936
rect 26108 3924 26114 3936
rect 27617 3927 27675 3933
rect 27617 3924 27629 3927
rect 26108 3896 27629 3924
rect 26108 3884 26114 3896
rect 27617 3893 27629 3896
rect 27663 3893 27675 3927
rect 27617 3887 27675 3893
rect 28077 3927 28135 3933
rect 28077 3893 28089 3927
rect 28123 3924 28135 3927
rect 28626 3924 28632 3936
rect 28123 3896 28632 3924
rect 28123 3893 28135 3896
rect 28077 3887 28135 3893
rect 28626 3884 28632 3896
rect 28684 3884 28690 3936
rect 1104 3834 32016 3856
rect 1104 3782 2136 3834
rect 2188 3782 12440 3834
rect 12492 3782 22744 3834
rect 22796 3782 32016 3834
rect 1104 3760 32016 3782
rect 2317 3723 2375 3729
rect 2317 3689 2329 3723
rect 2363 3720 2375 3723
rect 5074 3720 5080 3732
rect 2363 3692 5080 3720
rect 2363 3689 2375 3692
rect 2317 3683 2375 3689
rect 5074 3680 5080 3692
rect 5132 3680 5138 3732
rect 5442 3720 5448 3732
rect 5403 3692 5448 3720
rect 5442 3680 5448 3692
rect 5500 3680 5506 3732
rect 5718 3680 5724 3732
rect 5776 3720 5782 3732
rect 5813 3723 5871 3729
rect 5813 3720 5825 3723
rect 5776 3692 5825 3720
rect 5776 3680 5782 3692
rect 5813 3689 5825 3692
rect 5859 3720 5871 3723
rect 6086 3720 6092 3732
rect 5859 3692 6092 3720
rect 5859 3689 5871 3692
rect 5813 3683 5871 3689
rect 6086 3680 6092 3692
rect 6144 3680 6150 3732
rect 7929 3723 7987 3729
rect 7929 3689 7941 3723
rect 7975 3720 7987 3723
rect 12710 3720 12716 3732
rect 7975 3692 12716 3720
rect 7975 3689 7987 3692
rect 7929 3683 7987 3689
rect 12710 3680 12716 3692
rect 12768 3680 12774 3732
rect 12897 3723 12955 3729
rect 12897 3689 12909 3723
rect 12943 3720 12955 3723
rect 13814 3720 13820 3732
rect 12943 3692 13820 3720
rect 12943 3689 12955 3692
rect 12897 3683 12955 3689
rect 13814 3680 13820 3692
rect 13872 3680 13878 3732
rect 17034 3680 17040 3732
rect 17092 3720 17098 3732
rect 17313 3723 17371 3729
rect 17313 3720 17325 3723
rect 17092 3692 17325 3720
rect 17092 3680 17098 3692
rect 17313 3689 17325 3692
rect 17359 3689 17371 3723
rect 19245 3723 19303 3729
rect 19245 3720 19257 3723
rect 17313 3683 17371 3689
rect 18248 3692 19257 3720
rect 3142 3652 3148 3664
rect 3103 3624 3148 3652
rect 3142 3612 3148 3624
rect 3200 3612 3206 3664
rect 3513 3655 3571 3661
rect 3513 3621 3525 3655
rect 3559 3652 3571 3655
rect 3559 3624 6408 3652
rect 3559 3621 3571 3624
rect 3513 3615 3571 3621
rect 1949 3587 2007 3593
rect 1949 3553 1961 3587
rect 1995 3584 2007 3587
rect 2682 3584 2688 3596
rect 1995 3556 2688 3584
rect 1995 3553 2007 3556
rect 1949 3547 2007 3553
rect 2682 3544 2688 3556
rect 2740 3584 2746 3596
rect 2740 3556 3648 3584
rect 2740 3544 2746 3556
rect 2133 3519 2191 3525
rect 2133 3485 2145 3519
rect 2179 3516 2191 3519
rect 2406 3516 2412 3528
rect 2179 3488 2412 3516
rect 2179 3485 2191 3488
rect 2133 3479 2191 3485
rect 2406 3476 2412 3488
rect 2464 3476 2470 3528
rect 2961 3519 3019 3525
rect 2961 3485 2973 3519
rect 3007 3485 3019 3519
rect 2961 3479 3019 3485
rect 3237 3519 3295 3525
rect 3237 3485 3249 3519
rect 3283 3516 3295 3519
rect 3513 3519 3571 3525
rect 3513 3516 3525 3519
rect 3283 3488 3525 3516
rect 3283 3485 3295 3488
rect 3237 3479 3295 3485
rect 3513 3485 3525 3488
rect 3559 3485 3571 3519
rect 3620 3516 3648 3556
rect 3694 3544 3700 3596
rect 3752 3584 3758 3596
rect 4157 3587 4215 3593
rect 4157 3584 4169 3587
rect 3752 3556 4169 3584
rect 3752 3544 3758 3556
rect 4157 3553 4169 3556
rect 4203 3584 4215 3587
rect 4522 3584 4528 3596
rect 4203 3556 4528 3584
rect 4203 3553 4215 3556
rect 4157 3547 4215 3553
rect 4522 3544 4528 3556
rect 4580 3544 4586 3596
rect 5905 3587 5963 3593
rect 5905 3553 5917 3587
rect 5951 3584 5963 3587
rect 6270 3584 6276 3596
rect 5951 3556 6276 3584
rect 5951 3553 5963 3556
rect 5905 3547 5963 3553
rect 6270 3544 6276 3556
rect 6328 3544 6334 3596
rect 4338 3516 4344 3528
rect 3620 3488 4344 3516
rect 3513 3479 3571 3485
rect 2976 3448 3004 3479
rect 4338 3476 4344 3488
rect 4396 3516 4402 3528
rect 4433 3519 4491 3525
rect 4433 3516 4445 3519
rect 4396 3488 4445 3516
rect 4396 3476 4402 3488
rect 4433 3485 4445 3488
rect 4479 3485 4491 3519
rect 4433 3479 4491 3485
rect 5166 3476 5172 3528
rect 5224 3516 5230 3528
rect 5629 3519 5687 3525
rect 5629 3516 5641 3519
rect 5224 3488 5641 3516
rect 5224 3476 5230 3488
rect 5629 3485 5641 3488
rect 5675 3485 5687 3519
rect 5629 3479 5687 3485
rect 6086 3448 6092 3460
rect 2976 3420 5028 3448
rect 2777 3383 2835 3389
rect 2777 3349 2789 3383
rect 2823 3380 2835 3383
rect 4706 3380 4712 3392
rect 2823 3352 4712 3380
rect 2823 3349 2835 3352
rect 2777 3343 2835 3349
rect 4706 3340 4712 3352
rect 4764 3340 4770 3392
rect 5000 3380 5028 3420
rect 5184 3420 6092 3448
rect 5184 3380 5212 3420
rect 6086 3408 6092 3420
rect 6144 3408 6150 3460
rect 5000 3352 5212 3380
rect 6380 3380 6408 3624
rect 9214 3612 9220 3664
rect 9272 3652 9278 3664
rect 9272 3624 10364 3652
rect 9272 3612 9278 3624
rect 6822 3544 6828 3596
rect 6880 3544 6886 3596
rect 6914 3516 6920 3528
rect 6472 3488 6776 3516
rect 6875 3488 6920 3516
rect 6472 3460 6500 3488
rect 6454 3408 6460 3460
rect 6512 3408 6518 3460
rect 6638 3448 6644 3460
rect 6599 3420 6644 3448
rect 6638 3408 6644 3420
rect 6696 3408 6702 3460
rect 6748 3448 6776 3488
rect 6914 3476 6920 3488
rect 6972 3476 6978 3528
rect 9214 3516 9220 3528
rect 9175 3488 9220 3516
rect 9214 3476 9220 3488
rect 9272 3476 9278 3528
rect 9490 3516 9496 3528
rect 9451 3488 9496 3516
rect 9490 3476 9496 3488
rect 9548 3476 9554 3528
rect 9677 3519 9735 3525
rect 9677 3485 9689 3519
rect 9723 3516 9735 3519
rect 9766 3516 9772 3528
rect 9723 3488 9772 3516
rect 9723 3485 9735 3488
rect 9677 3479 9735 3485
rect 9766 3476 9772 3488
rect 9824 3476 9830 3528
rect 10336 3525 10364 3624
rect 10686 3612 10692 3664
rect 10744 3652 10750 3664
rect 13357 3655 13415 3661
rect 10744 3624 11100 3652
rect 10744 3612 10750 3624
rect 10321 3519 10379 3525
rect 10321 3485 10333 3519
rect 10367 3485 10379 3519
rect 10321 3479 10379 3485
rect 10410 3476 10416 3528
rect 10468 3516 10474 3528
rect 10597 3519 10655 3525
rect 10597 3516 10609 3519
rect 10468 3488 10609 3516
rect 10468 3476 10474 3488
rect 10597 3485 10609 3488
rect 10643 3516 10655 3519
rect 10686 3516 10692 3528
rect 10643 3488 10692 3516
rect 10643 3485 10655 3488
rect 10597 3479 10655 3485
rect 10686 3476 10692 3488
rect 10744 3476 10750 3528
rect 10781 3519 10839 3525
rect 10781 3485 10793 3519
rect 10827 3485 10839 3519
rect 10781 3479 10839 3485
rect 7009 3451 7067 3457
rect 7009 3448 7021 3451
rect 6748 3420 7021 3448
rect 7009 3417 7021 3420
rect 7055 3417 7067 3451
rect 7009 3411 7067 3417
rect 7377 3451 7435 3457
rect 7377 3417 7389 3451
rect 7423 3448 7435 3451
rect 7558 3448 7564 3460
rect 7423 3420 7564 3448
rect 7423 3417 7435 3420
rect 7377 3411 7435 3417
rect 7558 3408 7564 3420
rect 7616 3408 7622 3460
rect 7834 3408 7840 3460
rect 7892 3448 7898 3460
rect 10796 3448 10824 3479
rect 10962 3448 10968 3460
rect 7892 3420 10968 3448
rect 7892 3408 7898 3420
rect 10962 3408 10968 3420
rect 11020 3408 11026 3460
rect 11072 3448 11100 3624
rect 13357 3621 13369 3655
rect 13403 3652 13415 3655
rect 16850 3652 16856 3664
rect 13403 3624 16856 3652
rect 13403 3621 13415 3624
rect 13357 3615 13415 3621
rect 16850 3612 16856 3624
rect 16908 3652 16914 3664
rect 16908 3624 17081 3652
rect 16908 3612 16914 3624
rect 11330 3544 11336 3596
rect 11388 3584 11394 3596
rect 11517 3587 11575 3593
rect 11517 3584 11529 3587
rect 11388 3556 11529 3584
rect 11388 3544 11394 3556
rect 11517 3553 11529 3556
rect 11563 3553 11575 3587
rect 11517 3547 11575 3553
rect 13170 3544 13176 3596
rect 13228 3584 13234 3596
rect 15286 3584 15292 3596
rect 13228 3556 15292 3584
rect 13228 3544 13234 3556
rect 11790 3525 11796 3528
rect 11784 3516 11796 3525
rect 11751 3488 11796 3516
rect 11784 3479 11796 3488
rect 11790 3476 11796 3479
rect 11848 3476 11854 3528
rect 13372 3525 13400 3556
rect 15286 3544 15292 3556
rect 15344 3544 15350 3596
rect 15381 3587 15439 3593
rect 15381 3553 15393 3587
rect 15427 3584 15439 3587
rect 15470 3584 15476 3596
rect 15427 3556 15476 3584
rect 15427 3553 15439 3556
rect 15381 3547 15439 3553
rect 15470 3544 15476 3556
rect 15528 3544 15534 3596
rect 15562 3544 15568 3596
rect 15620 3584 15626 3596
rect 16482 3584 16488 3596
rect 15620 3556 16488 3584
rect 15620 3544 15626 3556
rect 16482 3544 16488 3556
rect 16540 3584 16546 3596
rect 16540 3556 16988 3584
rect 16540 3544 16546 3556
rect 13357 3519 13415 3525
rect 13357 3485 13369 3519
rect 13403 3485 13415 3519
rect 13538 3516 13544 3528
rect 13499 3488 13544 3516
rect 13357 3479 13415 3485
rect 13538 3476 13544 3488
rect 13596 3476 13602 3528
rect 14274 3516 14280 3528
rect 14235 3488 14280 3516
rect 14274 3476 14280 3488
rect 14332 3476 14338 3528
rect 14366 3476 14372 3528
rect 14424 3516 14430 3528
rect 14553 3519 14611 3525
rect 14553 3516 14565 3519
rect 14424 3488 14565 3516
rect 14424 3476 14430 3488
rect 14553 3485 14565 3488
rect 14599 3485 14611 3519
rect 14553 3479 14611 3485
rect 14737 3519 14795 3525
rect 14737 3485 14749 3519
rect 14783 3516 14795 3519
rect 14826 3516 14832 3528
rect 14783 3488 14832 3516
rect 14783 3485 14795 3488
rect 14737 3479 14795 3485
rect 14826 3476 14832 3488
rect 14884 3476 14890 3528
rect 15657 3519 15715 3525
rect 15657 3485 15669 3519
rect 15703 3516 15715 3519
rect 16022 3516 16028 3528
rect 15703 3488 16028 3516
rect 15703 3485 15715 3488
rect 15657 3479 15715 3485
rect 16022 3476 16028 3488
rect 16080 3476 16086 3528
rect 16574 3476 16580 3528
rect 16632 3516 16638 3528
rect 16669 3519 16727 3525
rect 16669 3516 16681 3519
rect 16632 3488 16681 3516
rect 16632 3476 16638 3488
rect 16669 3485 16681 3488
rect 16715 3485 16727 3519
rect 16669 3479 16727 3485
rect 16758 3476 16764 3528
rect 16816 3516 16822 3528
rect 16960 3525 16988 3556
rect 16945 3519 17003 3525
rect 16816 3488 16861 3516
rect 16816 3476 16822 3488
rect 16945 3485 16957 3519
rect 16991 3485 17003 3519
rect 17053 3516 17081 3624
rect 17134 3519 17192 3525
rect 17134 3516 17146 3519
rect 17053 3488 17146 3516
rect 16945 3479 17003 3485
rect 17134 3485 17146 3488
rect 17180 3485 17192 3519
rect 17134 3479 17192 3485
rect 17862 3476 17868 3528
rect 17920 3516 17926 3528
rect 18248 3525 18276 3692
rect 19245 3689 19257 3692
rect 19291 3689 19303 3723
rect 19886 3720 19892 3732
rect 19847 3692 19892 3720
rect 19245 3683 19303 3689
rect 19886 3680 19892 3692
rect 19944 3680 19950 3732
rect 20990 3720 20996 3732
rect 20951 3692 20996 3720
rect 20990 3680 20996 3692
rect 21048 3680 21054 3732
rect 23385 3723 23443 3729
rect 23385 3689 23397 3723
rect 23431 3720 23443 3723
rect 23658 3720 23664 3732
rect 23431 3692 23664 3720
rect 23431 3689 23443 3692
rect 23385 3683 23443 3689
rect 23658 3680 23664 3692
rect 23716 3680 23722 3732
rect 23750 3680 23756 3732
rect 23808 3720 23814 3732
rect 26234 3720 26240 3732
rect 23808 3692 26240 3720
rect 23808 3680 23814 3692
rect 26234 3680 26240 3692
rect 26292 3680 26298 3732
rect 26513 3723 26571 3729
rect 26513 3689 26525 3723
rect 26559 3720 26571 3723
rect 26602 3720 26608 3732
rect 26559 3692 26608 3720
rect 26559 3689 26571 3692
rect 26513 3683 26571 3689
rect 26602 3680 26608 3692
rect 26660 3680 26666 3732
rect 30650 3720 30656 3732
rect 30611 3692 30656 3720
rect 30650 3680 30656 3692
rect 30708 3680 30714 3732
rect 20898 3612 20904 3664
rect 20956 3652 20962 3664
rect 20956 3624 21496 3652
rect 20956 3612 20962 3624
rect 18322 3544 18328 3596
rect 18380 3584 18386 3596
rect 18380 3556 18736 3584
rect 18380 3544 18386 3556
rect 18708 3528 18736 3556
rect 19242 3544 19248 3596
rect 19300 3584 19306 3596
rect 21468 3584 21496 3624
rect 21542 3612 21548 3664
rect 21600 3652 21606 3664
rect 26418 3652 26424 3664
rect 21600 3624 26424 3652
rect 21600 3612 21606 3624
rect 26418 3612 26424 3624
rect 26476 3612 26482 3664
rect 29730 3612 29736 3664
rect 29788 3652 29794 3664
rect 31018 3652 31024 3664
rect 29788 3624 31024 3652
rect 29788 3612 29794 3624
rect 31018 3612 31024 3624
rect 31076 3612 31082 3664
rect 24118 3584 24124 3596
rect 19300 3556 21220 3584
rect 19300 3544 19306 3556
rect 18233 3519 18291 3525
rect 18233 3516 18245 3519
rect 17920 3488 18245 3516
rect 17920 3476 17926 3488
rect 18233 3485 18245 3488
rect 18279 3485 18291 3519
rect 18233 3479 18291 3485
rect 18509 3519 18567 3525
rect 18509 3485 18521 3519
rect 18555 3485 18567 3519
rect 18509 3479 18567 3485
rect 16482 3448 16488 3460
rect 11072 3420 16488 3448
rect 16482 3408 16488 3420
rect 16540 3408 16546 3460
rect 17034 3408 17040 3460
rect 17092 3448 17098 3460
rect 17092 3420 17137 3448
rect 17092 3408 17098 3420
rect 17218 3408 17224 3460
rect 17276 3448 17282 3460
rect 18524 3448 18552 3479
rect 18690 3476 18696 3528
rect 18748 3516 18754 3528
rect 18748 3488 18841 3516
rect 18748 3476 18754 3488
rect 19334 3476 19340 3528
rect 19392 3516 19398 3528
rect 20088 3525 20116 3556
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 19392 3488 19441 3516
rect 19392 3476 19398 3488
rect 19429 3485 19441 3488
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 20073 3519 20131 3525
rect 20073 3485 20085 3519
rect 20119 3516 20131 3519
rect 20254 3516 20260 3528
rect 20119 3488 20260 3516
rect 20119 3485 20131 3488
rect 20073 3479 20131 3485
rect 20254 3476 20260 3488
rect 20312 3476 20318 3528
rect 20349 3519 20407 3525
rect 20349 3485 20361 3519
rect 20395 3485 20407 3519
rect 20349 3479 20407 3485
rect 20533 3519 20591 3525
rect 20533 3485 20545 3519
rect 20579 3516 20591 3519
rect 20622 3516 20628 3528
rect 20579 3488 20628 3516
rect 20579 3485 20591 3488
rect 20533 3479 20591 3485
rect 18598 3448 18604 3460
rect 17276 3420 18604 3448
rect 17276 3408 17282 3420
rect 18598 3408 18604 3420
rect 18656 3408 18662 3460
rect 20364 3448 20392 3479
rect 20622 3476 20628 3488
rect 20680 3476 20686 3528
rect 21192 3525 21220 3556
rect 21468 3556 24124 3584
rect 21468 3525 21496 3556
rect 22572 3528 22600 3556
rect 24118 3544 24124 3556
rect 24176 3544 24182 3596
rect 28350 3584 28356 3596
rect 25976 3556 28356 3584
rect 21177 3519 21235 3525
rect 21177 3485 21189 3519
rect 21223 3485 21235 3519
rect 21177 3479 21235 3485
rect 21453 3519 21511 3525
rect 21453 3485 21465 3519
rect 21499 3485 21511 3519
rect 21453 3479 21511 3485
rect 21637 3519 21695 3525
rect 21637 3485 21649 3519
rect 21683 3516 21695 3519
rect 22186 3516 22192 3528
rect 21683 3488 22192 3516
rect 21683 3485 21695 3488
rect 21637 3479 21695 3485
rect 20898 3448 20904 3460
rect 20364 3420 20904 3448
rect 20898 3408 20904 3420
rect 20956 3408 20962 3460
rect 21192 3448 21220 3479
rect 22186 3476 22192 3488
rect 22244 3476 22250 3528
rect 22278 3476 22284 3528
rect 22336 3516 22342 3528
rect 22554 3516 22560 3528
rect 22336 3488 22429 3516
rect 22467 3488 22560 3516
rect 22336 3476 22342 3488
rect 22554 3476 22560 3488
rect 22612 3476 22618 3528
rect 22741 3519 22799 3525
rect 22741 3485 22753 3519
rect 22787 3516 22799 3519
rect 22830 3516 22836 3528
rect 22787 3488 22836 3516
rect 22787 3485 22799 3488
rect 22741 3479 22799 3485
rect 22830 3476 22836 3488
rect 22888 3476 22894 3528
rect 23566 3516 23572 3528
rect 23527 3488 23572 3516
rect 23566 3476 23572 3488
rect 23624 3476 23630 3528
rect 23845 3519 23903 3525
rect 23845 3485 23857 3519
rect 23891 3485 23903 3519
rect 23845 3479 23903 3485
rect 24949 3519 25007 3525
rect 24949 3485 24961 3519
rect 24995 3516 25007 3519
rect 25038 3516 25044 3528
rect 24995 3488 25044 3516
rect 24995 3485 25007 3488
rect 24949 3479 25007 3485
rect 22287 3448 22315 3476
rect 21192 3420 22315 3448
rect 23860 3448 23888 3479
rect 25038 3476 25044 3488
rect 25096 3476 25102 3528
rect 25222 3516 25228 3528
rect 25183 3488 25228 3516
rect 25222 3476 25228 3488
rect 25280 3476 25286 3528
rect 25409 3519 25467 3525
rect 25409 3485 25421 3519
rect 25455 3516 25467 3519
rect 25590 3516 25596 3528
rect 25455 3488 25596 3516
rect 25455 3485 25467 3488
rect 25409 3479 25467 3485
rect 25424 3448 25452 3479
rect 25590 3476 25596 3488
rect 25648 3476 25654 3528
rect 25976 3525 26004 3556
rect 28350 3544 28356 3556
rect 28408 3544 28414 3596
rect 28626 3544 28632 3596
rect 28684 3584 28690 3596
rect 31110 3584 31116 3596
rect 28684 3556 30880 3584
rect 31071 3556 31116 3584
rect 28684 3544 28690 3556
rect 25961 3519 26019 3525
rect 25961 3485 25973 3519
rect 26007 3485 26019 3519
rect 26142 3516 26148 3528
rect 26103 3488 26148 3516
rect 25961 3479 26019 3485
rect 26142 3476 26148 3488
rect 26200 3476 26206 3528
rect 26329 3519 26387 3525
rect 26329 3485 26341 3519
rect 26375 3516 26387 3519
rect 26510 3516 26516 3528
rect 26375 3488 26516 3516
rect 26375 3485 26387 3488
rect 26329 3479 26387 3485
rect 26510 3476 26516 3488
rect 26568 3476 26574 3528
rect 26970 3516 26976 3528
rect 26931 3488 26976 3516
rect 26970 3476 26976 3488
rect 27028 3476 27034 3528
rect 27706 3476 27712 3528
rect 27764 3516 27770 3528
rect 29730 3516 29736 3528
rect 27764 3488 29592 3516
rect 29691 3488 29736 3516
rect 27764 3476 27770 3488
rect 23860 3420 25452 3448
rect 26237 3451 26295 3457
rect 26237 3417 26249 3451
rect 26283 3417 26295 3451
rect 28718 3448 28724 3460
rect 28679 3420 28724 3448
rect 26237 3411 26295 3417
rect 7098 3380 7104 3392
rect 6380 3352 7104 3380
rect 7098 3340 7104 3352
rect 7156 3340 7162 3392
rect 7742 3380 7748 3392
rect 7703 3352 7748 3380
rect 7742 3340 7748 3352
rect 7800 3340 7806 3392
rect 9033 3383 9091 3389
rect 9033 3349 9045 3383
rect 9079 3380 9091 3383
rect 10042 3380 10048 3392
rect 9079 3352 10048 3380
rect 9079 3349 9091 3352
rect 9033 3343 9091 3349
rect 10042 3340 10048 3352
rect 10100 3340 10106 3392
rect 10137 3383 10195 3389
rect 10137 3349 10149 3383
rect 10183 3380 10195 3383
rect 11606 3380 11612 3392
rect 10183 3352 11612 3380
rect 10183 3349 10195 3352
rect 10137 3343 10195 3349
rect 11606 3340 11612 3352
rect 11664 3340 11670 3392
rect 13538 3340 13544 3392
rect 13596 3380 13602 3392
rect 14093 3383 14151 3389
rect 14093 3380 14105 3383
rect 13596 3352 14105 3380
rect 13596 3340 13602 3352
rect 14093 3349 14105 3352
rect 14139 3349 14151 3383
rect 14093 3343 14151 3349
rect 18049 3383 18107 3389
rect 18049 3349 18061 3383
rect 18095 3380 18107 3383
rect 18414 3380 18420 3392
rect 18095 3352 18420 3380
rect 18095 3349 18107 3352
rect 18049 3343 18107 3349
rect 18414 3340 18420 3352
rect 18472 3340 18478 3392
rect 19794 3340 19800 3392
rect 19852 3380 19858 3392
rect 22097 3383 22155 3389
rect 22097 3380 22109 3383
rect 19852 3352 22109 3380
rect 19852 3340 19858 3352
rect 22097 3349 22109 3352
rect 22143 3349 22155 3383
rect 22097 3343 22155 3349
rect 24765 3383 24823 3389
rect 24765 3349 24777 3383
rect 24811 3380 24823 3383
rect 24854 3380 24860 3392
rect 24811 3352 24860 3380
rect 24811 3349 24823 3352
rect 24765 3343 24823 3349
rect 24854 3340 24860 3352
rect 24912 3340 24918 3392
rect 25866 3340 25872 3392
rect 25924 3380 25930 3392
rect 26252 3380 26280 3411
rect 28718 3408 28724 3420
rect 28776 3408 28782 3460
rect 29564 3448 29592 3488
rect 29730 3476 29736 3488
rect 29788 3476 29794 3528
rect 30006 3516 30012 3528
rect 29967 3488 30012 3516
rect 30006 3476 30012 3488
rect 30064 3476 30070 3528
rect 30852 3525 30880 3556
rect 31110 3544 31116 3556
rect 31168 3544 31174 3596
rect 30193 3519 30251 3525
rect 30193 3485 30205 3519
rect 30239 3485 30251 3519
rect 30193 3479 30251 3485
rect 30837 3519 30895 3525
rect 30837 3485 30849 3519
rect 30883 3485 30895 3519
rect 30837 3479 30895 3485
rect 30208 3448 30236 3479
rect 30742 3448 30748 3460
rect 29564 3420 30748 3448
rect 30742 3408 30748 3420
rect 30800 3408 30806 3460
rect 25924 3352 26280 3380
rect 29549 3383 29607 3389
rect 25924 3340 25930 3352
rect 29549 3349 29561 3383
rect 29595 3380 29607 3383
rect 30558 3380 30564 3392
rect 29595 3352 30564 3380
rect 29595 3349 29607 3352
rect 29549 3343 29607 3349
rect 30558 3340 30564 3352
rect 30616 3340 30622 3392
rect 1104 3290 32016 3312
rect 1104 3238 7288 3290
rect 7340 3238 17592 3290
rect 17644 3238 27896 3290
rect 27948 3238 32016 3290
rect 1104 3216 32016 3238
rect 2774 3136 2780 3188
rect 2832 3176 2838 3188
rect 9674 3176 9680 3188
rect 2832 3148 9680 3176
rect 2832 3136 2838 3148
rect 9674 3136 9680 3148
rect 9732 3136 9738 3188
rect 11698 3176 11704 3188
rect 9784 3148 11704 3176
rect 2222 3108 2228 3120
rect 2135 3080 2228 3108
rect 2148 3049 2176 3080
rect 2222 3068 2228 3080
rect 2280 3108 2286 3120
rect 4338 3108 4344 3120
rect 2280 3080 2774 3108
rect 2280 3068 2286 3080
rect 2133 3043 2191 3049
rect 2133 3009 2145 3043
rect 2179 3009 2191 3043
rect 2133 3003 2191 3009
rect 2314 3000 2320 3052
rect 2372 3040 2378 3052
rect 2409 3043 2467 3049
rect 2409 3040 2421 3043
rect 2372 3012 2421 3040
rect 2372 3000 2378 3012
rect 2409 3009 2421 3012
rect 2455 3009 2467 3043
rect 2590 3040 2596 3052
rect 2551 3012 2596 3040
rect 2409 3003 2467 3009
rect 2424 2972 2452 3003
rect 2590 3000 2596 3012
rect 2648 3000 2654 3052
rect 2746 3040 2774 3080
rect 3712 3080 4344 3108
rect 3712 3049 3740 3080
rect 4338 3068 4344 3080
rect 4396 3068 4402 3120
rect 5997 3111 6055 3117
rect 5997 3108 6009 3111
rect 4540 3080 6009 3108
rect 3237 3043 3295 3049
rect 3237 3040 3249 3043
rect 2746 3012 3249 3040
rect 3237 3009 3249 3012
rect 3283 3009 3295 3043
rect 3237 3003 3295 3009
rect 3513 3043 3571 3049
rect 3513 3009 3525 3043
rect 3559 3009 3571 3043
rect 3513 3003 3571 3009
rect 3697 3043 3755 3049
rect 3697 3009 3709 3043
rect 3743 3009 3755 3043
rect 3697 3003 3755 3009
rect 3528 2972 3556 3003
rect 4154 3000 4160 3052
rect 4212 3040 4218 3052
rect 4433 3043 4491 3049
rect 4433 3040 4445 3043
rect 4212 3012 4445 3040
rect 4212 3000 4218 3012
rect 4433 3009 4445 3012
rect 4479 3009 4491 3043
rect 4433 3003 4491 3009
rect 2424 2944 3556 2972
rect 3970 2932 3976 2984
rect 4028 2972 4034 2984
rect 4540 2972 4568 3080
rect 5997 3077 6009 3080
rect 6043 3077 6055 3111
rect 5997 3071 6055 3077
rect 6086 3068 6092 3120
rect 6144 3108 6150 3120
rect 6365 3111 6423 3117
rect 6365 3108 6377 3111
rect 6144 3080 6377 3108
rect 6144 3068 6150 3080
rect 6365 3077 6377 3080
rect 6411 3077 6423 3111
rect 6365 3071 6423 3077
rect 7742 3068 7748 3120
rect 7800 3108 7806 3120
rect 9125 3111 9183 3117
rect 9125 3108 9137 3111
rect 7800 3080 9137 3108
rect 7800 3068 7806 3080
rect 9125 3077 9137 3080
rect 9171 3077 9183 3111
rect 9784 3108 9812 3148
rect 11698 3136 11704 3148
rect 11756 3136 11762 3188
rect 13814 3136 13820 3188
rect 13872 3176 13878 3188
rect 14185 3179 14243 3185
rect 14185 3176 14197 3179
rect 13872 3148 14197 3176
rect 13872 3136 13878 3148
rect 14185 3145 14197 3148
rect 14231 3176 14243 3179
rect 14826 3176 14832 3188
rect 14231 3148 14832 3176
rect 14231 3145 14243 3148
rect 14185 3139 14243 3145
rect 14826 3136 14832 3148
rect 14884 3136 14890 3188
rect 15562 3136 15568 3188
rect 15620 3176 15626 3188
rect 15841 3179 15899 3185
rect 15841 3176 15853 3179
rect 15620 3148 15853 3176
rect 15620 3136 15626 3148
rect 15841 3145 15853 3148
rect 15887 3145 15899 3179
rect 15841 3139 15899 3145
rect 17678 3136 17684 3188
rect 17736 3176 17742 3188
rect 18877 3179 18935 3185
rect 18877 3176 18889 3179
rect 17736 3148 18889 3176
rect 17736 3136 17742 3148
rect 18877 3145 18889 3148
rect 18923 3145 18935 3179
rect 18877 3139 18935 3145
rect 20070 3136 20076 3188
rect 20128 3176 20134 3188
rect 20441 3179 20499 3185
rect 20441 3176 20453 3179
rect 20128 3148 20453 3176
rect 20128 3136 20134 3148
rect 20441 3145 20453 3148
rect 20487 3145 20499 3179
rect 28721 3179 28779 3185
rect 28721 3176 28733 3179
rect 20441 3139 20499 3145
rect 20548 3148 28733 3176
rect 9125 3071 9183 3077
rect 9223 3080 9812 3108
rect 4700 3043 4758 3049
rect 4700 3009 4712 3043
rect 4746 3040 4758 3043
rect 6270 3040 6276 3052
rect 4746 3012 6276 3040
rect 4746 3009 4758 3012
rect 4700 3003 4758 3009
rect 6270 3000 6276 3012
rect 6328 3000 6334 3052
rect 6546 3040 6552 3052
rect 6507 3012 6552 3040
rect 6546 3000 6552 3012
rect 6604 3000 6610 3052
rect 6730 3000 6736 3052
rect 6788 3040 6794 3052
rect 6825 3043 6883 3049
rect 6825 3040 6837 3043
rect 6788 3012 6837 3040
rect 6788 3000 6794 3012
rect 6825 3009 6837 3012
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 6914 3000 6920 3052
rect 6972 3040 6978 3052
rect 7009 3043 7067 3049
rect 7009 3040 7021 3043
rect 6972 3012 7021 3040
rect 6972 3000 6978 3012
rect 7009 3009 7021 3012
rect 7055 3009 7067 3043
rect 7009 3003 7067 3009
rect 7377 3043 7435 3049
rect 7377 3009 7389 3043
rect 7423 3040 7435 3043
rect 7929 3043 7987 3049
rect 7929 3040 7941 3043
rect 7423 3012 7941 3040
rect 7423 3009 7435 3012
rect 7377 3003 7435 3009
rect 7929 3009 7941 3012
rect 7975 3040 7987 3043
rect 8662 3040 8668 3052
rect 7975 3012 8668 3040
rect 7975 3009 7987 3012
rect 7929 3003 7987 3009
rect 8662 3000 8668 3012
rect 8720 3000 8726 3052
rect 8938 3040 8944 3052
rect 8899 3012 8944 3040
rect 8938 3000 8944 3012
rect 8996 3040 9002 3052
rect 9223 3040 9251 3080
rect 10594 3068 10600 3120
rect 10652 3108 10658 3120
rect 11149 3111 11207 3117
rect 11149 3108 11161 3111
rect 10652 3080 11161 3108
rect 10652 3068 10658 3080
rect 11149 3077 11161 3080
rect 11195 3077 11207 3111
rect 11149 3071 11207 3077
rect 11330 3068 11336 3120
rect 11388 3108 11394 3120
rect 11388 3080 11836 3108
rect 11388 3068 11394 3080
rect 9582 3040 9588 3052
rect 8996 3012 9251 3040
rect 9543 3012 9588 3040
rect 8996 3000 9002 3012
rect 9582 3000 9588 3012
rect 9640 3000 9646 3052
rect 9852 3043 9910 3049
rect 9852 3009 9864 3043
rect 9898 3040 9910 3043
rect 9898 3012 10732 3040
rect 9898 3009 9910 3012
rect 9852 3003 9910 3009
rect 8021 2975 8079 2981
rect 8021 2972 8033 2975
rect 4028 2944 4568 2972
rect 5460 2944 8033 2972
rect 4028 2932 4034 2944
rect 3510 2864 3516 2916
rect 3568 2904 3574 2916
rect 4430 2904 4436 2916
rect 3568 2876 4436 2904
rect 3568 2864 3574 2876
rect 4430 2864 4436 2876
rect 4488 2864 4494 2916
rect 1949 2839 2007 2845
rect 1949 2805 1961 2839
rect 1995 2836 2007 2839
rect 2314 2836 2320 2848
rect 1995 2808 2320 2836
rect 1995 2805 2007 2808
rect 1949 2799 2007 2805
rect 2314 2796 2320 2808
rect 2372 2796 2378 2848
rect 3053 2839 3111 2845
rect 3053 2805 3065 2839
rect 3099 2836 3111 2839
rect 3326 2836 3332 2848
rect 3099 2808 3332 2836
rect 3099 2805 3111 2808
rect 3053 2799 3111 2805
rect 3326 2796 3332 2808
rect 3384 2796 3390 2848
rect 3786 2796 3792 2848
rect 3844 2836 3850 2848
rect 4798 2836 4804 2848
rect 3844 2808 4804 2836
rect 3844 2796 3850 2808
rect 4798 2796 4804 2808
rect 4856 2836 4862 2848
rect 5460 2836 5488 2944
rect 8021 2941 8033 2944
rect 8067 2941 8079 2975
rect 8202 2972 8208 2984
rect 8163 2944 8208 2972
rect 8021 2935 8079 2941
rect 8202 2932 8208 2944
rect 8260 2932 8266 2984
rect 8757 2975 8815 2981
rect 8757 2941 8769 2975
rect 8803 2941 8815 2975
rect 10704 2972 10732 3012
rect 11606 3000 11612 3052
rect 11664 3040 11670 3052
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 11664 3012 11713 3040
rect 11664 3000 11670 3012
rect 11701 3009 11713 3012
rect 11747 3009 11759 3043
rect 11808 3040 11836 3080
rect 12710 3068 12716 3120
rect 12768 3108 12774 3120
rect 12768 3080 13860 3108
rect 12768 3068 12774 3080
rect 12805 3043 12863 3049
rect 12805 3040 12817 3043
rect 11808 3012 12817 3040
rect 11701 3003 11759 3009
rect 12805 3009 12817 3012
rect 12851 3040 12863 3043
rect 12894 3040 12900 3052
rect 12851 3012 12900 3040
rect 12851 3009 12863 3012
rect 12805 3003 12863 3009
rect 12894 3000 12900 3012
rect 12952 3000 12958 3052
rect 13072 3043 13130 3049
rect 13072 3009 13084 3043
rect 13118 3040 13130 3043
rect 13354 3040 13360 3052
rect 13118 3012 13360 3040
rect 13118 3009 13130 3012
rect 13072 3003 13130 3009
rect 13354 3000 13360 3012
rect 13412 3000 13418 3052
rect 11517 2975 11575 2981
rect 11517 2972 11529 2975
rect 10704 2944 11529 2972
rect 8757 2935 8815 2941
rect 11517 2941 11529 2944
rect 11563 2941 11575 2975
rect 11517 2935 11575 2941
rect 11977 2975 12035 2981
rect 11977 2941 11989 2975
rect 12023 2941 12035 2975
rect 11977 2935 12035 2941
rect 5813 2907 5871 2913
rect 5813 2873 5825 2907
rect 5859 2904 5871 2907
rect 6178 2904 6184 2916
rect 5859 2876 6184 2904
rect 5859 2873 5871 2876
rect 5813 2867 5871 2873
rect 6178 2864 6184 2876
rect 6236 2904 6242 2916
rect 6454 2904 6460 2916
rect 6236 2876 6460 2904
rect 6236 2864 6242 2876
rect 6454 2864 6460 2876
rect 6512 2864 6518 2916
rect 7377 2907 7435 2913
rect 7377 2904 7389 2907
rect 7024 2876 7389 2904
rect 4856 2808 5488 2836
rect 5997 2839 6055 2845
rect 4856 2796 4862 2808
rect 5997 2805 6009 2839
rect 6043 2836 6055 2839
rect 7024 2836 7052 2876
rect 7377 2873 7389 2876
rect 7423 2873 7435 2907
rect 7558 2904 7564 2916
rect 7519 2876 7564 2904
rect 7377 2867 7435 2873
rect 7558 2864 7564 2876
rect 7616 2864 7622 2916
rect 8772 2904 8800 2935
rect 10962 2904 10968 2916
rect 8128 2876 8800 2904
rect 10923 2876 10968 2904
rect 8128 2848 8156 2876
rect 10962 2864 10968 2876
rect 11020 2864 11026 2916
rect 11054 2864 11060 2916
rect 11112 2904 11118 2916
rect 11992 2904 12020 2935
rect 11112 2876 12020 2904
rect 13832 2904 13860 3080
rect 14366 3068 14372 3120
rect 14424 3108 14430 3120
rect 15654 3108 15660 3120
rect 14424 3080 15148 3108
rect 14424 3068 14430 3080
rect 14274 3000 14280 3052
rect 14332 3040 14338 3052
rect 15120 3049 15148 3080
rect 15304 3080 15660 3108
rect 15304 3049 15332 3080
rect 15654 3068 15660 3080
rect 15712 3108 15718 3120
rect 16114 3108 16120 3120
rect 15712 3080 16120 3108
rect 15712 3068 15718 3080
rect 16114 3068 16120 3080
rect 16172 3068 16178 3120
rect 16482 3068 16488 3120
rect 16540 3108 16546 3120
rect 20548 3108 20576 3148
rect 28721 3145 28733 3148
rect 28767 3145 28779 3179
rect 30742 3176 30748 3188
rect 30703 3148 30748 3176
rect 28721 3139 28779 3145
rect 30742 3136 30748 3148
rect 30800 3176 30806 3188
rect 31110 3176 31116 3188
rect 30800 3148 31116 3176
rect 30800 3136 30806 3148
rect 31110 3136 31116 3148
rect 31168 3136 31174 3188
rect 16540 3080 20576 3108
rect 16540 3068 16546 3080
rect 25222 3068 25228 3120
rect 25280 3108 25286 3120
rect 28258 3108 28264 3120
rect 25280 3080 25820 3108
rect 25280 3068 25286 3080
rect 14829 3043 14887 3049
rect 14829 3040 14841 3043
rect 14332 3012 14841 3040
rect 14332 3000 14338 3012
rect 14829 3009 14841 3012
rect 14875 3009 14887 3043
rect 14829 3003 14887 3009
rect 15105 3043 15163 3049
rect 15105 3009 15117 3043
rect 15151 3009 15163 3043
rect 15105 3003 15163 3009
rect 15289 3043 15347 3049
rect 15289 3009 15301 3043
rect 15335 3009 15347 3043
rect 15746 3040 15752 3052
rect 15707 3012 15752 3040
rect 15289 3003 15347 3009
rect 15746 3000 15752 3012
rect 15804 3000 15810 3052
rect 15933 3043 15991 3049
rect 15933 3009 15945 3043
rect 15979 3009 15991 3043
rect 16850 3040 16856 3052
rect 16811 3012 16856 3040
rect 15933 3003 15991 3009
rect 14182 2932 14188 2984
rect 14240 2972 14246 2984
rect 15948 2972 15976 3003
rect 16850 3000 16856 3012
rect 16908 3000 16914 3052
rect 17126 3040 17132 3052
rect 17087 3012 17132 3040
rect 17126 3000 17132 3012
rect 17184 3000 17190 3052
rect 17310 3040 17316 3052
rect 17271 3012 17316 3040
rect 17310 3000 17316 3012
rect 17368 3000 17374 3052
rect 18049 3043 18107 3049
rect 18049 3009 18061 3043
rect 18095 3040 18107 3043
rect 18325 3043 18383 3049
rect 18325 3040 18337 3043
rect 18095 3012 18337 3040
rect 18095 3009 18107 3012
rect 18049 3003 18107 3009
rect 18325 3009 18337 3012
rect 18371 3009 18383 3043
rect 18598 3040 18604 3052
rect 18559 3012 18604 3040
rect 18325 3003 18383 3009
rect 18598 3000 18604 3012
rect 18656 3000 18662 3052
rect 18785 3043 18843 3049
rect 18785 3009 18797 3043
rect 18831 3040 18843 3043
rect 18877 3043 18935 3049
rect 18877 3040 18889 3043
rect 18831 3012 18889 3040
rect 18831 3009 18843 3012
rect 18785 3003 18843 3009
rect 18877 3009 18889 3012
rect 18923 3009 18935 3043
rect 18877 3003 18935 3009
rect 19705 3043 19763 3049
rect 19705 3009 19717 3043
rect 19751 3040 19763 3043
rect 19794 3040 19800 3052
rect 19751 3012 19800 3040
rect 19751 3009 19763 3012
rect 19705 3003 19763 3009
rect 19794 3000 19800 3012
rect 19852 3000 19858 3052
rect 20254 3000 20260 3052
rect 20312 3040 20318 3052
rect 20625 3043 20683 3049
rect 20625 3040 20637 3043
rect 20312 3012 20637 3040
rect 20312 3000 20318 3012
rect 20625 3009 20637 3012
rect 20671 3009 20683 3043
rect 20898 3040 20904 3052
rect 20859 3012 20904 3040
rect 20625 3003 20683 3009
rect 20898 3000 20904 3012
rect 20956 3000 20962 3052
rect 21085 3043 21143 3049
rect 21085 3009 21097 3043
rect 21131 3040 21143 3043
rect 21177 3043 21235 3049
rect 21177 3040 21189 3043
rect 21131 3012 21189 3040
rect 21131 3009 21143 3012
rect 21085 3003 21143 3009
rect 21177 3009 21189 3012
rect 21223 3009 21235 3043
rect 22278 3040 22284 3052
rect 22239 3012 22284 3040
rect 21177 3003 21235 3009
rect 22278 3000 22284 3012
rect 22336 3000 22342 3052
rect 22554 3040 22560 3052
rect 22515 3012 22560 3040
rect 22554 3000 22560 3012
rect 22612 3000 22618 3052
rect 22741 3043 22799 3049
rect 22741 3009 22753 3043
rect 22787 3040 22799 3043
rect 23014 3040 23020 3052
rect 22787 3012 23020 3040
rect 22787 3009 22799 3012
rect 22741 3003 22799 3009
rect 23014 3000 23020 3012
rect 23072 3000 23078 3052
rect 23106 3000 23112 3052
rect 23164 3040 23170 3052
rect 23201 3043 23259 3049
rect 23201 3040 23213 3043
rect 23164 3012 23213 3040
rect 23164 3000 23170 3012
rect 23201 3009 23213 3012
rect 23247 3009 23259 3043
rect 23201 3003 23259 3009
rect 23290 3000 23296 3052
rect 23348 3040 23354 3052
rect 23457 3043 23515 3049
rect 23457 3040 23469 3043
rect 23348 3012 23469 3040
rect 23348 3000 23354 3012
rect 23457 3009 23469 3012
rect 23503 3009 23515 3043
rect 23457 3003 23515 3009
rect 24486 3000 24492 3052
rect 24544 3040 24550 3052
rect 25038 3040 25044 3052
rect 24544 3012 25044 3040
rect 24544 3000 24550 3012
rect 25038 3000 25044 3012
rect 25096 3040 25102 3052
rect 25792 3049 25820 3080
rect 27632 3080 28264 3108
rect 25501 3043 25559 3049
rect 25501 3040 25513 3043
rect 25096 3012 25513 3040
rect 25096 3000 25102 3012
rect 25501 3009 25513 3012
rect 25547 3009 25559 3043
rect 25501 3003 25559 3009
rect 25777 3043 25835 3049
rect 25777 3009 25789 3043
rect 25823 3009 25835 3043
rect 25777 3003 25835 3009
rect 25866 3000 25872 3052
rect 25924 3040 25930 3052
rect 27632 3049 27660 3080
rect 28258 3068 28264 3080
rect 28316 3068 28322 3120
rect 31202 3108 31208 3120
rect 28920 3080 31208 3108
rect 25961 3043 26019 3049
rect 25961 3040 25973 3043
rect 25924 3012 25973 3040
rect 25924 3000 25930 3012
rect 25961 3009 25973 3012
rect 26007 3009 26019 3043
rect 25961 3003 26019 3009
rect 27617 3043 27675 3049
rect 27617 3009 27629 3043
rect 27663 3009 27675 3043
rect 27617 3003 27675 3009
rect 27893 3043 27951 3049
rect 27893 3009 27905 3043
rect 27939 3009 27951 3043
rect 27893 3003 27951 3009
rect 14240 2944 15976 2972
rect 14240 2932 14246 2944
rect 16942 2932 16948 2984
rect 17000 2972 17006 2984
rect 18966 2972 18972 2984
rect 17000 2944 18972 2972
rect 17000 2932 17006 2944
rect 18966 2932 18972 2944
rect 19024 2932 19030 2984
rect 19981 2975 20039 2981
rect 19981 2941 19993 2975
rect 20027 2972 20039 2975
rect 27908 2972 27936 3003
rect 27982 3000 27988 3052
rect 28040 3040 28046 3052
rect 28920 3049 28948 3080
rect 31202 3068 31208 3080
rect 31260 3068 31266 3120
rect 28077 3043 28135 3049
rect 28077 3040 28089 3043
rect 28040 3012 28089 3040
rect 28040 3000 28046 3012
rect 28077 3009 28089 3012
rect 28123 3009 28135 3043
rect 28077 3003 28135 3009
rect 28905 3043 28963 3049
rect 28905 3009 28917 3043
rect 28951 3009 28963 3043
rect 28905 3003 28963 3009
rect 29632 3043 29690 3049
rect 29632 3009 29644 3043
rect 29678 3040 29690 3043
rect 30650 3040 30656 3052
rect 29678 3012 30656 3040
rect 29678 3009 29690 3012
rect 29632 3003 29690 3009
rect 30650 3000 30656 3012
rect 30708 3000 30714 3052
rect 28534 2972 28540 2984
rect 20027 2944 21864 2972
rect 27908 2944 28540 2972
rect 20027 2941 20039 2944
rect 19981 2935 20039 2941
rect 13832 2876 16804 2904
rect 11112 2864 11118 2876
rect 6043 2808 7052 2836
rect 6043 2805 6055 2808
rect 5997 2799 6055 2805
rect 7098 2796 7104 2848
rect 7156 2836 7162 2848
rect 8110 2836 8116 2848
rect 7156 2808 8116 2836
rect 7156 2796 7162 2808
rect 8110 2796 8116 2808
rect 8168 2796 8174 2848
rect 11149 2839 11207 2845
rect 11149 2805 11161 2839
rect 11195 2836 11207 2839
rect 11885 2839 11943 2845
rect 11885 2836 11897 2839
rect 11195 2808 11897 2836
rect 11195 2805 11207 2808
rect 11149 2799 11207 2805
rect 11885 2805 11897 2808
rect 11931 2805 11943 2839
rect 11885 2799 11943 2805
rect 14645 2839 14703 2845
rect 14645 2805 14657 2839
rect 14691 2836 14703 2839
rect 14918 2836 14924 2848
rect 14691 2808 14924 2836
rect 14691 2805 14703 2808
rect 14645 2799 14703 2805
rect 14918 2796 14924 2808
rect 14976 2796 14982 2848
rect 15838 2796 15844 2848
rect 15896 2836 15902 2848
rect 16669 2839 16727 2845
rect 16669 2836 16681 2839
rect 15896 2808 16681 2836
rect 15896 2796 15902 2808
rect 16669 2805 16681 2808
rect 16715 2805 16727 2839
rect 16776 2836 16804 2876
rect 16850 2864 16856 2916
rect 16908 2904 16914 2916
rect 17862 2904 17868 2916
rect 16908 2876 17868 2904
rect 16908 2864 16914 2876
rect 17862 2864 17868 2876
rect 17920 2904 17926 2916
rect 18049 2907 18107 2913
rect 18049 2904 18061 2907
rect 17920 2876 18061 2904
rect 17920 2864 17926 2876
rect 18049 2873 18061 2876
rect 18095 2873 18107 2907
rect 18049 2867 18107 2873
rect 19889 2907 19947 2913
rect 19889 2873 19901 2907
rect 19935 2904 19947 2907
rect 21266 2904 21272 2916
rect 19935 2876 21272 2904
rect 19935 2873 19947 2876
rect 19889 2867 19947 2873
rect 21266 2864 21272 2876
rect 21324 2864 21330 2916
rect 21836 2904 21864 2944
rect 28534 2932 28540 2944
rect 28592 2932 28598 2984
rect 28718 2932 28724 2984
rect 28776 2972 28782 2984
rect 29365 2975 29423 2981
rect 29365 2972 29377 2975
rect 28776 2944 29377 2972
rect 28776 2932 28782 2944
rect 28920 2916 28948 2944
rect 29365 2941 29377 2944
rect 29411 2941 29423 2975
rect 29365 2935 29423 2941
rect 23014 2904 23020 2916
rect 21836 2876 23020 2904
rect 23014 2864 23020 2876
rect 23072 2864 23078 2916
rect 24578 2904 24584 2916
rect 24539 2876 24584 2904
rect 24578 2864 24584 2876
rect 24636 2864 24642 2916
rect 28902 2864 28908 2916
rect 28960 2864 28966 2916
rect 17770 2836 17776 2848
rect 16776 2808 17776 2836
rect 16669 2799 16727 2805
rect 17770 2796 17776 2808
rect 17828 2796 17834 2848
rect 18141 2839 18199 2845
rect 18141 2805 18153 2839
rect 18187 2836 18199 2839
rect 18230 2836 18236 2848
rect 18187 2808 18236 2836
rect 18187 2805 18199 2808
rect 18141 2799 18199 2805
rect 18230 2796 18236 2808
rect 18288 2796 18294 2848
rect 19521 2839 19579 2845
rect 19521 2805 19533 2839
rect 19567 2836 19579 2839
rect 19794 2836 19800 2848
rect 19567 2808 19800 2836
rect 19567 2805 19579 2808
rect 19521 2799 19579 2805
rect 19794 2796 19800 2808
rect 19852 2796 19858 2848
rect 20438 2796 20444 2848
rect 20496 2836 20502 2848
rect 21177 2839 21235 2845
rect 21177 2836 21189 2839
rect 20496 2808 21189 2836
rect 20496 2796 20502 2808
rect 21177 2805 21189 2808
rect 21223 2805 21235 2839
rect 21177 2799 21235 2805
rect 22097 2839 22155 2845
rect 22097 2805 22109 2839
rect 22143 2836 22155 2839
rect 22646 2836 22652 2848
rect 22143 2808 22652 2836
rect 22143 2805 22155 2808
rect 22097 2799 22155 2805
rect 22646 2796 22652 2808
rect 22704 2796 22710 2848
rect 25314 2836 25320 2848
rect 25275 2808 25320 2836
rect 25314 2796 25320 2808
rect 25372 2796 25378 2848
rect 26142 2796 26148 2848
rect 26200 2836 26206 2848
rect 27433 2839 27491 2845
rect 27433 2836 27445 2839
rect 26200 2808 27445 2836
rect 26200 2796 26206 2808
rect 27433 2805 27445 2808
rect 27479 2805 27491 2839
rect 27433 2799 27491 2805
rect 1104 2746 32016 2768
rect 0 2700 800 2714
rect 0 2672 888 2700
rect 1104 2694 2136 2746
rect 2188 2694 12440 2746
rect 12492 2694 22744 2746
rect 22796 2694 32016 2746
rect 32320 2700 33120 2714
rect 1104 2672 32016 2694
rect 32048 2672 33120 2700
rect 0 2658 800 2672
rect 860 2496 888 2672
rect 2590 2592 2596 2644
rect 2648 2632 2654 2644
rect 2961 2635 3019 2641
rect 2961 2632 2973 2635
rect 2648 2604 2973 2632
rect 2648 2592 2654 2604
rect 2961 2601 2973 2604
rect 3007 2601 3019 2635
rect 4154 2632 4160 2644
rect 2961 2595 3019 2601
rect 3804 2604 4160 2632
rect 768 2468 888 2496
rect 768 2020 796 2468
rect 1394 2456 1400 2508
rect 1452 2496 1458 2508
rect 3804 2505 3832 2604
rect 4154 2592 4160 2604
rect 4212 2592 4218 2644
rect 4522 2592 4528 2644
rect 4580 2632 4586 2644
rect 5169 2635 5227 2641
rect 5169 2632 5181 2635
rect 4580 2604 5181 2632
rect 4580 2592 4586 2604
rect 5169 2601 5181 2604
rect 5215 2601 5227 2635
rect 5169 2595 5227 2601
rect 6365 2635 6423 2641
rect 6365 2601 6377 2635
rect 6411 2632 6423 2635
rect 8938 2632 8944 2644
rect 6411 2604 8944 2632
rect 6411 2601 6423 2604
rect 6365 2595 6423 2601
rect 8938 2592 8944 2604
rect 8996 2592 9002 2644
rect 9858 2592 9864 2644
rect 9916 2592 9922 2644
rect 10686 2592 10692 2644
rect 10744 2632 10750 2644
rect 10965 2635 11023 2641
rect 10965 2632 10977 2635
rect 10744 2604 10977 2632
rect 10744 2592 10750 2604
rect 10965 2601 10977 2604
rect 11011 2601 11023 2635
rect 10965 2595 11023 2601
rect 12897 2635 12955 2641
rect 12897 2601 12909 2635
rect 12943 2632 12955 2635
rect 13078 2632 13084 2644
rect 12943 2604 13084 2632
rect 12943 2601 12955 2604
rect 12897 2595 12955 2601
rect 13078 2592 13084 2604
rect 13136 2592 13142 2644
rect 13357 2635 13415 2641
rect 13357 2601 13369 2635
rect 13403 2632 13415 2635
rect 14274 2632 14280 2644
rect 13403 2604 14280 2632
rect 13403 2601 13415 2604
rect 13357 2595 13415 2601
rect 14274 2592 14280 2604
rect 14332 2592 14338 2644
rect 16206 2592 16212 2644
rect 16264 2632 16270 2644
rect 16264 2604 18644 2632
rect 16264 2592 16270 2604
rect 9876 2564 9904 2592
rect 10321 2567 10379 2573
rect 10321 2564 10333 2567
rect 9876 2536 10333 2564
rect 10321 2533 10333 2536
rect 10367 2564 10379 2567
rect 10870 2564 10876 2576
rect 10367 2536 10876 2564
rect 10367 2533 10379 2536
rect 10321 2527 10379 2533
rect 10870 2524 10876 2536
rect 10928 2524 10934 2576
rect 18616 2564 18644 2604
rect 18690 2592 18696 2644
rect 18748 2632 18754 2644
rect 20625 2635 20683 2641
rect 20625 2632 20637 2635
rect 18748 2604 20637 2632
rect 18748 2592 18754 2604
rect 20625 2601 20637 2604
rect 20671 2601 20683 2635
rect 20625 2595 20683 2601
rect 22741 2635 22799 2641
rect 22741 2601 22753 2635
rect 22787 2632 22799 2635
rect 22830 2632 22836 2644
rect 22787 2604 22836 2632
rect 22787 2601 22799 2604
rect 22741 2595 22799 2601
rect 22830 2592 22836 2604
rect 22888 2592 22894 2644
rect 24397 2635 24455 2641
rect 24397 2601 24409 2635
rect 24443 2632 24455 2635
rect 25222 2632 25228 2644
rect 24443 2604 25228 2632
rect 24443 2601 24455 2604
rect 24397 2595 24455 2601
rect 25222 2592 25228 2604
rect 25280 2592 25286 2644
rect 27338 2592 27344 2644
rect 27396 2632 27402 2644
rect 28905 2635 28963 2641
rect 28905 2632 28917 2635
rect 27396 2604 28917 2632
rect 27396 2592 27402 2604
rect 28905 2601 28917 2604
rect 28951 2601 28963 2635
rect 28905 2595 28963 2601
rect 29086 2592 29092 2644
rect 29144 2632 29150 2644
rect 30650 2632 30656 2644
rect 29144 2604 30420 2632
rect 30611 2604 30656 2632
rect 29144 2592 29150 2604
rect 19242 2564 19248 2576
rect 18616 2536 19248 2564
rect 19242 2524 19248 2536
rect 19300 2524 19306 2576
rect 24486 2564 24492 2576
rect 23400 2536 24492 2564
rect 1581 2499 1639 2505
rect 1581 2496 1593 2499
rect 1452 2468 1593 2496
rect 1452 2456 1458 2468
rect 1581 2465 1593 2468
rect 1627 2465 1639 2499
rect 1581 2459 1639 2465
rect 3789 2499 3847 2505
rect 3789 2465 3801 2499
rect 3835 2465 3847 2499
rect 7837 2499 7895 2505
rect 7837 2496 7849 2499
rect 3789 2459 3847 2465
rect 7116 2468 7849 2496
rect 937 2431 995 2437
rect 937 2397 949 2431
rect 983 2428 995 2431
rect 5629 2431 5687 2437
rect 5629 2428 5641 2431
rect 983 2400 5641 2428
rect 983 2397 995 2400
rect 937 2391 995 2397
rect 5629 2397 5641 2400
rect 5675 2397 5687 2431
rect 5629 2391 5687 2397
rect 6546 2388 6552 2440
rect 6604 2428 6610 2440
rect 6641 2431 6699 2437
rect 6641 2428 6653 2431
rect 6604 2400 6653 2428
rect 6604 2388 6610 2400
rect 6641 2397 6653 2400
rect 6687 2397 6699 2431
rect 6641 2391 6699 2397
rect 6730 2388 6736 2440
rect 6788 2428 6794 2440
rect 7116 2437 7144 2468
rect 7837 2465 7849 2468
rect 7883 2496 7895 2499
rect 8110 2496 8116 2508
rect 7883 2468 8116 2496
rect 7883 2465 7895 2468
rect 7837 2459 7895 2465
rect 8110 2456 8116 2468
rect 8168 2456 8174 2508
rect 11330 2456 11336 2508
rect 11388 2496 11394 2508
rect 11517 2499 11575 2505
rect 11517 2496 11529 2499
rect 11388 2468 11529 2496
rect 11388 2456 11394 2468
rect 11517 2465 11529 2468
rect 11563 2465 11575 2499
rect 11517 2459 11575 2465
rect 12802 2456 12808 2508
rect 12860 2496 12866 2508
rect 14550 2496 14556 2508
rect 12860 2468 14556 2496
rect 12860 2456 12866 2468
rect 14550 2456 14556 2468
rect 14608 2456 14614 2508
rect 18693 2499 18751 2505
rect 18693 2465 18705 2499
rect 18739 2496 18751 2499
rect 18782 2496 18788 2508
rect 18739 2468 18788 2496
rect 18739 2465 18751 2468
rect 18693 2459 18751 2465
rect 18782 2456 18788 2468
rect 18840 2456 18846 2508
rect 6917 2431 6975 2437
rect 6917 2428 6929 2431
rect 6788 2400 6929 2428
rect 6788 2388 6794 2400
rect 6917 2397 6929 2400
rect 6963 2397 6975 2431
rect 6917 2391 6975 2397
rect 7101 2431 7159 2437
rect 7101 2397 7113 2431
rect 7147 2397 7159 2431
rect 7558 2428 7564 2440
rect 7519 2400 7564 2428
rect 7101 2391 7159 2397
rect 7558 2388 7564 2400
rect 7616 2388 7622 2440
rect 8941 2431 8999 2437
rect 8941 2397 8953 2431
rect 8987 2428 8999 2431
rect 9582 2428 9588 2440
rect 8987 2400 9588 2428
rect 8987 2397 8999 2400
rect 8941 2391 8999 2397
rect 9582 2388 9588 2400
rect 9640 2388 9646 2440
rect 10502 2388 10508 2440
rect 10560 2428 10566 2440
rect 10873 2431 10931 2437
rect 10873 2428 10885 2431
rect 10560 2400 10885 2428
rect 10560 2388 10566 2400
rect 10873 2397 10885 2400
rect 10919 2397 10931 2431
rect 10873 2391 10931 2397
rect 13541 2431 13599 2437
rect 13541 2397 13553 2431
rect 13587 2428 13599 2431
rect 16206 2428 16212 2440
rect 13587 2400 16212 2428
rect 13587 2397 13599 2400
rect 13541 2391 13599 2397
rect 16206 2388 16212 2400
rect 16264 2388 16270 2440
rect 16393 2431 16451 2437
rect 16393 2397 16405 2431
rect 16439 2428 16451 2431
rect 18138 2428 18144 2440
rect 16439 2400 18144 2428
rect 16439 2397 16451 2400
rect 16393 2391 16451 2397
rect 18138 2388 18144 2400
rect 18196 2388 18202 2440
rect 18414 2428 18420 2440
rect 18375 2400 18420 2428
rect 18414 2388 18420 2400
rect 18472 2388 18478 2440
rect 18598 2428 18604 2440
rect 18559 2400 18604 2428
rect 18598 2388 18604 2400
rect 18656 2388 18662 2440
rect 19245 2431 19303 2437
rect 19245 2397 19257 2431
rect 19291 2428 19303 2431
rect 21361 2431 21419 2437
rect 21361 2428 21373 2431
rect 19291 2400 21373 2428
rect 19291 2397 19303 2400
rect 19245 2391 19303 2397
rect 21361 2397 21373 2400
rect 21407 2428 21419 2431
rect 21910 2428 21916 2440
rect 21407 2400 21916 2428
rect 21407 2397 21419 2400
rect 21361 2391 21419 2397
rect 21910 2388 21916 2400
rect 21968 2428 21974 2440
rect 23106 2428 23112 2440
rect 21968 2400 23112 2428
rect 21968 2388 21974 2400
rect 23106 2388 23112 2400
rect 23164 2388 23170 2440
rect 23400 2437 23428 2536
rect 24486 2524 24492 2536
rect 24544 2524 24550 2576
rect 28350 2524 28356 2576
rect 28408 2564 28414 2576
rect 30285 2567 30343 2573
rect 30285 2564 30297 2567
rect 28408 2536 30297 2564
rect 28408 2524 28414 2536
rect 30285 2533 30297 2536
rect 30331 2533 30343 2567
rect 30392 2564 30420 2604
rect 30650 2592 30656 2604
rect 30708 2592 30714 2644
rect 32048 2564 32076 2672
rect 32320 2658 33120 2672
rect 30392 2536 32076 2564
rect 30285 2527 30343 2533
rect 24397 2499 24455 2505
rect 24397 2496 24409 2499
rect 23676 2468 24409 2496
rect 23676 2437 23704 2468
rect 24397 2465 24409 2468
rect 24443 2465 24455 2499
rect 24397 2459 24455 2465
rect 28368 2468 29500 2496
rect 23385 2431 23443 2437
rect 23385 2397 23397 2431
rect 23431 2397 23443 2431
rect 23385 2391 23443 2397
rect 23661 2431 23719 2437
rect 23661 2397 23673 2431
rect 23707 2397 23719 2431
rect 23661 2391 23719 2397
rect 23845 2431 23903 2437
rect 23845 2397 23857 2431
rect 23891 2397 23903 2431
rect 23845 2391 23903 2397
rect 1848 2363 1906 2369
rect 1848 2329 1860 2363
rect 1894 2360 1906 2363
rect 2038 2360 2044 2372
rect 1894 2332 2044 2360
rect 1894 2329 1906 2332
rect 1848 2323 1906 2329
rect 2038 2320 2044 2332
rect 2096 2320 2102 2372
rect 3142 2320 3148 2372
rect 3200 2360 3206 2372
rect 4034 2363 4092 2369
rect 4034 2360 4046 2363
rect 3200 2332 4046 2360
rect 3200 2320 3206 2332
rect 4034 2329 4046 2332
rect 4080 2329 4092 2363
rect 9208 2363 9266 2369
rect 4034 2323 4092 2329
rect 4264 2332 7512 2360
rect 3510 2252 3516 2304
rect 3568 2292 3574 2304
rect 4264 2292 4292 2332
rect 3568 2264 4292 2292
rect 3568 2252 3574 2264
rect 4430 2252 4436 2304
rect 4488 2292 4494 2304
rect 5813 2295 5871 2301
rect 5813 2292 5825 2295
rect 4488 2264 5825 2292
rect 4488 2252 4494 2264
rect 5813 2261 5825 2264
rect 5859 2292 5871 2295
rect 6365 2295 6423 2301
rect 6365 2292 6377 2295
rect 5859 2264 6377 2292
rect 5859 2261 5871 2264
rect 5813 2255 5871 2261
rect 6365 2261 6377 2264
rect 6411 2261 6423 2295
rect 6365 2255 6423 2261
rect 6457 2295 6515 2301
rect 6457 2261 6469 2295
rect 6503 2292 6515 2295
rect 7374 2292 7380 2304
rect 6503 2264 7380 2292
rect 6503 2261 6515 2264
rect 6457 2255 6515 2261
rect 7374 2252 7380 2264
rect 7432 2252 7438 2304
rect 7484 2292 7512 2332
rect 9208 2329 9220 2363
rect 9254 2360 9266 2363
rect 10226 2360 10232 2372
rect 9254 2332 10232 2360
rect 9254 2329 9266 2332
rect 9208 2323 9266 2329
rect 10226 2320 10232 2332
rect 10284 2320 10290 2372
rect 11784 2363 11842 2369
rect 11784 2329 11796 2363
rect 11830 2360 11842 2363
rect 13078 2360 13084 2372
rect 11830 2332 13084 2360
rect 11830 2329 11842 2332
rect 11784 2323 11842 2329
rect 13078 2320 13084 2332
rect 13136 2320 13142 2372
rect 14820 2363 14878 2369
rect 14820 2329 14832 2363
rect 14866 2360 14878 2363
rect 15654 2360 15660 2372
rect 14866 2332 15660 2360
rect 14866 2329 14878 2332
rect 14820 2323 14878 2329
rect 15654 2320 15660 2332
rect 15712 2320 15718 2372
rect 16666 2369 16672 2372
rect 16660 2323 16672 2369
rect 16724 2360 16730 2372
rect 18233 2363 18291 2369
rect 16724 2332 16760 2360
rect 16666 2320 16672 2323
rect 16724 2320 16730 2332
rect 18233 2329 18245 2363
rect 18279 2360 18291 2363
rect 19490 2363 19548 2369
rect 19490 2360 19502 2363
rect 18279 2332 19502 2360
rect 18279 2329 18291 2332
rect 18233 2323 18291 2329
rect 19490 2329 19502 2332
rect 19536 2329 19548 2363
rect 19490 2323 19548 2329
rect 19794 2320 19800 2372
rect 19852 2360 19858 2372
rect 21606 2363 21664 2369
rect 21606 2360 21618 2363
rect 19852 2332 21618 2360
rect 19852 2320 19858 2332
rect 21606 2329 21618 2332
rect 21652 2329 21664 2363
rect 21606 2323 21664 2329
rect 22922 2320 22928 2372
rect 22980 2360 22986 2372
rect 23860 2360 23888 2391
rect 24026 2388 24032 2440
rect 24084 2428 24090 2440
rect 24489 2431 24547 2437
rect 24489 2428 24501 2431
rect 24084 2400 24501 2428
rect 24084 2388 24090 2400
rect 24489 2397 24501 2400
rect 24535 2428 24547 2431
rect 26329 2431 26387 2437
rect 26329 2428 26341 2431
rect 24535 2400 26341 2428
rect 24535 2397 24547 2400
rect 24489 2391 24547 2397
rect 26329 2397 26341 2400
rect 26375 2428 26387 2431
rect 27614 2428 27620 2440
rect 26375 2400 27620 2428
rect 26375 2397 26387 2400
rect 26329 2391 26387 2397
rect 27614 2388 27620 2400
rect 27672 2388 27678 2440
rect 28258 2388 28264 2440
rect 28316 2428 28322 2440
rect 28368 2437 28396 2468
rect 28353 2431 28411 2437
rect 28353 2428 28365 2431
rect 28316 2400 28365 2428
rect 28316 2388 28322 2400
rect 28353 2397 28365 2400
rect 28399 2397 28411 2431
rect 28353 2391 28411 2397
rect 28534 2388 28540 2440
rect 28592 2428 28598 2440
rect 28629 2431 28687 2437
rect 28629 2428 28641 2431
rect 28592 2400 28641 2428
rect 28592 2388 28598 2400
rect 28629 2397 28641 2400
rect 28675 2397 28687 2431
rect 28629 2391 28687 2397
rect 24578 2360 24584 2372
rect 22980 2332 24584 2360
rect 22980 2320 22986 2332
rect 24578 2320 24584 2332
rect 24636 2320 24642 2372
rect 24756 2363 24814 2369
rect 24756 2329 24768 2363
rect 24802 2360 24814 2363
rect 25774 2360 25780 2372
rect 24802 2332 25780 2360
rect 24802 2329 24814 2332
rect 24756 2323 24814 2329
rect 25774 2320 25780 2332
rect 25832 2320 25838 2372
rect 25958 2320 25964 2372
rect 26016 2360 26022 2372
rect 26574 2363 26632 2369
rect 26574 2360 26586 2363
rect 26016 2332 26586 2360
rect 26016 2320 26022 2332
rect 26574 2329 26586 2332
rect 26620 2329 26632 2363
rect 28644 2360 28672 2391
rect 28810 2388 28816 2440
rect 28868 2428 28874 2440
rect 28905 2431 28963 2437
rect 28905 2428 28917 2431
rect 28868 2400 28917 2428
rect 28868 2388 28874 2400
rect 28905 2397 28917 2400
rect 28951 2397 28963 2431
rect 29472 2428 29500 2468
rect 30098 2456 30104 2508
rect 30156 2496 30162 2508
rect 31113 2499 31171 2505
rect 31113 2496 31125 2499
rect 30156 2468 31125 2496
rect 30156 2456 30162 2468
rect 31113 2465 31125 2468
rect 31159 2465 31171 2499
rect 31113 2459 31171 2465
rect 29730 2437 29736 2440
rect 29726 2428 29736 2437
rect 29472 2400 29736 2428
rect 28905 2391 28963 2397
rect 29726 2391 29736 2400
rect 29730 2388 29736 2391
rect 29788 2388 29794 2440
rect 30006 2428 30012 2440
rect 29919 2400 30012 2428
rect 30006 2388 30012 2400
rect 30064 2388 30070 2440
rect 30193 2431 30251 2437
rect 30193 2397 30205 2431
rect 30239 2428 30251 2431
rect 30282 2428 30288 2440
rect 30239 2400 30288 2428
rect 30239 2397 30251 2400
rect 30193 2391 30251 2397
rect 30282 2388 30288 2400
rect 30340 2388 30346 2440
rect 30558 2388 30564 2440
rect 30616 2428 30622 2440
rect 30837 2431 30895 2437
rect 30837 2428 30849 2431
rect 30616 2400 30849 2428
rect 30616 2388 30622 2400
rect 30837 2397 30849 2400
rect 30883 2397 30895 2431
rect 31018 2428 31024 2440
rect 30979 2400 31024 2428
rect 30837 2391 30895 2397
rect 31018 2388 31024 2400
rect 31076 2388 31082 2440
rect 30024 2360 30052 2388
rect 28644 2332 30052 2360
rect 26574 2323 26632 2329
rect 11054 2292 11060 2304
rect 7484 2264 11060 2292
rect 11054 2252 11060 2264
rect 11112 2252 11118 2304
rect 12066 2252 12072 2304
rect 12124 2292 12130 2304
rect 14090 2292 14096 2304
rect 12124 2264 14096 2292
rect 12124 2252 12130 2264
rect 14090 2252 14096 2264
rect 14148 2252 14154 2304
rect 15930 2292 15936 2304
rect 15891 2264 15936 2292
rect 15930 2252 15936 2264
rect 15988 2292 15994 2304
rect 17034 2292 17040 2304
rect 15988 2264 17040 2292
rect 15988 2252 15994 2264
rect 17034 2252 17040 2264
rect 17092 2292 17098 2304
rect 17310 2292 17316 2304
rect 17092 2264 17316 2292
rect 17092 2252 17098 2264
rect 17310 2252 17316 2264
rect 17368 2252 17374 2304
rect 17770 2292 17776 2304
rect 17731 2264 17776 2292
rect 17770 2252 17776 2264
rect 17828 2252 17834 2304
rect 17862 2252 17868 2304
rect 17920 2292 17926 2304
rect 21450 2292 21456 2304
rect 17920 2264 21456 2292
rect 17920 2252 17926 2264
rect 21450 2252 21456 2264
rect 21508 2252 21514 2304
rect 23201 2295 23259 2301
rect 23201 2261 23213 2295
rect 23247 2292 23259 2295
rect 23566 2292 23572 2304
rect 23247 2264 23572 2292
rect 23247 2261 23259 2264
rect 23201 2255 23259 2261
rect 23566 2252 23572 2264
rect 23624 2252 23630 2304
rect 25130 2252 25136 2304
rect 25188 2292 25194 2304
rect 25866 2292 25872 2304
rect 25188 2264 25872 2292
rect 25188 2252 25194 2264
rect 25866 2252 25872 2264
rect 25924 2252 25930 2304
rect 26234 2252 26240 2304
rect 26292 2292 26298 2304
rect 27062 2292 27068 2304
rect 26292 2264 27068 2292
rect 26292 2252 26298 2264
rect 27062 2252 27068 2264
rect 27120 2292 27126 2304
rect 27709 2295 27767 2301
rect 27709 2292 27721 2295
rect 27120 2264 27721 2292
rect 27120 2252 27126 2264
rect 27709 2261 27721 2264
rect 27755 2292 27767 2295
rect 27982 2292 27988 2304
rect 27755 2264 27988 2292
rect 27755 2261 27767 2264
rect 27709 2255 27767 2261
rect 27982 2252 27988 2264
rect 28040 2252 28046 2304
rect 28074 2252 28080 2304
rect 28132 2292 28138 2304
rect 28169 2295 28227 2301
rect 28169 2292 28181 2295
rect 28132 2264 28181 2292
rect 28132 2252 28138 2264
rect 28169 2261 28181 2264
rect 28215 2261 28227 2295
rect 28169 2255 28227 2261
rect 29549 2295 29607 2301
rect 29549 2261 29561 2295
rect 29595 2292 29607 2295
rect 30834 2292 30840 2304
rect 29595 2264 30840 2292
rect 29595 2261 29607 2264
rect 29549 2255 29607 2261
rect 30834 2252 30840 2264
rect 30892 2252 30898 2304
rect 1104 2202 32016 2224
rect 1104 2150 7288 2202
rect 7340 2150 17592 2202
rect 17644 2150 27896 2202
rect 27948 2150 32016 2202
rect 1104 2128 32016 2150
rect 2038 2048 2044 2100
rect 2096 2088 2102 2100
rect 2133 2091 2191 2097
rect 2133 2088 2145 2091
rect 2096 2060 2145 2088
rect 2096 2048 2102 2060
rect 2133 2057 2145 2060
rect 2179 2057 2191 2091
rect 3142 2088 3148 2100
rect 3103 2060 3148 2088
rect 2133 2051 2191 2057
rect 3142 2048 3148 2060
rect 3200 2048 3206 2100
rect 5813 2091 5871 2097
rect 5813 2057 5825 2091
rect 5859 2088 5871 2091
rect 6822 2088 6828 2100
rect 5859 2060 6828 2088
rect 5859 2057 5871 2060
rect 5813 2051 5871 2057
rect 6822 2048 6828 2060
rect 6880 2048 6886 2100
rect 7558 2048 7564 2100
rect 7616 2088 7622 2100
rect 8202 2088 8208 2100
rect 7616 2060 8208 2088
rect 7616 2048 7622 2060
rect 8202 2048 8208 2060
rect 8260 2088 8266 2100
rect 8573 2091 8631 2097
rect 8573 2088 8585 2091
rect 8260 2060 8585 2088
rect 8260 2048 8266 2060
rect 8573 2057 8585 2060
rect 8619 2057 8631 2091
rect 8573 2051 8631 2057
rect 10965 2091 11023 2097
rect 10965 2057 10977 2091
rect 11011 2057 11023 2091
rect 10965 2051 11023 2057
rect 4706 2029 4712 2032
rect 1489 2023 1547 2029
rect 1489 2020 1501 2023
rect 768 1992 1501 2020
rect 1489 1989 1501 1992
rect 1535 1989 1547 2023
rect 4700 2020 4712 2029
rect 4667 1992 4712 2020
rect 1489 1983 1547 1989
rect 4700 1983 4712 1992
rect 4706 1980 4712 1983
rect 4764 1980 4770 2032
rect 7006 2020 7012 2032
rect 5460 1992 7012 2020
rect 2314 1952 2320 1964
rect 2275 1924 2320 1952
rect 2314 1912 2320 1924
rect 2372 1912 2378 1964
rect 2501 1955 2559 1961
rect 2501 1921 2513 1955
rect 2547 1952 2559 1955
rect 3326 1952 3332 1964
rect 2547 1924 2820 1952
rect 3287 1924 3332 1952
rect 2547 1921 2559 1924
rect 2501 1915 2559 1921
rect 2593 1887 2651 1893
rect 2593 1853 2605 1887
rect 2639 1884 2651 1887
rect 2682 1884 2688 1896
rect 2639 1856 2688 1884
rect 2639 1853 2651 1856
rect 2593 1847 2651 1853
rect 2682 1844 2688 1856
rect 2740 1844 2746 1896
rect 2792 1884 2820 1924
rect 3326 1912 3332 1924
rect 3384 1912 3390 1964
rect 3605 1955 3663 1961
rect 3605 1921 3617 1955
rect 3651 1952 3663 1955
rect 4062 1952 4068 1964
rect 3651 1924 4068 1952
rect 3651 1921 3663 1924
rect 3605 1915 3663 1921
rect 4062 1912 4068 1924
rect 4120 1912 4126 1964
rect 4154 1912 4160 1964
rect 4212 1952 4218 1964
rect 4433 1955 4491 1961
rect 4433 1952 4445 1955
rect 4212 1924 4445 1952
rect 4212 1912 4218 1924
rect 4433 1921 4445 1924
rect 4479 1921 4491 1955
rect 4433 1915 4491 1921
rect 3050 1884 3056 1896
rect 2792 1856 3056 1884
rect 3050 1844 3056 1856
rect 3108 1884 3114 1896
rect 3513 1887 3571 1893
rect 3513 1884 3525 1887
rect 3108 1856 3525 1884
rect 3108 1844 3114 1856
rect 3513 1853 3525 1856
rect 3559 1853 3571 1887
rect 3513 1847 3571 1853
rect 1581 1751 1639 1757
rect 1581 1717 1593 1751
rect 1627 1748 1639 1751
rect 5460 1748 5488 1992
rect 7006 1980 7012 1992
rect 7064 1980 7070 2032
rect 10980 2020 11008 2051
rect 11054 2048 11060 2100
rect 11112 2088 11118 2100
rect 11112 2060 20024 2088
rect 11112 2048 11118 2060
rect 11762 2023 11820 2029
rect 11762 2020 11774 2023
rect 10980 1992 11774 2020
rect 11762 1989 11774 1992
rect 11808 1989 11820 2023
rect 13354 2020 13360 2032
rect 13315 1992 13360 2020
rect 11762 1983 11820 1989
rect 13354 1980 13360 1992
rect 13412 1980 13418 2032
rect 17862 2020 17868 2032
rect 13648 1992 17868 2020
rect 6733 1955 6791 1961
rect 6733 1921 6745 1955
rect 6779 1921 6791 1955
rect 7190 1952 7196 1964
rect 7151 1924 7196 1952
rect 6733 1915 6791 1921
rect 6546 1748 6552 1760
rect 1627 1720 5488 1748
rect 6507 1720 6552 1748
rect 1627 1717 1639 1720
rect 1581 1711 1639 1717
rect 6546 1708 6552 1720
rect 6604 1708 6610 1760
rect 6748 1748 6776 1915
rect 7190 1912 7196 1924
rect 7248 1912 7254 1964
rect 7466 1961 7472 1964
rect 7460 1915 7472 1961
rect 7524 1952 7530 1964
rect 9582 1952 9588 1964
rect 7524 1924 7560 1952
rect 9543 1924 9588 1952
rect 7466 1912 7472 1915
rect 7524 1912 7530 1924
rect 9582 1912 9588 1924
rect 9640 1912 9646 1964
rect 9674 1912 9680 1964
rect 9732 1952 9738 1964
rect 9841 1955 9899 1961
rect 9841 1952 9853 1955
rect 9732 1924 9853 1952
rect 9732 1912 9738 1924
rect 9841 1921 9853 1924
rect 9887 1921 9899 1955
rect 9841 1915 9899 1921
rect 11330 1912 11336 1964
rect 11388 1952 11394 1964
rect 11517 1955 11575 1961
rect 11517 1952 11529 1955
rect 11388 1924 11529 1952
rect 11388 1912 11394 1924
rect 11517 1921 11529 1924
rect 11563 1921 11575 1955
rect 13538 1952 13544 1964
rect 13499 1924 13544 1952
rect 11517 1915 11575 1921
rect 13538 1912 13544 1924
rect 13596 1912 13602 1964
rect 12894 1816 12900 1828
rect 12855 1788 12900 1816
rect 12894 1776 12900 1788
rect 12952 1776 12958 1828
rect 13648 1816 13676 1992
rect 17862 1980 17868 1992
rect 17920 1980 17926 2032
rect 18138 2020 18144 2032
rect 18051 1992 18144 2020
rect 14550 1952 14556 1964
rect 14511 1924 14556 1952
rect 14550 1912 14556 1924
rect 14608 1912 14614 1964
rect 14826 1961 14832 1964
rect 14820 1915 14832 1961
rect 14884 1952 14890 1964
rect 14884 1924 14920 1952
rect 14826 1912 14832 1915
rect 14884 1912 14890 1924
rect 16850 1912 16856 1964
rect 16908 1952 16914 1964
rect 17037 1955 17095 1961
rect 17037 1952 17049 1955
rect 16908 1924 17049 1952
rect 16908 1912 16914 1924
rect 17037 1921 17049 1924
rect 17083 1921 17095 1955
rect 17037 1915 17095 1921
rect 17126 1912 17132 1964
rect 17184 1952 17190 1964
rect 17313 1955 17371 1961
rect 17313 1952 17325 1955
rect 17184 1924 17325 1952
rect 17184 1912 17190 1924
rect 17313 1921 17325 1924
rect 17359 1921 17371 1955
rect 17313 1915 17371 1921
rect 17497 1955 17555 1961
rect 17497 1921 17509 1955
rect 17543 1952 17555 1955
rect 17770 1952 17776 1964
rect 17543 1924 17776 1952
rect 17543 1921 17555 1924
rect 17497 1915 17555 1921
rect 13817 1887 13875 1893
rect 13817 1853 13829 1887
rect 13863 1853 13875 1887
rect 13817 1847 13875 1853
rect 13464 1788 13676 1816
rect 13464 1748 13492 1788
rect 6748 1720 13492 1748
rect 13538 1708 13544 1760
rect 13596 1748 13602 1760
rect 13725 1751 13783 1757
rect 13725 1748 13737 1751
rect 13596 1720 13737 1748
rect 13596 1708 13602 1720
rect 13725 1717 13737 1720
rect 13771 1717 13783 1751
rect 13832 1748 13860 1847
rect 16574 1844 16580 1896
rect 16632 1884 16638 1896
rect 16758 1884 16764 1896
rect 16632 1856 16764 1884
rect 16632 1844 16638 1856
rect 16758 1844 16764 1856
rect 16816 1884 16822 1896
rect 17512 1884 17540 1915
rect 17770 1912 17776 1924
rect 17828 1912 17834 1964
rect 18064 1961 18092 1992
rect 18138 1980 18144 1992
rect 18196 2020 18202 2032
rect 19996 2020 20024 2060
rect 20622 2048 20628 2100
rect 20680 2088 20686 2100
rect 21269 2091 21327 2097
rect 21269 2088 21281 2091
rect 20680 2060 21281 2088
rect 20680 2048 20686 2060
rect 21269 2057 21281 2060
rect 21315 2057 21327 2091
rect 21269 2051 21327 2057
rect 23014 2048 23020 2100
rect 23072 2088 23078 2100
rect 23293 2091 23351 2097
rect 23293 2088 23305 2091
rect 23072 2060 23305 2088
rect 23072 2048 23078 2060
rect 23293 2057 23305 2060
rect 23339 2057 23351 2091
rect 23293 2051 23351 2057
rect 25409 2091 25467 2097
rect 25409 2057 25421 2091
rect 25455 2088 25467 2091
rect 25590 2088 25596 2100
rect 25455 2060 25596 2088
rect 25455 2057 25467 2060
rect 25409 2051 25467 2057
rect 25590 2048 25596 2060
rect 25648 2048 25654 2100
rect 25958 2088 25964 2100
rect 25919 2060 25964 2088
rect 25958 2048 25964 2060
rect 26016 2048 26022 2100
rect 31113 2091 31171 2097
rect 31113 2088 31125 2091
rect 26620 2060 31125 2088
rect 26620 2020 26648 2060
rect 31113 2057 31125 2060
rect 31159 2057 31171 2091
rect 31113 2051 31171 2057
rect 27614 2020 27620 2032
rect 18196 1992 19932 2020
rect 19996 1992 26648 2020
rect 27448 1992 27620 2020
rect 18196 1980 18202 1992
rect 18322 1961 18328 1964
rect 18049 1955 18107 1961
rect 18049 1921 18061 1955
rect 18095 1921 18107 1955
rect 18049 1915 18107 1921
rect 18316 1915 18328 1961
rect 18380 1952 18386 1964
rect 19904 1961 19932 1992
rect 19889 1955 19947 1961
rect 18380 1924 18416 1952
rect 18322 1912 18328 1915
rect 18380 1912 18386 1924
rect 19889 1921 19901 1955
rect 19935 1921 19947 1955
rect 19889 1915 19947 1921
rect 19978 1912 19984 1964
rect 20036 1952 20042 1964
rect 20145 1955 20203 1961
rect 20145 1952 20157 1955
rect 20036 1924 20157 1952
rect 20036 1912 20042 1924
rect 20145 1921 20157 1924
rect 20191 1921 20203 1955
rect 21910 1952 21916 1964
rect 21871 1924 21916 1952
rect 20145 1915 20203 1921
rect 21910 1912 21916 1924
rect 21968 1912 21974 1964
rect 22180 1955 22238 1961
rect 22180 1921 22192 1955
rect 22226 1952 22238 1955
rect 22462 1952 22468 1964
rect 22226 1924 22468 1952
rect 22226 1921 22238 1924
rect 22180 1915 22238 1921
rect 22462 1912 22468 1924
rect 22520 1912 22526 1964
rect 24026 1952 24032 1964
rect 23987 1924 24032 1952
rect 24026 1912 24032 1924
rect 24084 1912 24090 1964
rect 24296 1955 24354 1961
rect 24296 1921 24308 1955
rect 24342 1952 24354 1955
rect 24670 1952 24676 1964
rect 24342 1924 24676 1952
rect 24342 1921 24354 1924
rect 24296 1915 24354 1921
rect 24670 1912 24676 1924
rect 24728 1912 24734 1964
rect 26142 1952 26148 1964
rect 26103 1924 26148 1952
rect 26142 1912 26148 1924
rect 26200 1912 26206 1964
rect 26326 1952 26332 1964
rect 26287 1924 26332 1952
rect 26326 1912 26332 1924
rect 26384 1912 26390 1964
rect 26421 1955 26479 1961
rect 26421 1921 26433 1955
rect 26467 1952 26479 1955
rect 27338 1952 27344 1964
rect 26467 1924 27344 1952
rect 26467 1921 26479 1924
rect 26421 1915 26479 1921
rect 27338 1912 27344 1924
rect 27396 1912 27402 1964
rect 27448 1961 27476 1992
rect 27614 1980 27620 1992
rect 27672 2020 27678 2032
rect 28902 2020 28908 2032
rect 27672 1992 28908 2020
rect 27672 1980 27678 1992
rect 28902 1980 28908 1992
rect 28960 2020 28966 2032
rect 28960 1992 29316 2020
rect 28960 1980 28966 1992
rect 27706 1961 27712 1964
rect 27433 1955 27491 1961
rect 27433 1921 27445 1955
rect 27479 1921 27491 1955
rect 27433 1915 27491 1921
rect 27700 1915 27712 1961
rect 27764 1952 27770 1964
rect 29288 1961 29316 1992
rect 29273 1955 29331 1961
rect 27764 1924 27800 1952
rect 27706 1912 27712 1915
rect 27764 1912 27770 1924
rect 29273 1921 29285 1955
rect 29319 1921 29331 1955
rect 29273 1915 29331 1921
rect 29540 1955 29598 1961
rect 29540 1921 29552 1955
rect 29586 1952 29598 1955
rect 30650 1952 30656 1964
rect 29586 1924 30656 1952
rect 29586 1921 29598 1924
rect 29540 1915 29598 1921
rect 30650 1912 30656 1924
rect 30708 1912 30714 1964
rect 31294 1952 31300 1964
rect 31255 1924 31300 1952
rect 31294 1912 31300 1924
rect 31352 1912 31358 1964
rect 16816 1856 17540 1884
rect 16816 1844 16822 1856
rect 28810 1816 28816 1828
rect 28771 1788 28816 1816
rect 28810 1776 28816 1788
rect 28868 1776 28874 1828
rect 30282 1776 30288 1828
rect 30340 1816 30346 1828
rect 30653 1819 30711 1825
rect 30653 1816 30665 1819
rect 30340 1788 30665 1816
rect 30340 1776 30346 1788
rect 30653 1785 30665 1788
rect 30699 1785 30711 1819
rect 30653 1779 30711 1785
rect 15746 1748 15752 1760
rect 13832 1720 15752 1748
rect 13725 1711 13783 1717
rect 15746 1708 15752 1720
rect 15804 1748 15810 1760
rect 15933 1751 15991 1757
rect 15933 1748 15945 1751
rect 15804 1720 15945 1748
rect 15804 1708 15810 1720
rect 15933 1717 15945 1720
rect 15979 1717 15991 1751
rect 16850 1748 16856 1760
rect 16811 1720 16856 1748
rect 15933 1711 15991 1717
rect 16850 1708 16856 1720
rect 16908 1708 16914 1760
rect 17678 1708 17684 1760
rect 17736 1748 17742 1760
rect 19429 1751 19487 1757
rect 19429 1748 19441 1751
rect 17736 1720 19441 1748
rect 17736 1708 17742 1720
rect 19429 1717 19441 1720
rect 19475 1717 19487 1751
rect 19429 1711 19487 1717
rect 1104 1658 32016 1680
rect 1104 1606 2136 1658
rect 2188 1606 12440 1658
rect 12492 1606 22744 1658
rect 22796 1606 32016 1658
rect 1104 1584 32016 1606
rect 1854 1504 1860 1556
rect 1912 1544 1918 1556
rect 1949 1547 2007 1553
rect 1949 1544 1961 1547
rect 1912 1516 1961 1544
rect 1912 1504 1918 1516
rect 1949 1513 1961 1516
rect 1995 1513 2007 1547
rect 1949 1507 2007 1513
rect 2685 1547 2743 1553
rect 2685 1513 2697 1547
rect 2731 1544 2743 1547
rect 2866 1544 2872 1556
rect 2731 1516 2872 1544
rect 2731 1513 2743 1516
rect 2685 1507 2743 1513
rect 2866 1504 2872 1516
rect 2924 1504 2930 1556
rect 6270 1504 6276 1556
rect 6328 1544 6334 1556
rect 6365 1547 6423 1553
rect 6365 1544 6377 1547
rect 6328 1516 6377 1544
rect 6328 1504 6334 1516
rect 6365 1513 6377 1516
rect 6411 1513 6423 1547
rect 6365 1507 6423 1513
rect 7285 1547 7343 1553
rect 7285 1513 7297 1547
rect 7331 1544 7343 1547
rect 7466 1544 7472 1556
rect 7331 1516 7472 1544
rect 7331 1513 7343 1516
rect 7285 1507 7343 1513
rect 7466 1504 7472 1516
rect 7524 1504 7530 1556
rect 10226 1544 10232 1556
rect 10187 1516 10232 1544
rect 10226 1504 10232 1516
rect 10284 1504 10290 1556
rect 13078 1544 13084 1556
rect 13039 1516 13084 1544
rect 13078 1504 13084 1516
rect 13136 1504 13142 1556
rect 13449 1547 13507 1553
rect 13449 1513 13461 1547
rect 13495 1544 13507 1547
rect 13538 1544 13544 1556
rect 13495 1516 13544 1544
rect 13495 1513 13507 1516
rect 13449 1507 13507 1513
rect 13538 1504 13544 1516
rect 13596 1544 13602 1556
rect 14369 1547 14427 1553
rect 14369 1544 14381 1547
rect 13596 1516 14381 1544
rect 13596 1504 13602 1516
rect 14369 1513 14381 1516
rect 14415 1513 14427 1547
rect 14369 1507 14427 1513
rect 14737 1547 14795 1553
rect 14737 1513 14749 1547
rect 14783 1544 14795 1547
rect 14826 1544 14832 1556
rect 14783 1516 14832 1544
rect 14783 1513 14795 1516
rect 14737 1507 14795 1513
rect 14826 1504 14832 1516
rect 14884 1504 14890 1556
rect 15654 1544 15660 1556
rect 15615 1516 15660 1544
rect 15654 1504 15660 1516
rect 15712 1504 15718 1556
rect 16666 1544 16672 1556
rect 16627 1516 16672 1544
rect 16666 1504 16672 1516
rect 16724 1504 16730 1556
rect 18233 1547 18291 1553
rect 18233 1513 18245 1547
rect 18279 1544 18291 1547
rect 18322 1544 18328 1556
rect 18279 1516 18328 1544
rect 18279 1513 18291 1516
rect 18233 1507 18291 1513
rect 18322 1504 18328 1516
rect 18380 1504 18386 1556
rect 18598 1544 18604 1556
rect 18559 1516 18604 1544
rect 18598 1504 18604 1516
rect 18656 1504 18662 1556
rect 22462 1544 22468 1556
rect 22423 1516 22468 1544
rect 22462 1504 22468 1516
rect 22520 1504 22526 1556
rect 24670 1544 24676 1556
rect 22848 1516 23980 1544
rect 24631 1516 24676 1544
rect 2958 1436 2964 1488
rect 3016 1476 3022 1488
rect 4801 1479 4859 1485
rect 4801 1476 4813 1479
rect 3016 1448 4813 1476
rect 3016 1436 3022 1448
rect 4801 1445 4813 1448
rect 4847 1445 4859 1479
rect 4801 1439 4859 1445
rect 6546 1436 6552 1488
rect 6604 1476 6610 1488
rect 22848 1476 22876 1516
rect 6604 1448 22876 1476
rect 23952 1476 23980 1516
rect 24670 1504 24676 1516
rect 24728 1504 24734 1556
rect 25774 1544 25780 1556
rect 25735 1516 25780 1544
rect 25774 1504 25780 1516
rect 25832 1504 25838 1556
rect 26145 1547 26203 1553
rect 26145 1513 26157 1547
rect 26191 1544 26203 1547
rect 26326 1544 26332 1556
rect 26191 1516 26332 1544
rect 26191 1513 26203 1516
rect 26145 1507 26203 1513
rect 26326 1504 26332 1516
rect 26384 1504 26390 1556
rect 26436 1516 27660 1544
rect 26436 1476 26464 1516
rect 23952 1448 26464 1476
rect 27249 1479 27307 1485
rect 6604 1436 6610 1448
rect 27249 1445 27261 1479
rect 27295 1476 27307 1479
rect 27525 1479 27583 1485
rect 27525 1476 27537 1479
rect 27295 1448 27537 1476
rect 27295 1445 27307 1448
rect 27249 1439 27307 1445
rect 27525 1445 27537 1448
rect 27571 1445 27583 1479
rect 27632 1476 27660 1516
rect 27706 1504 27712 1556
rect 27764 1544 27770 1556
rect 27893 1547 27951 1553
rect 27893 1544 27905 1547
rect 27764 1516 27905 1544
rect 27764 1504 27770 1516
rect 27893 1513 27905 1516
rect 27939 1513 27951 1547
rect 28810 1544 28816 1556
rect 28771 1516 28816 1544
rect 27893 1507 27951 1513
rect 28810 1504 28816 1516
rect 28868 1504 28874 1556
rect 30650 1544 30656 1556
rect 30611 1516 30656 1544
rect 30650 1504 30656 1516
rect 30708 1504 30714 1556
rect 29638 1476 29644 1488
rect 27632 1448 29644 1476
rect 27525 1439 27583 1445
rect 29638 1436 29644 1448
rect 29696 1436 29702 1488
rect 6822 1408 6828 1420
rect 6783 1380 6828 1408
rect 6822 1368 6828 1380
rect 6880 1368 6886 1420
rect 9950 1368 9956 1420
rect 10008 1408 10014 1420
rect 11517 1411 11575 1417
rect 11517 1408 11529 1411
rect 10008 1380 11529 1408
rect 10008 1368 10014 1380
rect 2498 1340 2504 1352
rect 2459 1312 2504 1340
rect 2498 1300 2504 1312
rect 2556 1300 2562 1352
rect 3878 1340 3884 1352
rect 3839 1312 3884 1340
rect 3878 1300 3884 1312
rect 3936 1300 3942 1352
rect 4617 1343 4675 1349
rect 4617 1309 4629 1343
rect 4663 1340 4675 1343
rect 4890 1340 4896 1352
rect 4663 1312 4896 1340
rect 4663 1309 4675 1312
rect 4617 1303 4675 1309
rect 4890 1300 4896 1312
rect 4948 1300 4954 1352
rect 5810 1340 5816 1352
rect 5771 1312 5816 1340
rect 5810 1300 5816 1312
rect 5868 1300 5874 1352
rect 6362 1300 6368 1352
rect 6420 1340 6426 1352
rect 6549 1343 6607 1349
rect 6549 1340 6561 1343
rect 6420 1312 6561 1340
rect 6420 1300 6426 1312
rect 6549 1309 6561 1312
rect 6595 1309 6607 1343
rect 6549 1303 6607 1309
rect 6733 1343 6791 1349
rect 6733 1309 6745 1343
rect 6779 1309 6791 1343
rect 6733 1303 6791 1309
rect 1857 1275 1915 1281
rect 1857 1272 1869 1275
rect 768 1244 1869 1272
rect 768 1068 796 1244
rect 1857 1241 1869 1244
rect 1903 1241 1915 1275
rect 1857 1235 1915 1241
rect 5718 1232 5724 1284
rect 5776 1272 5782 1284
rect 6748 1272 6776 1303
rect 7374 1300 7380 1352
rect 7432 1340 7438 1352
rect 7469 1343 7527 1349
rect 7469 1340 7481 1343
rect 7432 1312 7481 1340
rect 7432 1300 7438 1312
rect 7469 1309 7481 1312
rect 7515 1309 7527 1343
rect 7469 1303 7527 1309
rect 7653 1343 7711 1349
rect 7653 1309 7665 1343
rect 7699 1309 7711 1343
rect 7653 1303 7711 1309
rect 7745 1343 7803 1349
rect 7745 1309 7757 1343
rect 7791 1340 7803 1343
rect 7834 1340 7840 1352
rect 7791 1312 7840 1340
rect 7791 1309 7803 1312
rect 7745 1303 7803 1309
rect 7668 1272 7696 1303
rect 7834 1300 7840 1312
rect 7892 1300 7898 1352
rect 8386 1340 8392 1352
rect 8347 1312 8392 1340
rect 8386 1300 8392 1312
rect 8444 1300 8450 1352
rect 8941 1343 8999 1349
rect 8941 1309 8953 1343
rect 8987 1309 8999 1343
rect 9214 1340 9220 1352
rect 9175 1312 9220 1340
rect 8941 1303 8999 1309
rect 5776 1244 7696 1272
rect 5776 1232 5782 1244
rect 8294 1232 8300 1284
rect 8352 1272 8358 1284
rect 8956 1272 8984 1303
rect 9214 1300 9220 1312
rect 9272 1300 9278 1352
rect 10042 1300 10048 1352
rect 10100 1340 10106 1352
rect 10413 1343 10471 1349
rect 10413 1340 10425 1343
rect 10100 1312 10425 1340
rect 10100 1300 10106 1312
rect 10413 1309 10425 1312
rect 10459 1309 10471 1343
rect 10594 1340 10600 1352
rect 10555 1312 10600 1340
rect 10413 1303 10471 1309
rect 10594 1300 10600 1312
rect 10652 1300 10658 1352
rect 10704 1349 10732 1380
rect 11517 1377 11529 1380
rect 11563 1377 11575 1411
rect 13814 1408 13820 1420
rect 11517 1371 11575 1377
rect 13556 1380 13820 1408
rect 10689 1343 10747 1349
rect 10689 1309 10701 1343
rect 10735 1309 10747 1343
rect 11698 1340 11704 1352
rect 11659 1312 11704 1340
rect 10689 1303 10747 1309
rect 11698 1300 11704 1312
rect 11756 1300 11762 1352
rect 12529 1343 12587 1349
rect 12529 1309 12541 1343
rect 12575 1340 12587 1343
rect 12989 1343 13047 1349
rect 12989 1340 13001 1343
rect 12575 1312 13001 1340
rect 12575 1309 12587 1312
rect 12529 1303 12587 1309
rect 12989 1309 13001 1312
rect 13035 1309 13047 1343
rect 13262 1340 13268 1352
rect 13223 1312 13268 1340
rect 12989 1303 13047 1309
rect 13262 1300 13268 1312
rect 13320 1300 13326 1352
rect 13556 1349 13584 1380
rect 13814 1368 13820 1380
rect 13872 1368 13878 1420
rect 15197 1411 15255 1417
rect 15197 1377 15209 1411
rect 15243 1408 15255 1411
rect 15930 1408 15936 1420
rect 15243 1380 15936 1408
rect 15243 1377 15255 1380
rect 15197 1371 15255 1377
rect 15930 1368 15936 1380
rect 15988 1368 15994 1420
rect 17129 1411 17187 1417
rect 17129 1377 17141 1411
rect 17175 1408 17187 1411
rect 17678 1408 17684 1420
rect 17175 1380 17684 1408
rect 17175 1377 17187 1380
rect 17129 1371 17187 1377
rect 17678 1368 17684 1380
rect 17736 1368 17742 1420
rect 20901 1411 20959 1417
rect 20901 1377 20913 1411
rect 20947 1408 20959 1411
rect 21542 1408 21548 1420
rect 20947 1380 21548 1408
rect 20947 1377 20959 1380
rect 20901 1371 20959 1377
rect 21542 1368 21548 1380
rect 21600 1368 21606 1420
rect 22833 1411 22891 1417
rect 22833 1377 22845 1411
rect 22879 1408 22891 1411
rect 23198 1408 23204 1420
rect 22879 1380 23204 1408
rect 22879 1377 22891 1380
rect 22833 1371 22891 1377
rect 23198 1368 23204 1380
rect 23256 1408 23262 1420
rect 23753 1411 23811 1417
rect 23753 1408 23765 1411
rect 23256 1380 23765 1408
rect 23256 1368 23262 1380
rect 23753 1377 23765 1380
rect 23799 1377 23811 1411
rect 24946 1408 24952 1420
rect 23753 1371 23811 1377
rect 24688 1380 24952 1408
rect 13541 1343 13599 1349
rect 13541 1309 13553 1343
rect 13587 1309 13599 1343
rect 13541 1303 13599 1309
rect 13630 1300 13636 1352
rect 13688 1340 13694 1352
rect 14277 1343 14335 1349
rect 14277 1340 14289 1343
rect 13688 1312 14289 1340
rect 13688 1300 13694 1312
rect 14277 1309 14289 1312
rect 14323 1309 14335 1343
rect 14918 1340 14924 1352
rect 14879 1312 14924 1340
rect 14277 1303 14335 1309
rect 14918 1300 14924 1312
rect 14976 1300 14982 1352
rect 15105 1343 15163 1349
rect 15105 1309 15117 1343
rect 15151 1340 15163 1343
rect 15289 1343 15347 1349
rect 15289 1340 15301 1343
rect 15151 1312 15301 1340
rect 15151 1309 15163 1312
rect 15105 1303 15163 1309
rect 15289 1309 15301 1312
rect 15335 1309 15347 1343
rect 15838 1340 15844 1352
rect 15799 1312 15844 1340
rect 15289 1303 15347 1309
rect 15838 1300 15844 1312
rect 15896 1300 15902 1352
rect 16022 1340 16028 1352
rect 15983 1312 16028 1340
rect 16022 1300 16028 1312
rect 16080 1300 16086 1352
rect 16117 1343 16175 1349
rect 16117 1309 16129 1343
rect 16163 1340 16175 1343
rect 16574 1340 16580 1352
rect 16163 1312 16580 1340
rect 16163 1309 16175 1312
rect 16117 1303 16175 1309
rect 16574 1300 16580 1312
rect 16632 1300 16638 1352
rect 16850 1340 16856 1352
rect 16811 1312 16856 1340
rect 16850 1300 16856 1312
rect 16908 1300 16914 1352
rect 17037 1343 17095 1349
rect 17037 1309 17049 1343
rect 17083 1340 17095 1343
rect 17221 1343 17279 1349
rect 17221 1340 17233 1343
rect 17083 1312 17233 1340
rect 17083 1309 17095 1312
rect 17037 1303 17095 1309
rect 17221 1309 17233 1312
rect 17267 1309 17279 1343
rect 17221 1303 17279 1309
rect 17773 1343 17831 1349
rect 17773 1309 17785 1343
rect 17819 1340 17831 1343
rect 17954 1340 17960 1352
rect 17819 1312 17960 1340
rect 17819 1309 17831 1312
rect 17773 1303 17831 1309
rect 17954 1300 17960 1312
rect 18012 1300 18018 1352
rect 18230 1300 18236 1352
rect 18288 1340 18294 1352
rect 18417 1343 18475 1349
rect 18417 1340 18429 1343
rect 18288 1312 18429 1340
rect 18288 1300 18294 1312
rect 18417 1309 18429 1312
rect 18463 1309 18475 1343
rect 18690 1340 18696 1352
rect 18651 1312 18696 1340
rect 18417 1303 18475 1309
rect 18690 1300 18696 1312
rect 18748 1300 18754 1352
rect 19334 1300 19340 1352
rect 19392 1340 19398 1352
rect 19613 1343 19671 1349
rect 19613 1340 19625 1343
rect 19392 1312 19625 1340
rect 19392 1300 19398 1312
rect 19613 1309 19625 1312
rect 19659 1309 19671 1343
rect 19613 1303 19671 1309
rect 20257 1343 20315 1349
rect 20257 1309 20269 1343
rect 20303 1340 20315 1343
rect 20714 1340 20720 1352
rect 20303 1312 20720 1340
rect 20303 1309 20315 1312
rect 20257 1303 20315 1309
rect 20714 1300 20720 1312
rect 20772 1300 20778 1352
rect 21085 1343 21143 1349
rect 21085 1309 21097 1343
rect 21131 1340 21143 1343
rect 21361 1343 21419 1349
rect 21361 1340 21373 1343
rect 21131 1312 21373 1340
rect 21131 1309 21143 1312
rect 21085 1303 21143 1309
rect 21361 1309 21373 1312
rect 21407 1309 21419 1343
rect 22002 1340 22008 1352
rect 21963 1312 22008 1340
rect 21361 1303 21419 1309
rect 22002 1300 22008 1312
rect 22060 1300 22066 1352
rect 22646 1340 22652 1352
rect 22607 1312 22652 1340
rect 22646 1300 22652 1312
rect 22704 1300 22710 1352
rect 22922 1340 22928 1352
rect 22883 1312 22928 1340
rect 22922 1300 22928 1312
rect 22980 1300 22986 1352
rect 23566 1340 23572 1352
rect 23527 1312 23572 1340
rect 23566 1300 23572 1312
rect 23624 1300 23630 1352
rect 23845 1343 23903 1349
rect 23845 1309 23857 1343
rect 23891 1340 23903 1343
rect 24688 1340 24716 1380
rect 24946 1368 24952 1380
rect 25004 1368 25010 1420
rect 25130 1408 25136 1420
rect 25091 1380 25136 1408
rect 25130 1368 25136 1380
rect 25188 1368 25194 1420
rect 26234 1408 26240 1420
rect 26195 1380 26240 1408
rect 26234 1368 26240 1380
rect 26292 1368 26298 1420
rect 31018 1408 31024 1420
rect 28920 1380 29868 1408
rect 24854 1340 24860 1352
rect 23891 1312 24716 1340
rect 24815 1312 24860 1340
rect 23891 1309 23903 1312
rect 23845 1303 23903 1309
rect 24854 1300 24860 1312
rect 24912 1300 24918 1352
rect 25041 1343 25099 1349
rect 25041 1309 25053 1343
rect 25087 1340 25099 1343
rect 25225 1343 25283 1349
rect 25225 1340 25237 1343
rect 25087 1312 25237 1340
rect 25087 1309 25099 1312
rect 25041 1303 25099 1309
rect 25225 1309 25237 1312
rect 25271 1309 25283 1343
rect 25225 1303 25283 1309
rect 25314 1300 25320 1352
rect 25372 1340 25378 1352
rect 25961 1343 26019 1349
rect 25961 1340 25973 1343
rect 25372 1312 25973 1340
rect 25372 1300 25378 1312
rect 25961 1309 25973 1312
rect 26007 1309 26019 1343
rect 25961 1303 26019 1309
rect 27430 1300 27436 1352
rect 27488 1340 27494 1352
rect 28074 1340 28080 1352
rect 27488 1312 27533 1340
rect 28035 1312 28080 1340
rect 27488 1300 27494 1312
rect 28074 1300 28080 1312
rect 28132 1300 28138 1352
rect 28261 1343 28319 1349
rect 28261 1309 28273 1343
rect 28307 1309 28319 1343
rect 28261 1303 28319 1309
rect 8352 1244 8984 1272
rect 8352 1232 8358 1244
rect 9398 1232 9404 1284
rect 9456 1272 9462 1284
rect 11885 1275 11943 1281
rect 11885 1272 11897 1275
rect 9456 1244 11897 1272
rect 9456 1232 9462 1244
rect 11885 1241 11897 1244
rect 11931 1241 11943 1275
rect 11885 1235 11943 1241
rect 11974 1232 11980 1284
rect 12032 1272 12038 1284
rect 27525 1275 27583 1281
rect 12032 1244 26464 1272
rect 12032 1232 12038 1244
rect 3234 1164 3240 1216
rect 3292 1204 3298 1216
rect 3973 1207 4031 1213
rect 3973 1204 3985 1207
rect 3292 1176 3985 1204
rect 3292 1164 3298 1176
rect 3973 1173 3985 1176
rect 4019 1173 4031 1207
rect 5626 1204 5632 1216
rect 5587 1176 5632 1204
rect 3973 1167 4031 1173
rect 5626 1164 5632 1176
rect 5684 1164 5690 1216
rect 8205 1207 8263 1213
rect 8205 1173 8217 1207
rect 8251 1204 8263 1207
rect 9674 1204 9680 1216
rect 8251 1176 9680 1204
rect 8251 1173 8263 1176
rect 8205 1167 8263 1173
rect 9674 1164 9680 1176
rect 9732 1164 9738 1216
rect 12342 1204 12348 1216
rect 12303 1176 12348 1204
rect 12342 1164 12348 1176
rect 12400 1164 12406 1216
rect 12989 1207 13047 1213
rect 12989 1173 13001 1207
rect 13035 1204 13047 1207
rect 13722 1204 13728 1216
rect 13035 1176 13728 1204
rect 13035 1173 13047 1176
rect 12989 1167 13047 1173
rect 13722 1164 13728 1176
rect 13780 1164 13786 1216
rect 14090 1204 14096 1216
rect 14051 1176 14096 1204
rect 14090 1164 14096 1176
rect 14148 1164 14154 1216
rect 14369 1207 14427 1213
rect 14369 1173 14381 1207
rect 14415 1204 14427 1207
rect 15289 1207 15347 1213
rect 15289 1204 15301 1207
rect 14415 1176 15301 1204
rect 14415 1173 14427 1176
rect 14369 1167 14427 1173
rect 15289 1173 15301 1176
rect 15335 1204 15347 1207
rect 16022 1204 16028 1216
rect 15335 1176 16028 1204
rect 15335 1173 15347 1176
rect 15289 1167 15347 1173
rect 16022 1164 16028 1176
rect 16080 1204 16086 1216
rect 17221 1207 17279 1213
rect 17221 1204 17233 1207
rect 16080 1176 17233 1204
rect 16080 1164 16086 1176
rect 17221 1173 17233 1176
rect 17267 1173 17279 1207
rect 17221 1167 17279 1173
rect 17494 1164 17500 1216
rect 17552 1204 17558 1216
rect 17589 1207 17647 1213
rect 17589 1204 17601 1207
rect 17552 1176 17601 1204
rect 17552 1164 17558 1176
rect 17589 1173 17601 1176
rect 17635 1173 17647 1207
rect 17589 1167 17647 1173
rect 19058 1164 19064 1216
rect 19116 1204 19122 1216
rect 19429 1207 19487 1213
rect 19429 1204 19441 1207
rect 19116 1176 19441 1204
rect 19116 1164 19122 1176
rect 19429 1173 19441 1176
rect 19475 1173 19487 1207
rect 19429 1167 19487 1173
rect 19702 1164 19708 1216
rect 19760 1204 19766 1216
rect 20073 1207 20131 1213
rect 20073 1204 20085 1207
rect 19760 1176 20085 1204
rect 19760 1164 19766 1176
rect 20073 1173 20085 1176
rect 20119 1173 20131 1207
rect 20073 1167 20131 1173
rect 20898 1164 20904 1216
rect 20956 1204 20962 1216
rect 21269 1207 21327 1213
rect 21269 1204 21281 1207
rect 20956 1176 21281 1204
rect 20956 1164 20962 1176
rect 21269 1173 21281 1176
rect 21315 1173 21327 1207
rect 21269 1167 21327 1173
rect 21361 1207 21419 1213
rect 21361 1173 21373 1207
rect 21407 1204 21419 1207
rect 21821 1207 21879 1213
rect 21821 1204 21833 1207
rect 21407 1176 21833 1204
rect 21407 1173 21419 1176
rect 21361 1167 21419 1173
rect 21821 1173 21833 1176
rect 21867 1173 21879 1207
rect 21821 1167 21879 1173
rect 23290 1164 23296 1216
rect 23348 1204 23354 1216
rect 23385 1207 23443 1213
rect 23385 1204 23397 1207
rect 23348 1176 23397 1204
rect 23348 1164 23354 1176
rect 23385 1173 23397 1176
rect 23431 1173 23443 1207
rect 23385 1167 23443 1173
rect 25225 1207 25283 1213
rect 25225 1173 25237 1207
rect 25271 1204 25283 1207
rect 26326 1204 26332 1216
rect 25271 1176 26332 1204
rect 25271 1173 25283 1176
rect 25225 1167 25283 1173
rect 26326 1164 26332 1176
rect 26384 1164 26390 1216
rect 26436 1204 26464 1244
rect 27525 1241 27537 1275
rect 27571 1272 27583 1275
rect 28166 1272 28172 1284
rect 27571 1244 28172 1272
rect 27571 1241 27583 1244
rect 27525 1235 27583 1241
rect 28166 1232 28172 1244
rect 28224 1232 28230 1284
rect 28276 1272 28304 1303
rect 28350 1300 28356 1352
rect 28408 1340 28414 1352
rect 28920 1340 28948 1380
rect 28408 1312 28453 1340
rect 28736 1312 28948 1340
rect 28408 1300 28414 1312
rect 28736 1272 28764 1312
rect 28994 1300 29000 1352
rect 29052 1340 29058 1352
rect 29730 1340 29736 1352
rect 29052 1312 29097 1340
rect 29691 1312 29736 1340
rect 29052 1300 29058 1312
rect 29730 1300 29736 1312
rect 29788 1300 29794 1352
rect 29840 1340 29868 1380
rect 30392 1380 31024 1408
rect 30392 1340 30420 1380
rect 31018 1368 31024 1380
rect 31076 1368 31082 1420
rect 30834 1340 30840 1352
rect 29840 1312 30420 1340
rect 30795 1312 30840 1340
rect 30834 1300 30840 1312
rect 30892 1300 30898 1352
rect 31110 1300 31116 1352
rect 31168 1340 31174 1352
rect 31168 1312 31213 1340
rect 31168 1300 31174 1312
rect 28276 1244 28764 1272
rect 28810 1232 28816 1284
rect 28868 1272 28874 1284
rect 28868 1244 32352 1272
rect 28868 1232 28874 1244
rect 29549 1207 29607 1213
rect 29549 1204 29561 1207
rect 26436 1176 29561 1204
rect 29549 1173 29561 1176
rect 29595 1173 29607 1207
rect 29549 1167 29607 1173
rect 1104 1114 32016 1136
rect 768 1040 888 1068
rect 1104 1062 7288 1114
rect 7340 1062 17592 1114
rect 17644 1062 27896 1114
rect 27948 1062 32016 1114
rect 32324 1068 32352 1244
rect 1104 1040 32016 1062
rect 32232 1040 32352 1068
rect 0 932 800 946
rect 860 932 888 1040
rect 5810 960 5816 1012
rect 5868 1000 5874 1012
rect 17221 1003 17279 1009
rect 17221 1000 17233 1003
rect 5868 972 17233 1000
rect 5868 960 5874 972
rect 17221 969 17233 972
rect 17267 969 17279 1003
rect 17221 963 17279 969
rect 17402 960 17408 1012
rect 17460 1000 17466 1012
rect 29730 1000 29736 1012
rect 17460 972 29736 1000
rect 17460 960 17466 972
rect 29730 960 29736 972
rect 29788 960 29794 1012
rect 0 904 888 932
rect 0 890 800 904
rect 8386 892 8392 944
rect 8444 932 8450 944
rect 13814 932 13820 944
rect 8444 904 13820 932
rect 8444 892 8450 904
rect 13814 892 13820 904
rect 13872 892 13878 944
rect 22002 892 22008 944
rect 22060 932 22066 944
rect 24854 932 24860 944
rect 22060 904 24860 932
rect 22060 892 22066 904
rect 24854 892 24860 904
rect 24912 892 24918 944
rect 32232 932 32260 1040
rect 32320 932 33120 946
rect 32232 904 33120 932
rect 32320 890 33120 904
rect 9214 824 9220 876
rect 9272 864 9278 876
rect 19610 864 19616 876
rect 9272 836 19616 864
rect 9272 824 9278 836
rect 19610 824 19616 836
rect 19668 824 19674 876
rect 24762 824 24768 876
rect 24820 864 24826 876
rect 28994 864 29000 876
rect 24820 836 29000 864
rect 24820 824 24826 836
rect 28994 824 29000 836
rect 29052 824 29058 876
rect 5626 756 5632 808
rect 5684 796 5690 808
rect 5684 768 22094 796
rect 5684 756 5690 768
rect 6270 688 6276 740
rect 6328 728 6334 740
rect 11974 728 11980 740
rect 6328 700 11980 728
rect 6328 688 6334 700
rect 11974 688 11980 700
rect 12032 688 12038 740
rect 22066 728 22094 768
rect 24302 756 24308 808
rect 24360 796 24366 808
rect 27430 796 27436 808
rect 24360 768 27436 796
rect 24360 756 24366 768
rect 27430 756 27436 768
rect 27488 796 27494 808
rect 31294 796 31300 808
rect 27488 768 31300 796
rect 27488 756 27494 768
rect 31294 756 31300 768
rect 31352 756 31358 808
rect 29086 728 29092 740
rect 22066 700 29092 728
rect 29086 688 29092 700
rect 29144 688 29150 740
rect 17221 663 17279 669
rect 17221 629 17233 663
rect 17267 660 17279 663
rect 28442 660 28448 672
rect 17267 632 28448 660
rect 17267 629 17279 632
rect 17221 623 17279 629
rect 28442 620 28448 632
rect 28500 620 28506 672
<< via1 >>
rect 25780 42576 25832 42628
rect 29736 42576 29788 42628
rect 25596 42508 25648 42560
rect 30104 42508 30156 42560
rect 7288 42406 7340 42458
rect 17592 42406 17644 42458
rect 27896 42406 27948 42458
rect 1216 42304 1268 42356
rect 8208 42304 8260 42356
rect 20444 42304 20496 42356
rect 1492 42168 1544 42220
rect 2872 42211 2924 42220
rect 2872 42177 2881 42211
rect 2881 42177 2915 42211
rect 2915 42177 2924 42211
rect 2872 42168 2924 42177
rect 7656 42211 7708 42220
rect 7656 42177 7665 42211
rect 7665 42177 7699 42211
rect 7699 42177 7708 42211
rect 7656 42168 7708 42177
rect 8116 42168 8168 42220
rect 9128 42211 9180 42220
rect 9128 42177 9137 42211
rect 9137 42177 9171 42211
rect 9171 42177 9180 42211
rect 9128 42168 9180 42177
rect 10232 42168 10284 42220
rect 12716 42211 12768 42220
rect 12716 42177 12725 42211
rect 12725 42177 12759 42211
rect 12759 42177 12768 42211
rect 12716 42168 12768 42177
rect 18144 42211 18196 42220
rect 3240 42100 3292 42152
rect 8392 42100 8444 42152
rect 12992 42143 13044 42152
rect 12992 42109 13001 42143
rect 13001 42109 13035 42143
rect 13035 42109 13044 42143
rect 12992 42100 13044 42109
rect 16396 42100 16448 42152
rect 18144 42177 18153 42211
rect 18153 42177 18187 42211
rect 18187 42177 18196 42211
rect 18144 42168 18196 42177
rect 19892 42168 19944 42220
rect 20444 42168 20496 42220
rect 17224 42100 17276 42152
rect 18052 42100 18104 42152
rect 19340 42100 19392 42152
rect 25412 42168 25464 42220
rect 25780 42211 25832 42220
rect 25780 42177 25789 42211
rect 25789 42177 25823 42211
rect 25823 42177 25832 42211
rect 25780 42168 25832 42177
rect 27160 42211 27212 42220
rect 27160 42177 27169 42211
rect 27169 42177 27203 42211
rect 27203 42177 27212 42211
rect 27160 42168 27212 42177
rect 28632 42211 28684 42220
rect 2596 42032 2648 42084
rect 9036 42032 9088 42084
rect 16028 42032 16080 42084
rect 18604 42032 18656 42084
rect 23020 42032 23072 42084
rect 26608 42100 26660 42152
rect 27344 42100 27396 42152
rect 28632 42177 28641 42211
rect 28641 42177 28675 42211
rect 28675 42177 28684 42211
rect 28632 42168 28684 42177
rect 29736 42211 29788 42220
rect 28816 42100 28868 42152
rect 29736 42177 29745 42211
rect 29745 42177 29779 42211
rect 29779 42177 29788 42211
rect 29736 42168 29788 42177
rect 31392 42168 31444 42220
rect 1584 41964 1636 42016
rect 2688 42007 2740 42016
rect 2688 41973 2697 42007
rect 2697 41973 2731 42007
rect 2731 41973 2740 42007
rect 2688 41964 2740 41973
rect 8576 41964 8628 42016
rect 8944 42007 8996 42016
rect 8944 41973 8953 42007
rect 8953 41973 8987 42007
rect 8987 41973 8996 42007
rect 8944 41964 8996 41973
rect 10784 41964 10836 42016
rect 12348 41964 12400 42016
rect 12900 42007 12952 42016
rect 12900 41973 12909 42007
rect 12909 41973 12943 42007
rect 12943 41973 12952 42007
rect 12900 41964 12952 41973
rect 16212 41964 16264 42016
rect 16672 42007 16724 42016
rect 16672 41973 16681 42007
rect 16681 41973 16715 42007
rect 16715 41973 16724 42007
rect 16672 41964 16724 41973
rect 19064 41964 19116 42016
rect 23572 41964 23624 42016
rect 23664 41964 23716 42016
rect 25596 42007 25648 42016
rect 25596 41973 25605 42007
rect 25605 41973 25639 42007
rect 25639 41973 25648 42007
rect 25596 41964 25648 41973
rect 26240 42007 26292 42016
rect 26240 41973 26249 42007
rect 26249 41973 26283 42007
rect 26283 41973 26292 42007
rect 26240 41964 26292 41973
rect 27252 41964 27304 42016
rect 27620 42032 27672 42084
rect 28540 42032 28592 42084
rect 28448 42007 28500 42016
rect 28448 41973 28457 42007
rect 28457 41973 28491 42007
rect 28491 41973 28500 42007
rect 28448 41964 28500 41973
rect 29368 42032 29420 42084
rect 31484 42100 31536 42152
rect 2136 41862 2188 41914
rect 12440 41862 12492 41914
rect 22744 41862 22796 41914
rect 8392 41803 8444 41812
rect 8392 41769 8401 41803
rect 8401 41769 8435 41803
rect 8435 41769 8444 41803
rect 8392 41760 8444 41769
rect 19064 41760 19116 41812
rect 27620 41760 27672 41812
rect 1400 41556 1452 41608
rect 2688 41556 2740 41608
rect 3976 41599 4028 41608
rect 3976 41565 3985 41599
rect 3985 41565 4019 41599
rect 4019 41565 4028 41599
rect 3976 41556 4028 41565
rect 8576 41692 8628 41744
rect 19432 41692 19484 41744
rect 5264 41624 5316 41676
rect 8760 41624 8812 41676
rect 4344 41556 4396 41608
rect 2688 41420 2740 41472
rect 3884 41420 3936 41472
rect 4068 41420 4120 41472
rect 4988 41556 5040 41608
rect 5356 41599 5408 41608
rect 5356 41565 5365 41599
rect 5365 41565 5399 41599
rect 5399 41565 5408 41599
rect 5356 41556 5408 41565
rect 7012 41599 7064 41608
rect 7012 41565 7021 41599
rect 7021 41565 7055 41599
rect 7055 41565 7064 41599
rect 7012 41556 7064 41565
rect 8392 41556 8444 41608
rect 11888 41556 11940 41608
rect 12348 41599 12400 41608
rect 12348 41565 12382 41599
rect 12382 41565 12400 41599
rect 12348 41556 12400 41565
rect 14004 41556 14056 41608
rect 16672 41556 16724 41608
rect 18236 41599 18288 41608
rect 18236 41565 18245 41599
rect 18245 41565 18279 41599
rect 18279 41565 18288 41599
rect 18236 41556 18288 41565
rect 18512 41599 18564 41608
rect 18512 41565 18521 41599
rect 18521 41565 18555 41599
rect 18555 41565 18564 41599
rect 18512 41556 18564 41565
rect 19524 41624 19576 41676
rect 23572 41624 23624 41676
rect 10324 41531 10376 41540
rect 10324 41497 10358 41531
rect 10358 41497 10376 41531
rect 10324 41488 10376 41497
rect 15108 41488 15160 41540
rect 19340 41488 19392 41540
rect 21640 41556 21692 41608
rect 24400 41599 24452 41608
rect 24400 41565 24409 41599
rect 24409 41565 24443 41599
rect 24443 41565 24452 41599
rect 24400 41556 24452 41565
rect 25596 41624 25648 41676
rect 31024 41624 31076 41676
rect 26424 41599 26476 41608
rect 21824 41488 21876 41540
rect 23296 41488 23348 41540
rect 24768 41488 24820 41540
rect 26424 41565 26433 41599
rect 26433 41565 26467 41599
rect 26467 41565 26476 41599
rect 26424 41556 26476 41565
rect 27620 41599 27672 41608
rect 27620 41565 27629 41599
rect 27629 41565 27663 41599
rect 27663 41565 27672 41599
rect 27620 41556 27672 41565
rect 28448 41556 28500 41608
rect 29736 41599 29788 41608
rect 29736 41565 29745 41599
rect 29745 41565 29779 41599
rect 29779 41565 29788 41599
rect 29736 41556 29788 41565
rect 29828 41556 29880 41608
rect 31300 41599 31352 41608
rect 28356 41488 28408 41540
rect 31300 41565 31309 41599
rect 31309 41565 31343 41599
rect 31343 41565 31352 41599
rect 31300 41556 31352 41565
rect 31392 41488 31444 41540
rect 5816 41463 5868 41472
rect 5816 41429 5825 41463
rect 5825 41429 5859 41463
rect 5859 41429 5868 41463
rect 5816 41420 5868 41429
rect 12256 41420 12308 41472
rect 14280 41420 14332 41472
rect 15752 41420 15804 41472
rect 17316 41463 17368 41472
rect 17316 41429 17325 41463
rect 17325 41429 17359 41463
rect 17359 41429 17368 41463
rect 17316 41420 17368 41429
rect 19156 41420 19208 41472
rect 23572 41420 23624 41472
rect 23848 41463 23900 41472
rect 23848 41429 23857 41463
rect 23857 41429 23891 41463
rect 23891 41429 23900 41463
rect 23848 41420 23900 41429
rect 26056 41420 26108 41472
rect 29644 41420 29696 41472
rect 30288 41420 30340 41472
rect 31116 41463 31168 41472
rect 31116 41429 31125 41463
rect 31125 41429 31159 41463
rect 31159 41429 31168 41463
rect 31116 41420 31168 41429
rect 7288 41318 7340 41370
rect 17592 41318 17644 41370
rect 27896 41318 27948 41370
rect 10324 41259 10376 41268
rect 10324 41225 10333 41259
rect 10333 41225 10367 41259
rect 10367 41225 10376 41259
rect 10324 41216 10376 41225
rect 11888 41216 11940 41268
rect 12716 41216 12768 41268
rect 15108 41216 15160 41268
rect 22284 41216 22336 41268
rect 1400 41123 1452 41132
rect 1400 41089 1409 41123
rect 1409 41089 1443 41123
rect 1443 41089 1452 41123
rect 1400 41080 1452 41089
rect 1676 41123 1728 41132
rect 1676 41089 1710 41123
rect 1710 41089 1728 41123
rect 4436 41148 4488 41200
rect 1676 41080 1728 41089
rect 3884 41080 3936 41132
rect 7012 41148 7064 41200
rect 8944 41148 8996 41200
rect 6920 41080 6972 41132
rect 11520 41080 11572 41132
rect 12624 41080 12676 41132
rect 13084 41080 13136 41132
rect 14096 41123 14148 41132
rect 11060 41012 11112 41064
rect 14096 41089 14105 41123
rect 14105 41089 14139 41123
rect 14139 41089 14148 41123
rect 14096 41080 14148 41089
rect 14740 41123 14792 41132
rect 14740 41089 14749 41123
rect 14749 41089 14783 41123
rect 14783 41089 14792 41123
rect 14740 41080 14792 41089
rect 14648 41012 14700 41064
rect 15752 41080 15804 41132
rect 18328 41148 18380 41200
rect 16764 41080 16816 41132
rect 18604 41148 18656 41200
rect 26056 41148 26108 41200
rect 27252 41191 27304 41200
rect 27252 41157 27286 41191
rect 27286 41157 27304 41191
rect 27252 41148 27304 41157
rect 31300 41148 31352 41200
rect 19248 41080 19300 41132
rect 20260 41080 20312 41132
rect 21272 41123 21324 41132
rect 21272 41089 21281 41123
rect 21281 41089 21315 41123
rect 21315 41089 21324 41123
rect 21272 41080 21324 41089
rect 14096 40944 14148 40996
rect 21640 41012 21692 41064
rect 22836 41012 22888 41064
rect 25780 41080 25832 41132
rect 27620 41080 27672 41132
rect 28724 41080 28776 41132
rect 28908 41080 28960 41132
rect 19800 40944 19852 40996
rect 23572 40944 23624 40996
rect 24308 41012 24360 41064
rect 25044 41055 25096 41064
rect 25044 41021 25053 41055
rect 25053 41021 25087 41055
rect 25087 41021 25096 41055
rect 25044 41012 25096 41021
rect 29920 41012 29972 41064
rect 3240 40876 3292 40928
rect 5264 40876 5316 40928
rect 8208 40876 8260 40928
rect 9680 40876 9732 40928
rect 10784 40876 10836 40928
rect 12992 40919 13044 40928
rect 12992 40885 13001 40919
rect 13001 40885 13035 40919
rect 13035 40885 13044 40919
rect 12992 40876 13044 40885
rect 13452 40876 13504 40928
rect 15660 40876 15712 40928
rect 16028 40919 16080 40928
rect 16028 40885 16037 40919
rect 16037 40885 16071 40919
rect 16071 40885 16080 40919
rect 16028 40876 16080 40885
rect 18052 40919 18104 40928
rect 18052 40885 18061 40919
rect 18061 40885 18095 40919
rect 18095 40885 18104 40919
rect 18052 40876 18104 40885
rect 19524 40876 19576 40928
rect 21088 40919 21140 40928
rect 21088 40885 21097 40919
rect 21097 40885 21131 40919
rect 21131 40885 21140 40919
rect 21088 40876 21140 40885
rect 23756 40876 23808 40928
rect 24032 40919 24084 40928
rect 24032 40885 24041 40919
rect 24041 40885 24075 40919
rect 24075 40885 24084 40919
rect 24032 40876 24084 40885
rect 26332 40876 26384 40928
rect 27344 40876 27396 40928
rect 27712 40876 27764 40928
rect 28816 40876 28868 40928
rect 29000 40876 29052 40928
rect 30472 40876 30524 40928
rect 2136 40774 2188 40826
rect 12440 40774 12492 40826
rect 22744 40774 22796 40826
rect 1492 40672 1544 40724
rect 1676 40715 1728 40724
rect 1676 40681 1685 40715
rect 1685 40681 1719 40715
rect 1719 40681 1728 40715
rect 1676 40672 1728 40681
rect 2872 40672 2924 40724
rect 7012 40715 7064 40724
rect 7012 40681 7021 40715
rect 7021 40681 7055 40715
rect 7055 40681 7064 40715
rect 7012 40672 7064 40681
rect 6920 40604 6972 40656
rect 2872 40536 2924 40588
rect 2688 40468 2740 40520
rect 3240 40511 3292 40520
rect 3240 40477 3249 40511
rect 3249 40477 3283 40511
rect 3283 40477 3292 40511
rect 3240 40468 3292 40477
rect 3516 40468 3568 40520
rect 4068 40468 4120 40520
rect 4620 40536 4672 40588
rect 4988 40536 5040 40588
rect 5356 40536 5408 40588
rect 11888 40672 11940 40724
rect 16396 40715 16448 40724
rect 16396 40681 16405 40715
rect 16405 40681 16439 40715
rect 16439 40681 16448 40715
rect 16396 40672 16448 40681
rect 22836 40672 22888 40724
rect 23296 40715 23348 40724
rect 23296 40681 23305 40715
rect 23305 40681 23339 40715
rect 23339 40681 23348 40715
rect 23296 40672 23348 40681
rect 26424 40672 26476 40724
rect 28908 40672 28960 40724
rect 4344 40468 4396 40520
rect 5172 40468 5224 40520
rect 7564 40468 7616 40520
rect 8576 40468 8628 40520
rect 8944 40468 8996 40520
rect 11428 40511 11480 40520
rect 11428 40477 11437 40511
rect 11437 40477 11471 40511
rect 11471 40477 11480 40511
rect 11428 40468 11480 40477
rect 11796 40468 11848 40520
rect 9956 40400 10008 40452
rect 10600 40332 10652 40384
rect 11060 40400 11112 40452
rect 11612 40400 11664 40452
rect 13084 40468 13136 40520
rect 13452 40511 13504 40520
rect 13452 40477 13461 40511
rect 13461 40477 13495 40511
rect 13495 40477 13504 40511
rect 13452 40468 13504 40477
rect 14004 40468 14056 40520
rect 14648 40400 14700 40452
rect 15292 40400 15344 40452
rect 10876 40332 10928 40384
rect 12808 40375 12860 40384
rect 12808 40341 12817 40375
rect 12817 40341 12851 40375
rect 12851 40341 12860 40375
rect 12808 40332 12860 40341
rect 15476 40332 15528 40384
rect 17224 40604 17276 40656
rect 25596 40604 25648 40656
rect 26056 40604 26108 40656
rect 16580 40511 16632 40520
rect 16580 40477 16589 40511
rect 16589 40477 16623 40511
rect 16623 40477 16632 40511
rect 16580 40468 16632 40477
rect 17316 40468 17368 40520
rect 18236 40536 18288 40588
rect 19248 40579 19300 40588
rect 19248 40545 19257 40579
rect 19257 40545 19291 40579
rect 19291 40545 19300 40579
rect 19248 40536 19300 40545
rect 17132 40400 17184 40452
rect 18052 40468 18104 40520
rect 19156 40468 19208 40520
rect 20720 40468 20772 40520
rect 22284 40468 22336 40520
rect 23020 40536 23072 40588
rect 23480 40511 23532 40520
rect 18512 40400 18564 40452
rect 22192 40400 22244 40452
rect 23480 40477 23489 40511
rect 23489 40477 23523 40511
rect 23523 40477 23532 40511
rect 23480 40468 23532 40477
rect 23572 40468 23624 40520
rect 24032 40536 24084 40588
rect 23756 40511 23808 40520
rect 23756 40477 23765 40511
rect 23765 40477 23799 40511
rect 23799 40477 23808 40511
rect 24400 40511 24452 40520
rect 23756 40468 23808 40477
rect 24400 40477 24409 40511
rect 24409 40477 24443 40511
rect 24443 40477 24452 40511
rect 24400 40468 24452 40477
rect 25044 40468 25096 40520
rect 25780 40468 25832 40520
rect 26240 40468 26292 40520
rect 26700 40511 26752 40520
rect 26700 40477 26709 40511
rect 26709 40477 26743 40511
rect 26743 40477 26752 40511
rect 26700 40468 26752 40477
rect 26976 40604 27028 40656
rect 29920 40672 29972 40724
rect 30288 40672 30340 40724
rect 27344 40536 27396 40588
rect 26976 40468 27028 40520
rect 27804 40511 27856 40520
rect 27804 40477 27813 40511
rect 27813 40477 27847 40511
rect 27847 40477 27856 40511
rect 27804 40468 27856 40477
rect 28724 40536 28776 40588
rect 29552 40579 29604 40588
rect 29552 40545 29561 40579
rect 29561 40545 29595 40579
rect 29595 40545 29604 40579
rect 29552 40536 29604 40545
rect 28264 40468 28316 40520
rect 28448 40468 28500 40520
rect 24492 40400 24544 40452
rect 28080 40400 28132 40452
rect 28816 40511 28868 40520
rect 28816 40477 28825 40511
rect 28825 40477 28859 40511
rect 28859 40477 28868 40511
rect 28816 40468 28868 40477
rect 28908 40511 28960 40520
rect 28908 40477 28917 40511
rect 28917 40477 28951 40511
rect 28951 40477 28960 40511
rect 28908 40468 28960 40477
rect 29644 40468 29696 40520
rect 16948 40332 17000 40384
rect 19432 40332 19484 40384
rect 22008 40332 22060 40384
rect 25872 40332 25924 40384
rect 28448 40332 28500 40384
rect 30932 40375 30984 40384
rect 30932 40341 30941 40375
rect 30941 40341 30975 40375
rect 30975 40341 30984 40375
rect 30932 40332 30984 40341
rect 7288 40230 7340 40282
rect 17592 40230 17644 40282
rect 27896 40230 27948 40282
rect 3976 40128 4028 40180
rect 5356 40128 5408 40180
rect 7564 40171 7616 40180
rect 2596 39992 2648 40044
rect 3516 40035 3568 40044
rect 3516 40001 3525 40035
rect 3525 40001 3559 40035
rect 3559 40001 3568 40035
rect 3516 39992 3568 40001
rect 5264 40060 5316 40112
rect 7564 40137 7573 40171
rect 7573 40137 7607 40171
rect 7607 40137 7616 40171
rect 7564 40128 7616 40137
rect 9128 40128 9180 40180
rect 9956 40171 10008 40180
rect 9956 40137 9965 40171
rect 9965 40137 9999 40171
rect 9999 40137 10008 40171
rect 9956 40128 10008 40137
rect 11520 40171 11572 40180
rect 11520 40137 11529 40171
rect 11529 40137 11563 40171
rect 11563 40137 11572 40171
rect 11520 40128 11572 40137
rect 4436 40035 4488 40044
rect 1400 39967 1452 39976
rect 1400 39933 1409 39967
rect 1409 39933 1443 39967
rect 1443 39933 1452 39967
rect 1400 39924 1452 39933
rect 4436 40001 4445 40035
rect 4445 40001 4479 40035
rect 4479 40001 4488 40035
rect 4436 39992 4488 40001
rect 4528 39992 4580 40044
rect 5816 39992 5868 40044
rect 6736 40035 6788 40044
rect 6736 40001 6745 40035
rect 6745 40001 6779 40035
rect 6779 40001 6788 40035
rect 6736 39992 6788 40001
rect 7104 39992 7156 40044
rect 7932 40060 7984 40112
rect 10232 40060 10284 40112
rect 10416 40060 10468 40112
rect 8208 40035 8260 40044
rect 8208 40001 8217 40035
rect 8217 40001 8251 40035
rect 8251 40001 8260 40035
rect 8208 39992 8260 40001
rect 9036 40035 9088 40044
rect 9036 40001 9045 40035
rect 9045 40001 9079 40035
rect 9079 40001 9088 40035
rect 9036 39992 9088 40001
rect 8300 39924 8352 39976
rect 9680 39992 9732 40044
rect 10876 39992 10928 40044
rect 11428 39992 11480 40044
rect 8208 39856 8260 39908
rect 11796 39992 11848 40044
rect 12256 39992 12308 40044
rect 12624 40035 12676 40044
rect 12624 40001 12633 40035
rect 12633 40001 12667 40035
rect 12667 40001 12676 40035
rect 12624 39992 12676 40001
rect 12808 40035 12860 40044
rect 12808 40001 12817 40035
rect 12817 40001 12851 40035
rect 12851 40001 12860 40035
rect 12808 39992 12860 40001
rect 15384 40060 15436 40112
rect 14648 40035 14700 40044
rect 12348 39924 12400 39976
rect 13820 39924 13872 39976
rect 12532 39856 12584 39908
rect 14648 40001 14657 40035
rect 14657 40001 14691 40035
rect 14691 40001 14700 40035
rect 14648 39992 14700 40001
rect 15292 40035 15344 40044
rect 15292 40001 15301 40035
rect 15301 40001 15335 40035
rect 15335 40001 15344 40035
rect 15292 39992 15344 40001
rect 17224 40060 17276 40112
rect 18236 40128 18288 40180
rect 23480 40128 23532 40180
rect 16580 39992 16632 40044
rect 17132 40035 17184 40044
rect 17132 40001 17141 40035
rect 17141 40001 17175 40035
rect 17175 40001 17184 40035
rect 17132 39992 17184 40001
rect 18512 39992 18564 40044
rect 22192 40060 22244 40112
rect 24584 40060 24636 40112
rect 26240 40128 26292 40180
rect 26884 40128 26936 40180
rect 27160 40128 27212 40180
rect 28080 40171 28132 40180
rect 28080 40137 28089 40171
rect 28089 40137 28123 40171
rect 28123 40137 28132 40171
rect 28080 40128 28132 40137
rect 28632 40128 28684 40180
rect 21824 40035 21876 40044
rect 21824 40001 21833 40035
rect 21833 40001 21867 40035
rect 21867 40001 21876 40035
rect 21824 39992 21876 40001
rect 22836 39992 22888 40044
rect 23020 40035 23072 40044
rect 23020 40001 23029 40035
rect 23029 40001 23063 40035
rect 23063 40001 23072 40035
rect 23020 39992 23072 40001
rect 23296 40035 23348 40044
rect 23296 40001 23305 40035
rect 23305 40001 23339 40035
rect 23339 40001 23348 40035
rect 23296 39992 23348 40001
rect 23848 39992 23900 40044
rect 26700 40060 26752 40112
rect 25964 39992 26016 40044
rect 27804 40060 27856 40112
rect 15200 39924 15252 39976
rect 16212 39924 16264 39976
rect 18420 39967 18472 39976
rect 14740 39856 14792 39908
rect 18420 39933 18429 39967
rect 18429 39933 18463 39967
rect 18463 39933 18472 39967
rect 18420 39924 18472 39933
rect 19708 39924 19760 39976
rect 22192 39924 22244 39976
rect 22928 39924 22980 39976
rect 23664 39924 23716 39976
rect 27712 39992 27764 40044
rect 30656 40060 30708 40112
rect 28724 40035 28776 40044
rect 28724 40001 28733 40035
rect 28733 40001 28767 40035
rect 28767 40001 28776 40035
rect 28724 39992 28776 40001
rect 28908 39992 28960 40044
rect 29644 40035 29696 40044
rect 29644 40001 29653 40035
rect 29653 40001 29687 40035
rect 29687 40001 29696 40035
rect 29644 39992 29696 40001
rect 29828 40035 29880 40044
rect 29828 40001 29837 40035
rect 29837 40001 29871 40035
rect 29871 40001 29880 40035
rect 29828 39992 29880 40001
rect 30472 40035 30524 40044
rect 30472 40001 30481 40035
rect 30481 40001 30515 40035
rect 30515 40001 30524 40035
rect 30472 39992 30524 40001
rect 24860 39856 24912 39908
rect 29460 39924 29512 39976
rect 28264 39856 28316 39908
rect 28816 39856 28868 39908
rect 29644 39856 29696 39908
rect 31300 39992 31352 40044
rect 2872 39788 2924 39840
rect 3792 39788 3844 39840
rect 5908 39788 5960 39840
rect 7196 39788 7248 39840
rect 9036 39788 9088 39840
rect 10784 39788 10836 39840
rect 12624 39788 12676 39840
rect 12900 39788 12952 39840
rect 15660 39831 15712 39840
rect 15660 39797 15669 39831
rect 15669 39797 15703 39831
rect 15703 39797 15712 39831
rect 15660 39788 15712 39797
rect 22468 39788 22520 39840
rect 23572 39788 23624 39840
rect 2136 39686 2188 39738
rect 12440 39686 12492 39738
rect 22744 39686 22796 39738
rect 2596 39627 2648 39636
rect 2596 39593 2605 39627
rect 2605 39593 2639 39627
rect 2639 39593 2648 39627
rect 2596 39584 2648 39593
rect 7196 39584 7248 39636
rect 8392 39584 8444 39636
rect 12624 39584 12676 39636
rect 16764 39627 16816 39636
rect 16764 39593 16773 39627
rect 16773 39593 16807 39627
rect 16807 39593 16816 39627
rect 16764 39584 16816 39593
rect 18144 39584 18196 39636
rect 22836 39627 22888 39636
rect 22836 39593 22845 39627
rect 22845 39593 22879 39627
rect 22879 39593 22888 39627
rect 22836 39584 22888 39593
rect 24492 39584 24544 39636
rect 12072 39516 12124 39568
rect 15660 39516 15712 39568
rect 23572 39516 23624 39568
rect 25964 39516 26016 39568
rect 2688 39448 2740 39500
rect 3240 39448 3292 39500
rect 4620 39491 4672 39500
rect 2780 39423 2832 39432
rect 2780 39389 2789 39423
rect 2789 39389 2823 39423
rect 2823 39389 2832 39423
rect 3056 39423 3108 39432
rect 2780 39380 2832 39389
rect 3056 39389 3065 39423
rect 3065 39389 3099 39423
rect 3099 39389 3108 39423
rect 3056 39380 3108 39389
rect 4252 39423 4304 39432
rect 4252 39389 4261 39423
rect 4261 39389 4295 39423
rect 4295 39389 4304 39423
rect 4252 39380 4304 39389
rect 4620 39457 4629 39491
rect 4629 39457 4663 39491
rect 4663 39457 4672 39491
rect 4620 39448 4672 39457
rect 3792 39312 3844 39364
rect 7104 39423 7156 39432
rect 6644 39312 6696 39364
rect 1860 39287 1912 39296
rect 1860 39253 1869 39287
rect 1869 39253 1903 39287
rect 1903 39253 1912 39287
rect 1860 39244 1912 39253
rect 5448 39244 5500 39296
rect 7104 39389 7113 39423
rect 7113 39389 7147 39423
rect 7147 39389 7156 39423
rect 7104 39380 7156 39389
rect 7932 39423 7984 39432
rect 7932 39389 7941 39423
rect 7941 39389 7975 39423
rect 7975 39389 7984 39423
rect 7932 39380 7984 39389
rect 8300 39380 8352 39432
rect 6828 39312 6880 39364
rect 8484 39380 8536 39432
rect 9036 39380 9088 39432
rect 10324 39380 10376 39432
rect 10784 39423 10836 39432
rect 10784 39389 10793 39423
rect 10793 39389 10827 39423
rect 10827 39389 10836 39423
rect 10784 39380 10836 39389
rect 12256 39312 12308 39364
rect 9680 39244 9732 39296
rect 9772 39244 9824 39296
rect 11980 39244 12032 39296
rect 13084 39380 13136 39432
rect 14648 39448 14700 39500
rect 17316 39448 17368 39500
rect 17500 39448 17552 39500
rect 13820 39380 13872 39432
rect 15384 39380 15436 39432
rect 15844 39423 15896 39432
rect 15844 39389 15853 39423
rect 15853 39389 15887 39423
rect 15887 39389 15896 39423
rect 16948 39423 17000 39432
rect 15844 39380 15896 39389
rect 16948 39389 16957 39423
rect 16957 39389 16991 39423
rect 16991 39389 17000 39423
rect 16948 39380 17000 39389
rect 18420 39448 18472 39500
rect 20996 39448 21048 39500
rect 23848 39448 23900 39500
rect 24676 39448 24728 39500
rect 27804 39448 27856 39500
rect 29552 39448 29604 39500
rect 18236 39423 18288 39432
rect 18236 39389 18245 39423
rect 18245 39389 18279 39423
rect 18279 39389 18288 39423
rect 18236 39380 18288 39389
rect 18512 39423 18564 39432
rect 18512 39389 18521 39423
rect 18521 39389 18555 39423
rect 18555 39389 18564 39423
rect 18512 39380 18564 39389
rect 19432 39423 19484 39432
rect 17408 39312 17460 39364
rect 19432 39389 19441 39423
rect 19441 39389 19475 39423
rect 19475 39389 19484 39423
rect 19432 39380 19484 39389
rect 21180 39380 21232 39432
rect 23020 39423 23072 39432
rect 23020 39389 23029 39423
rect 23029 39389 23063 39423
rect 23063 39389 23072 39423
rect 23020 39380 23072 39389
rect 23296 39423 23348 39432
rect 23296 39389 23305 39423
rect 23305 39389 23339 39423
rect 23339 39389 23348 39423
rect 23296 39380 23348 39389
rect 24308 39380 24360 39432
rect 24584 39423 24636 39432
rect 24584 39389 24593 39423
rect 24593 39389 24627 39423
rect 24627 39389 24636 39423
rect 24584 39380 24636 39389
rect 25872 39423 25924 39432
rect 25872 39389 25881 39423
rect 25881 39389 25915 39423
rect 25915 39389 25924 39423
rect 25872 39380 25924 39389
rect 26240 39423 26292 39432
rect 26240 39389 26249 39423
rect 26249 39389 26283 39423
rect 26283 39389 26292 39423
rect 26240 39380 26292 39389
rect 28632 39423 28684 39432
rect 19524 39312 19576 39364
rect 20628 39355 20680 39364
rect 20628 39321 20637 39355
rect 20637 39321 20671 39355
rect 20671 39321 20680 39355
rect 20628 39312 20680 39321
rect 25596 39312 25648 39364
rect 26332 39312 26384 39364
rect 28632 39389 28641 39423
rect 28641 39389 28675 39423
rect 28675 39389 28684 39423
rect 28632 39380 28684 39389
rect 29184 39312 29236 39364
rect 30472 39312 30524 39364
rect 13360 39244 13412 39296
rect 15384 39287 15436 39296
rect 15384 39253 15393 39287
rect 15393 39253 15427 39287
rect 15427 39253 15436 39287
rect 15384 39244 15436 39253
rect 20076 39244 20128 39296
rect 21640 39244 21692 39296
rect 27160 39244 27212 39296
rect 31300 39287 31352 39296
rect 31300 39253 31309 39287
rect 31309 39253 31343 39287
rect 31343 39253 31352 39287
rect 31300 39244 31352 39253
rect 7288 39142 7340 39194
rect 17592 39142 17644 39194
rect 27896 39142 27948 39194
rect 2780 39040 2832 39092
rect 2412 38947 2464 38956
rect 2412 38913 2421 38947
rect 2421 38913 2455 38947
rect 2455 38913 2464 38947
rect 2412 38904 2464 38913
rect 3516 39040 3568 39092
rect 4620 38972 4672 39024
rect 3792 38947 3844 38956
rect 3792 38913 3801 38947
rect 3801 38913 3835 38947
rect 3835 38913 3844 38947
rect 3792 38904 3844 38913
rect 5908 38972 5960 39024
rect 2780 38836 2832 38888
rect 5172 38947 5224 38956
rect 5172 38913 5182 38947
rect 5182 38913 5216 38947
rect 5216 38913 5224 38947
rect 5356 38947 5408 38956
rect 5172 38904 5224 38913
rect 5356 38913 5365 38947
rect 5365 38913 5399 38947
rect 5399 38913 5408 38947
rect 5356 38904 5408 38913
rect 2228 38743 2280 38752
rect 2228 38709 2237 38743
rect 2237 38709 2271 38743
rect 2271 38709 2280 38743
rect 2228 38700 2280 38709
rect 2688 38700 2740 38752
rect 5264 38836 5316 38888
rect 5632 38904 5684 38956
rect 6552 38947 6604 38956
rect 6552 38913 6561 38947
rect 6561 38913 6595 38947
rect 6595 38913 6604 38947
rect 6552 38904 6604 38913
rect 8116 39040 8168 39092
rect 8208 39040 8260 39092
rect 10324 39083 10376 39092
rect 7656 38947 7708 38956
rect 7656 38913 7665 38947
rect 7665 38913 7699 38947
rect 7699 38913 7708 38947
rect 7656 38904 7708 38913
rect 7932 38904 7984 38956
rect 8760 38947 8812 38956
rect 8392 38836 8444 38888
rect 8760 38913 8769 38947
rect 8769 38913 8803 38947
rect 8803 38913 8812 38947
rect 8760 38904 8812 38913
rect 10324 39049 10333 39083
rect 10333 39049 10367 39083
rect 10367 39049 10376 39083
rect 10324 39040 10376 39049
rect 10784 39040 10836 39092
rect 19432 39040 19484 39092
rect 12532 38972 12584 39024
rect 15384 38972 15436 39024
rect 10968 38947 11020 38956
rect 10968 38913 10977 38947
rect 10977 38913 11011 38947
rect 11011 38913 11020 38947
rect 10968 38904 11020 38913
rect 11888 38947 11940 38956
rect 11888 38913 11897 38947
rect 11897 38913 11931 38947
rect 11931 38913 11940 38947
rect 11888 38904 11940 38913
rect 11980 38904 12032 38956
rect 15292 38904 15344 38956
rect 18052 38972 18104 39024
rect 15936 38947 15988 38956
rect 15936 38913 15945 38947
rect 15945 38913 15979 38947
rect 15979 38913 15988 38947
rect 15936 38904 15988 38913
rect 17224 38947 17276 38956
rect 17224 38913 17233 38947
rect 17233 38913 17267 38947
rect 17267 38913 17276 38947
rect 17224 38904 17276 38913
rect 17408 38904 17460 38956
rect 7932 38768 7984 38820
rect 8208 38768 8260 38820
rect 8944 38768 8996 38820
rect 5724 38743 5776 38752
rect 5724 38709 5733 38743
rect 5733 38709 5767 38743
rect 5767 38709 5776 38743
rect 5724 38700 5776 38709
rect 7748 38700 7800 38752
rect 8300 38700 8352 38752
rect 11796 38836 11848 38888
rect 14004 38879 14056 38888
rect 14004 38845 14013 38879
rect 14013 38845 14047 38879
rect 14047 38845 14056 38879
rect 14004 38836 14056 38845
rect 15568 38836 15620 38888
rect 15200 38768 15252 38820
rect 17408 38768 17460 38820
rect 18328 38904 18380 38956
rect 18880 38904 18932 38956
rect 21548 38972 21600 39024
rect 23296 39040 23348 39092
rect 20444 38947 20496 38956
rect 20444 38913 20453 38947
rect 20453 38913 20487 38947
rect 20487 38913 20496 38947
rect 20444 38904 20496 38913
rect 22284 38947 22336 38956
rect 22284 38913 22293 38947
rect 22293 38913 22327 38947
rect 22327 38913 22336 38947
rect 22284 38904 22336 38913
rect 22928 38972 22980 39024
rect 23020 38904 23072 38956
rect 23388 38947 23440 38956
rect 23388 38913 23397 38947
rect 23397 38913 23431 38947
rect 23431 38913 23440 38947
rect 23388 38904 23440 38913
rect 28724 39040 28776 39092
rect 30472 39083 30524 39092
rect 30472 39049 30481 39083
rect 30481 39049 30515 39083
rect 30515 39049 30524 39083
rect 30472 39040 30524 39049
rect 25596 38972 25648 39024
rect 31300 38972 31352 39024
rect 24584 38904 24636 38956
rect 27620 38947 27672 38956
rect 20628 38836 20680 38888
rect 27620 38913 27629 38947
rect 27629 38913 27663 38947
rect 27663 38913 27672 38947
rect 27620 38904 27672 38913
rect 28448 38947 28500 38956
rect 28448 38913 28457 38947
rect 28457 38913 28491 38947
rect 28491 38913 28500 38947
rect 28448 38904 28500 38913
rect 28816 38904 28868 38956
rect 30656 38947 30708 38956
rect 30656 38913 30665 38947
rect 30665 38913 30699 38947
rect 30699 38913 30708 38947
rect 30656 38904 30708 38913
rect 31024 38904 31076 38956
rect 25872 38836 25924 38888
rect 29184 38879 29236 38888
rect 29184 38845 29193 38879
rect 29193 38845 29227 38879
rect 29227 38845 29236 38879
rect 29184 38836 29236 38845
rect 29644 38836 29696 38888
rect 30012 38836 30064 38888
rect 30932 38879 30984 38888
rect 30932 38845 30941 38879
rect 30941 38845 30975 38879
rect 30975 38845 30984 38879
rect 30932 38836 30984 38845
rect 20904 38768 20956 38820
rect 21916 38768 21968 38820
rect 23664 38768 23716 38820
rect 24768 38768 24820 38820
rect 28356 38768 28408 38820
rect 11520 38700 11572 38752
rect 12164 38700 12216 38752
rect 13820 38700 13872 38752
rect 14648 38700 14700 38752
rect 16580 38700 16632 38752
rect 18512 38700 18564 38752
rect 22284 38700 22336 38752
rect 24216 38700 24268 38752
rect 25780 38700 25832 38752
rect 27804 38743 27856 38752
rect 27804 38709 27813 38743
rect 27813 38709 27847 38743
rect 27847 38709 27856 38743
rect 27804 38700 27856 38709
rect 2136 38598 2188 38650
rect 12440 38598 12492 38650
rect 22744 38598 22796 38650
rect 3056 38496 3108 38548
rect 5448 38539 5500 38548
rect 5448 38505 5457 38539
rect 5457 38505 5491 38539
rect 5491 38505 5500 38539
rect 5448 38496 5500 38505
rect 6552 38496 6604 38548
rect 11888 38539 11940 38548
rect 11888 38505 11897 38539
rect 11897 38505 11931 38539
rect 11931 38505 11940 38539
rect 11888 38496 11940 38505
rect 12072 38496 12124 38548
rect 14280 38496 14332 38548
rect 4436 38428 4488 38480
rect 4528 38428 4580 38480
rect 5356 38428 5408 38480
rect 7656 38471 7708 38480
rect 7656 38437 7665 38471
rect 7665 38437 7699 38471
rect 7699 38437 7708 38471
rect 7656 38428 7708 38437
rect 8760 38428 8812 38480
rect 1400 38292 1452 38344
rect 2872 38292 2924 38344
rect 5448 38360 5500 38412
rect 8024 38360 8076 38412
rect 4436 38335 4488 38344
rect 4436 38301 4445 38335
rect 4445 38301 4479 38335
rect 4479 38301 4488 38335
rect 4436 38292 4488 38301
rect 2228 38224 2280 38276
rect 4528 38224 4580 38276
rect 5540 38335 5592 38344
rect 5540 38301 5549 38335
rect 5549 38301 5583 38335
rect 5583 38301 5592 38335
rect 5540 38292 5592 38301
rect 8300 38292 8352 38344
rect 11704 38428 11756 38480
rect 14004 38428 14056 38480
rect 17224 38496 17276 38548
rect 19064 38496 19116 38548
rect 22928 38496 22980 38548
rect 19340 38428 19392 38480
rect 9312 38335 9364 38344
rect 9312 38301 9321 38335
rect 9321 38301 9355 38335
rect 9355 38301 9364 38335
rect 9312 38292 9364 38301
rect 8208 38267 8260 38276
rect 8208 38233 8217 38267
rect 8217 38233 8251 38267
rect 8251 38233 8260 38267
rect 8208 38224 8260 38233
rect 8392 38224 8444 38276
rect 12072 38292 12124 38344
rect 12532 38292 12584 38344
rect 13084 38292 13136 38344
rect 13360 38292 13412 38344
rect 14188 38335 14240 38344
rect 14188 38301 14197 38335
rect 14197 38301 14231 38335
rect 14231 38301 14240 38335
rect 14188 38292 14240 38301
rect 10232 38224 10284 38276
rect 10600 38267 10652 38276
rect 10600 38233 10609 38267
rect 10609 38233 10643 38267
rect 10643 38233 10652 38267
rect 10600 38224 10652 38233
rect 17040 38360 17092 38412
rect 18512 38360 18564 38412
rect 23756 38360 23808 38412
rect 17500 38335 17552 38344
rect 17500 38301 17509 38335
rect 17509 38301 17543 38335
rect 17543 38301 17552 38335
rect 17500 38292 17552 38301
rect 17684 38292 17736 38344
rect 17776 38292 17828 38344
rect 19616 38292 19668 38344
rect 21640 38335 21692 38344
rect 21640 38301 21649 38335
rect 21649 38301 21683 38335
rect 21683 38301 21692 38335
rect 21640 38292 21692 38301
rect 23664 38335 23716 38344
rect 23664 38301 23673 38335
rect 23673 38301 23707 38335
rect 23707 38301 23716 38335
rect 23664 38292 23716 38301
rect 24400 38335 24452 38344
rect 24400 38301 24409 38335
rect 24409 38301 24443 38335
rect 24443 38301 24452 38335
rect 24400 38292 24452 38301
rect 24676 38360 24728 38412
rect 24860 38335 24912 38344
rect 24860 38301 24874 38335
rect 24874 38301 24908 38335
rect 24908 38301 24912 38335
rect 24860 38292 24912 38301
rect 20076 38267 20128 38276
rect 8116 38156 8168 38208
rect 9956 38199 10008 38208
rect 9956 38165 9965 38199
rect 9965 38165 9999 38199
rect 9999 38165 10008 38199
rect 9956 38156 10008 38165
rect 11796 38156 11848 38208
rect 13820 38156 13872 38208
rect 18236 38199 18288 38208
rect 18236 38165 18245 38199
rect 18245 38165 18279 38199
rect 18279 38165 18288 38199
rect 18236 38156 18288 38165
rect 20076 38233 20110 38267
rect 20110 38233 20128 38267
rect 20076 38224 20128 38233
rect 20996 38224 21048 38276
rect 20904 38156 20956 38208
rect 22100 38224 22152 38276
rect 26240 38428 26292 38480
rect 26148 38335 26200 38344
rect 26148 38301 26157 38335
rect 26157 38301 26191 38335
rect 26191 38301 26200 38335
rect 26148 38292 26200 38301
rect 27620 38496 27672 38548
rect 27804 38496 27856 38548
rect 29736 38496 29788 38548
rect 31024 38539 31076 38548
rect 31024 38505 31033 38539
rect 31033 38505 31067 38539
rect 31067 38505 31076 38539
rect 31024 38496 31076 38505
rect 27712 38428 27764 38480
rect 27068 38335 27120 38344
rect 27068 38301 27077 38335
rect 27077 38301 27111 38335
rect 27111 38301 27120 38335
rect 27068 38292 27120 38301
rect 27160 38335 27212 38344
rect 27160 38301 27169 38335
rect 27169 38301 27203 38335
rect 27203 38301 27212 38335
rect 27160 38292 27212 38301
rect 25320 38224 25372 38276
rect 25872 38267 25924 38276
rect 25872 38233 25881 38267
rect 25881 38233 25915 38267
rect 25915 38233 25924 38267
rect 25872 38224 25924 38233
rect 27804 38335 27856 38344
rect 27804 38301 27813 38335
rect 27813 38301 27847 38335
rect 27847 38301 27856 38335
rect 27804 38292 27856 38301
rect 27988 38335 28040 38344
rect 27988 38301 27997 38335
rect 27997 38301 28031 38335
rect 28031 38301 28040 38335
rect 27988 38292 28040 38301
rect 28724 38335 28776 38344
rect 28724 38301 28733 38335
rect 28733 38301 28767 38335
rect 28767 38301 28776 38335
rect 28724 38292 28776 38301
rect 29460 38292 29512 38344
rect 29736 38335 29788 38344
rect 29736 38301 29745 38335
rect 29745 38301 29779 38335
rect 29779 38301 29788 38335
rect 29736 38292 29788 38301
rect 30012 38335 30064 38344
rect 30012 38301 30021 38335
rect 30021 38301 30055 38335
rect 30055 38301 30064 38335
rect 30012 38292 30064 38301
rect 30932 38360 30984 38412
rect 31300 38360 31352 38412
rect 24492 38156 24544 38208
rect 25688 38156 25740 38208
rect 26332 38156 26384 38208
rect 27436 38156 27488 38208
rect 29828 38224 29880 38276
rect 30288 38292 30340 38344
rect 30656 38199 30708 38208
rect 30656 38165 30665 38199
rect 30665 38165 30699 38199
rect 30699 38165 30708 38199
rect 30656 38156 30708 38165
rect 7288 38054 7340 38106
rect 17592 38054 17644 38106
rect 27896 38054 27948 38106
rect 2412 37952 2464 38004
rect 5540 37952 5592 38004
rect 8760 37952 8812 38004
rect 10968 37952 11020 38004
rect 11888 37952 11940 38004
rect 3056 37884 3108 37936
rect 1308 37816 1360 37868
rect 4436 37884 4488 37936
rect 5632 37884 5684 37936
rect 9312 37884 9364 37936
rect 2320 37612 2372 37664
rect 4252 37816 4304 37868
rect 5540 37859 5592 37868
rect 5540 37825 5549 37859
rect 5549 37825 5583 37859
rect 5583 37825 5592 37859
rect 5540 37816 5592 37825
rect 5816 37816 5868 37868
rect 6552 37859 6604 37868
rect 6552 37825 6561 37859
rect 6561 37825 6595 37859
rect 6595 37825 6604 37859
rect 6552 37816 6604 37825
rect 7564 37816 7616 37868
rect 9772 37859 9824 37868
rect 9772 37825 9806 37859
rect 9806 37825 9824 37859
rect 9772 37816 9824 37825
rect 11796 37816 11848 37868
rect 4160 37748 4212 37800
rect 5448 37748 5500 37800
rect 5540 37680 5592 37732
rect 6092 37680 6144 37732
rect 14188 37952 14240 38004
rect 18880 37995 18932 38004
rect 12072 37884 12124 37936
rect 15844 37884 15896 37936
rect 18236 37884 18288 37936
rect 18880 37961 18889 37995
rect 18889 37961 18923 37995
rect 18923 37961 18932 37995
rect 18880 37952 18932 37961
rect 21180 37995 21232 38004
rect 21180 37961 21189 37995
rect 21189 37961 21223 37995
rect 21223 37961 21232 37995
rect 21180 37952 21232 37961
rect 22100 37995 22152 38004
rect 22100 37961 22109 37995
rect 22109 37961 22143 37995
rect 22143 37961 22152 37995
rect 22100 37952 22152 37961
rect 24400 37952 24452 38004
rect 26148 37952 26200 38004
rect 26516 37952 26568 38004
rect 13636 37816 13688 37868
rect 14280 37859 14332 37868
rect 14280 37825 14289 37859
rect 14289 37825 14323 37859
rect 14323 37825 14332 37859
rect 14280 37816 14332 37825
rect 12072 37748 12124 37800
rect 3792 37612 3844 37664
rect 11980 37612 12032 37664
rect 12624 37680 12676 37732
rect 12716 37680 12768 37732
rect 13728 37748 13780 37800
rect 14188 37748 14240 37800
rect 14464 37680 14516 37732
rect 15200 37859 15252 37868
rect 15200 37825 15210 37859
rect 15210 37825 15244 37859
rect 15244 37825 15252 37859
rect 15200 37816 15252 37825
rect 15384 37859 15436 37868
rect 15384 37825 15393 37859
rect 15393 37825 15427 37859
rect 15427 37825 15436 37859
rect 15384 37816 15436 37825
rect 15568 37859 15620 37868
rect 15568 37825 15582 37859
rect 15582 37825 15616 37859
rect 15616 37825 15620 37859
rect 19064 37859 19116 37868
rect 15568 37816 15620 37825
rect 19064 37825 19073 37859
rect 19073 37825 19107 37859
rect 19107 37825 19116 37859
rect 19064 37816 19116 37825
rect 19340 37859 19392 37868
rect 19340 37825 19349 37859
rect 19349 37825 19383 37859
rect 19383 37825 19392 37859
rect 19340 37816 19392 37825
rect 19616 37816 19668 37868
rect 20536 37816 20588 37868
rect 15200 37680 15252 37732
rect 16856 37748 16908 37800
rect 19156 37748 19208 37800
rect 22928 37884 22980 37936
rect 24768 37884 24820 37936
rect 22284 37859 22336 37868
rect 22284 37825 22293 37859
rect 22293 37825 22327 37859
rect 22327 37825 22336 37859
rect 22284 37816 22336 37825
rect 22468 37859 22520 37868
rect 22468 37825 22477 37859
rect 22477 37825 22511 37859
rect 22511 37825 22520 37859
rect 22468 37816 22520 37825
rect 24216 37859 24268 37868
rect 24216 37825 24225 37859
rect 24225 37825 24259 37859
rect 24259 37825 24268 37859
rect 24216 37816 24268 37825
rect 24308 37859 24360 37868
rect 24308 37825 24317 37859
rect 24317 37825 24351 37859
rect 24351 37825 24360 37859
rect 24492 37859 24544 37868
rect 24308 37816 24360 37825
rect 24492 37825 24501 37859
rect 24501 37825 24535 37859
rect 24535 37825 24544 37859
rect 24492 37816 24544 37825
rect 25320 37816 25372 37868
rect 26332 37884 26384 37936
rect 25964 37859 26016 37868
rect 25964 37825 25973 37859
rect 25973 37825 26007 37859
rect 26007 37825 26016 37859
rect 25964 37816 26016 37825
rect 26976 37859 27028 37868
rect 26976 37825 26985 37859
rect 26985 37825 27019 37859
rect 27019 37825 27028 37859
rect 26976 37816 27028 37825
rect 27436 37952 27488 38004
rect 27252 37859 27304 37868
rect 27252 37825 27261 37859
rect 27261 37825 27295 37859
rect 27295 37825 27304 37859
rect 27252 37816 27304 37825
rect 27344 37859 27396 37902
rect 27344 37850 27361 37859
rect 27361 37850 27395 37859
rect 27395 37850 27396 37859
rect 27620 37816 27672 37868
rect 22928 37748 22980 37800
rect 25872 37748 25924 37800
rect 27804 37748 27856 37800
rect 31116 37952 31168 38004
rect 29552 37884 29604 37936
rect 30656 37884 30708 37936
rect 29552 37748 29604 37800
rect 29644 37748 29696 37800
rect 13268 37612 13320 37664
rect 15476 37612 15528 37664
rect 15752 37655 15804 37664
rect 15752 37621 15761 37655
rect 15761 37621 15795 37655
rect 15795 37621 15804 37655
rect 15752 37612 15804 37621
rect 18052 37612 18104 37664
rect 18420 37655 18472 37664
rect 18420 37621 18429 37655
rect 18429 37621 18463 37655
rect 18463 37621 18472 37655
rect 18420 37612 18472 37621
rect 23296 37655 23348 37664
rect 23296 37621 23305 37655
rect 23305 37621 23339 37655
rect 23339 37621 23348 37655
rect 23296 37612 23348 37621
rect 24400 37612 24452 37664
rect 28724 37612 28776 37664
rect 29000 37612 29052 37664
rect 31300 37655 31352 37664
rect 31300 37621 31309 37655
rect 31309 37621 31343 37655
rect 31343 37621 31352 37655
rect 31300 37612 31352 37621
rect 2136 37510 2188 37562
rect 12440 37510 12492 37562
rect 22744 37510 22796 37562
rect 2780 37451 2832 37460
rect 2780 37417 2789 37451
rect 2789 37417 2823 37451
rect 2823 37417 2832 37451
rect 7564 37451 7616 37460
rect 2780 37408 2832 37417
rect 7564 37417 7573 37451
rect 7573 37417 7607 37451
rect 7607 37417 7616 37451
rect 7564 37408 7616 37417
rect 12348 37408 12400 37460
rect 13084 37408 13136 37460
rect 13636 37408 13688 37460
rect 15936 37408 15988 37460
rect 20536 37408 20588 37460
rect 23296 37408 23348 37460
rect 23480 37408 23532 37460
rect 6828 37340 6880 37392
rect 6092 37315 6144 37324
rect 1400 37247 1452 37256
rect 1400 37213 1409 37247
rect 1409 37213 1443 37247
rect 1443 37213 1452 37247
rect 1400 37204 1452 37213
rect 4344 37247 4396 37256
rect 4344 37213 4353 37247
rect 4353 37213 4387 37247
rect 4387 37213 4396 37247
rect 4344 37204 4396 37213
rect 1308 37136 1360 37188
rect 1492 37136 1544 37188
rect 3240 37136 3292 37188
rect 5724 37204 5776 37256
rect 6092 37281 6101 37315
rect 6101 37281 6135 37315
rect 6135 37281 6144 37315
rect 6092 37272 6144 37281
rect 11704 37340 11756 37392
rect 13360 37340 13412 37392
rect 8024 37315 8076 37324
rect 8024 37281 8033 37315
rect 8033 37281 8067 37315
rect 8067 37281 8076 37315
rect 8024 37272 8076 37281
rect 8116 37272 8168 37324
rect 11888 37272 11940 37324
rect 4712 37179 4764 37188
rect 4712 37145 4721 37179
rect 4721 37145 4755 37179
rect 4755 37145 4764 37179
rect 4712 37136 4764 37145
rect 6460 37204 6512 37256
rect 7012 37247 7064 37256
rect 7012 37213 7021 37247
rect 7021 37213 7055 37247
rect 7055 37213 7064 37247
rect 7748 37247 7800 37256
rect 7012 37204 7064 37213
rect 7748 37213 7757 37247
rect 7757 37213 7791 37247
rect 7791 37213 7800 37247
rect 7748 37204 7800 37213
rect 8944 37204 8996 37256
rect 9220 37247 9272 37256
rect 8668 37136 8720 37188
rect 9220 37213 9229 37247
rect 9229 37213 9263 37247
rect 9263 37213 9272 37247
rect 9220 37204 9272 37213
rect 9404 37204 9456 37256
rect 10048 37136 10100 37188
rect 6276 37068 6328 37120
rect 6644 37111 6696 37120
rect 6644 37077 6653 37111
rect 6653 37077 6687 37111
rect 6687 37077 6696 37111
rect 6644 37068 6696 37077
rect 7104 37068 7156 37120
rect 10324 37111 10376 37120
rect 10324 37077 10333 37111
rect 10333 37077 10367 37111
rect 10367 37077 10376 37111
rect 10324 37068 10376 37077
rect 10692 37204 10744 37256
rect 11520 37179 11572 37188
rect 11520 37145 11529 37179
rect 11529 37145 11563 37179
rect 11563 37145 11572 37179
rect 11520 37136 11572 37145
rect 11244 37068 11296 37120
rect 12072 37204 12124 37256
rect 14556 37247 14608 37256
rect 11980 37136 12032 37188
rect 13820 37136 13872 37188
rect 14556 37213 14565 37247
rect 14565 37213 14599 37247
rect 14599 37213 14608 37247
rect 14556 37204 14608 37213
rect 14648 37247 14700 37256
rect 14648 37213 14658 37247
rect 14658 37213 14692 37247
rect 14692 37213 14700 37247
rect 14924 37340 14976 37392
rect 15292 37340 15344 37392
rect 16488 37340 16540 37392
rect 19156 37340 19208 37392
rect 24676 37408 24728 37460
rect 27068 37408 27120 37460
rect 27160 37408 27212 37460
rect 24584 37340 24636 37392
rect 26240 37340 26292 37392
rect 27252 37340 27304 37392
rect 27620 37340 27672 37392
rect 28724 37340 28776 37392
rect 15660 37315 15712 37324
rect 15660 37281 15669 37315
rect 15669 37281 15703 37315
rect 15703 37281 15712 37315
rect 15660 37272 15712 37281
rect 19708 37272 19760 37324
rect 21732 37272 21784 37324
rect 24216 37272 24268 37324
rect 14648 37204 14700 37213
rect 15200 37204 15252 37256
rect 15292 37204 15344 37256
rect 17776 37247 17828 37256
rect 17776 37213 17785 37247
rect 17785 37213 17819 37247
rect 17819 37213 17828 37247
rect 17776 37204 17828 37213
rect 17868 37204 17920 37256
rect 18236 37247 18288 37256
rect 18236 37213 18245 37247
rect 18245 37213 18279 37247
rect 18279 37213 18288 37247
rect 18236 37204 18288 37213
rect 18420 37247 18472 37256
rect 18420 37213 18441 37247
rect 18441 37213 18472 37247
rect 18420 37204 18472 37213
rect 14832 37179 14884 37188
rect 14832 37145 14841 37179
rect 14841 37145 14875 37179
rect 14875 37145 14884 37179
rect 14832 37136 14884 37145
rect 17316 37136 17368 37188
rect 19984 37204 20036 37256
rect 20996 37247 21048 37256
rect 20996 37213 21005 37247
rect 21005 37213 21039 37247
rect 21039 37213 21048 37247
rect 20996 37204 21048 37213
rect 21548 37204 21600 37256
rect 23020 37247 23072 37256
rect 15844 37068 15896 37120
rect 16948 37068 17000 37120
rect 17684 37068 17736 37120
rect 23020 37213 23029 37247
rect 23029 37213 23063 37247
rect 23063 37213 23072 37247
rect 23020 37204 23072 37213
rect 24032 37204 24084 37256
rect 25964 37247 26016 37256
rect 23388 37136 23440 37188
rect 25964 37213 25973 37247
rect 25973 37213 26007 37247
rect 26007 37213 26016 37247
rect 25964 37204 26016 37213
rect 26056 37204 26108 37256
rect 24768 37136 24820 37188
rect 26792 37204 26844 37256
rect 27436 37204 27488 37256
rect 27988 37272 28040 37324
rect 29184 37408 29236 37460
rect 29828 37408 29880 37460
rect 29736 37340 29788 37392
rect 28816 37247 28868 37256
rect 28816 37213 28825 37247
rect 28825 37213 28859 37247
rect 28859 37213 28868 37247
rect 28816 37204 28868 37213
rect 29000 37247 29052 37256
rect 29000 37213 29021 37247
rect 29021 37213 29052 37247
rect 29000 37204 29052 37213
rect 24032 37068 24084 37120
rect 25596 37068 25648 37120
rect 27620 37179 27672 37188
rect 27620 37145 27629 37179
rect 27629 37145 27663 37179
rect 27663 37145 27672 37179
rect 27620 37136 27672 37145
rect 27804 37136 27856 37188
rect 30104 37136 30156 37188
rect 27160 37068 27212 37120
rect 28954 37068 29006 37120
rect 29644 37068 29696 37120
rect 7288 36966 7340 37018
rect 17592 36966 17644 37018
rect 27896 36966 27948 37018
rect 1492 36864 1544 36916
rect 3792 36864 3844 36916
rect 4344 36864 4396 36916
rect 2872 36728 2924 36780
rect 3792 36771 3844 36780
rect 3792 36737 3801 36771
rect 3801 36737 3835 36771
rect 3835 36737 3844 36771
rect 3792 36728 3844 36737
rect 4160 36728 4212 36780
rect 4344 36728 4396 36780
rect 4620 36728 4672 36780
rect 3240 36660 3292 36712
rect 5632 36728 5684 36780
rect 5356 36660 5408 36712
rect 8392 36864 8444 36916
rect 6828 36796 6880 36848
rect 6552 36771 6604 36780
rect 6552 36737 6561 36771
rect 6561 36737 6595 36771
rect 6595 36737 6604 36771
rect 6552 36728 6604 36737
rect 6828 36703 6880 36712
rect 6828 36669 6837 36703
rect 6837 36669 6871 36703
rect 6871 36669 6880 36703
rect 6828 36660 6880 36669
rect 3332 36592 3384 36644
rect 7012 36592 7064 36644
rect 9220 36796 9272 36848
rect 10324 36864 10376 36916
rect 12256 36864 12308 36916
rect 14372 36864 14424 36916
rect 14556 36864 14608 36916
rect 15752 36907 15804 36916
rect 15752 36873 15761 36907
rect 15761 36873 15795 36907
rect 15795 36873 15804 36907
rect 15752 36864 15804 36873
rect 15844 36907 15896 36916
rect 15844 36873 15853 36907
rect 15853 36873 15887 36907
rect 15887 36873 15896 36907
rect 15844 36864 15896 36873
rect 18512 36907 18564 36916
rect 18512 36873 18521 36907
rect 18521 36873 18555 36907
rect 18555 36873 18564 36907
rect 18512 36864 18564 36873
rect 19064 36864 19116 36916
rect 19984 36864 20036 36916
rect 20904 36864 20956 36916
rect 21180 36864 21232 36916
rect 8668 36771 8720 36780
rect 8668 36737 8677 36771
rect 8677 36737 8711 36771
rect 8711 36737 8720 36771
rect 8668 36728 8720 36737
rect 9588 36771 9640 36780
rect 9588 36737 9597 36771
rect 9597 36737 9631 36771
rect 9631 36737 9640 36771
rect 9588 36728 9640 36737
rect 15292 36796 15344 36848
rect 11060 36728 11112 36780
rect 11612 36728 11664 36780
rect 11796 36728 11848 36780
rect 12532 36728 12584 36780
rect 13084 36771 13136 36780
rect 13084 36737 13093 36771
rect 13093 36737 13127 36771
rect 13127 36737 13136 36771
rect 13084 36728 13136 36737
rect 13268 36771 13320 36780
rect 13268 36737 13277 36771
rect 13277 36737 13311 36771
rect 13311 36737 13320 36771
rect 13268 36728 13320 36737
rect 9128 36660 9180 36712
rect 9312 36660 9364 36712
rect 13452 36728 13504 36780
rect 14280 36771 14332 36780
rect 14280 36737 14289 36771
rect 14289 36737 14323 36771
rect 14323 36737 14332 36771
rect 14280 36728 14332 36737
rect 14464 36771 14516 36780
rect 14464 36737 14473 36771
rect 14473 36737 14507 36771
rect 14507 36737 14516 36771
rect 14464 36728 14516 36737
rect 14924 36728 14976 36780
rect 16672 36771 16724 36780
rect 16672 36737 16681 36771
rect 16681 36737 16715 36771
rect 16715 36737 16724 36771
rect 16672 36728 16724 36737
rect 16948 36771 17000 36780
rect 16948 36737 16957 36771
rect 16957 36737 16991 36771
rect 16991 36737 17000 36771
rect 16948 36728 17000 36737
rect 10232 36592 10284 36644
rect 14556 36660 14608 36712
rect 15660 36660 15712 36712
rect 17040 36660 17092 36712
rect 23388 36796 23440 36848
rect 17776 36728 17828 36780
rect 17500 36660 17552 36712
rect 18052 36660 18104 36712
rect 17684 36592 17736 36644
rect 19248 36771 19300 36780
rect 18236 36660 18288 36712
rect 19248 36737 19257 36771
rect 19257 36737 19291 36771
rect 19291 36737 19300 36771
rect 19248 36728 19300 36737
rect 19524 36728 19576 36780
rect 21180 36728 21232 36780
rect 22652 36728 22704 36780
rect 23020 36728 23072 36780
rect 25228 36771 25280 36780
rect 25228 36737 25237 36771
rect 25237 36737 25271 36771
rect 25271 36737 25280 36771
rect 25228 36728 25280 36737
rect 27344 36864 27396 36916
rect 28816 36864 28868 36916
rect 30288 36864 30340 36916
rect 26148 36771 26200 36780
rect 26148 36737 26157 36771
rect 26157 36737 26191 36771
rect 26191 36737 26200 36771
rect 26148 36728 26200 36737
rect 27160 36728 27212 36780
rect 29000 36796 29052 36848
rect 30012 36796 30064 36848
rect 22376 36660 22428 36712
rect 24032 36660 24084 36712
rect 26792 36660 26844 36712
rect 29276 36771 29328 36780
rect 29276 36737 29285 36771
rect 29285 36737 29319 36771
rect 29319 36737 29328 36771
rect 29276 36728 29328 36737
rect 29736 36728 29788 36780
rect 19248 36592 19300 36644
rect 21364 36592 21416 36644
rect 25596 36592 25648 36644
rect 2228 36524 2280 36576
rect 2412 36524 2464 36576
rect 6368 36567 6420 36576
rect 6368 36533 6377 36567
rect 6377 36533 6411 36567
rect 6411 36533 6420 36567
rect 6368 36524 6420 36533
rect 8116 36524 8168 36576
rect 8392 36524 8444 36576
rect 11704 36524 11756 36576
rect 13544 36524 13596 36576
rect 15384 36567 15436 36576
rect 15384 36533 15393 36567
rect 15393 36533 15427 36567
rect 15427 36533 15436 36567
rect 15384 36524 15436 36533
rect 15752 36524 15804 36576
rect 17408 36567 17460 36576
rect 17408 36533 17417 36567
rect 17417 36533 17451 36567
rect 17451 36533 17460 36567
rect 17408 36524 17460 36533
rect 19156 36524 19208 36576
rect 19708 36524 19760 36576
rect 21180 36524 21232 36576
rect 21916 36567 21968 36576
rect 21916 36533 21925 36567
rect 21925 36533 21959 36567
rect 21959 36533 21968 36567
rect 21916 36524 21968 36533
rect 24676 36524 24728 36576
rect 26056 36524 26108 36576
rect 26792 36524 26844 36576
rect 27436 36524 27488 36576
rect 31300 36728 31352 36780
rect 28908 36592 28960 36644
rect 31024 36592 31076 36644
rect 28632 36567 28684 36576
rect 28632 36533 28641 36567
rect 28641 36533 28675 36567
rect 28675 36533 28684 36567
rect 28632 36524 28684 36533
rect 29552 36524 29604 36576
rect 2136 36422 2188 36474
rect 12440 36422 12492 36474
rect 22744 36422 22796 36474
rect 2504 36320 2556 36372
rect 4620 36320 4672 36372
rect 6276 36320 6328 36372
rect 2596 36252 2648 36304
rect 5448 36184 5500 36236
rect 8392 36363 8444 36372
rect 8392 36329 8401 36363
rect 8401 36329 8435 36363
rect 8435 36329 8444 36363
rect 8392 36320 8444 36329
rect 9128 36320 9180 36372
rect 10324 36320 10376 36372
rect 10692 36320 10744 36372
rect 10784 36320 10836 36372
rect 11060 36320 11112 36372
rect 11612 36252 11664 36304
rect 9312 36227 9364 36236
rect 3240 36116 3292 36168
rect 3792 36116 3844 36168
rect 4160 36116 4212 36168
rect 4712 36116 4764 36168
rect 5172 36116 5224 36168
rect 6644 36116 6696 36168
rect 9312 36193 9321 36227
rect 9321 36193 9355 36227
rect 9355 36193 9364 36227
rect 9312 36184 9364 36193
rect 9588 36184 9640 36236
rect 10968 36227 11020 36236
rect 9404 36116 9456 36168
rect 9680 36116 9732 36168
rect 10692 36159 10744 36168
rect 10692 36125 10701 36159
rect 10701 36125 10735 36159
rect 10735 36125 10744 36159
rect 10692 36116 10744 36125
rect 10968 36193 10977 36227
rect 10977 36193 11011 36227
rect 11011 36193 11020 36227
rect 10968 36184 11020 36193
rect 11428 36159 11480 36168
rect 11428 36125 11437 36159
rect 11437 36125 11471 36159
rect 11471 36125 11480 36159
rect 11428 36116 11480 36125
rect 22192 36320 22244 36372
rect 24768 36320 24820 36372
rect 26148 36320 26200 36372
rect 28908 36363 28960 36372
rect 13268 36252 13320 36304
rect 14280 36252 14332 36304
rect 15200 36252 15252 36304
rect 16672 36252 16724 36304
rect 17776 36295 17828 36304
rect 17776 36261 17785 36295
rect 17785 36261 17819 36295
rect 17819 36261 17828 36295
rect 17776 36252 17828 36261
rect 27344 36252 27396 36304
rect 2044 35980 2096 36032
rect 2964 35980 3016 36032
rect 4620 35980 4672 36032
rect 7012 35980 7064 36032
rect 10324 35980 10376 36032
rect 10508 36023 10560 36032
rect 10508 35989 10517 36023
rect 10517 35989 10551 36023
rect 10551 35989 10560 36023
rect 10508 35980 10560 35989
rect 11060 36048 11112 36100
rect 13176 36116 13228 36168
rect 14004 36116 14056 36168
rect 14556 36159 14608 36168
rect 14556 36125 14565 36159
rect 14565 36125 14599 36159
rect 14599 36125 14608 36159
rect 14556 36116 14608 36125
rect 14648 36116 14700 36168
rect 15752 36159 15804 36168
rect 15752 36125 15761 36159
rect 15761 36125 15795 36159
rect 15795 36125 15804 36159
rect 15752 36116 15804 36125
rect 16580 36116 16632 36168
rect 17500 36184 17552 36236
rect 16948 36159 17000 36168
rect 16948 36125 16957 36159
rect 16957 36125 16991 36159
rect 16991 36125 17000 36159
rect 16948 36116 17000 36125
rect 17040 36159 17092 36168
rect 17040 36125 17049 36159
rect 17049 36125 17083 36159
rect 17083 36125 17092 36159
rect 17040 36116 17092 36125
rect 17868 36116 17920 36168
rect 19524 36184 19576 36236
rect 18236 36159 18288 36168
rect 18236 36125 18245 36159
rect 18245 36125 18279 36159
rect 18279 36125 18288 36159
rect 18236 36116 18288 36125
rect 18328 36116 18380 36168
rect 13360 36048 13412 36100
rect 19984 36116 20036 36168
rect 20812 36159 20864 36168
rect 20812 36125 20821 36159
rect 20821 36125 20855 36159
rect 20855 36125 20864 36159
rect 20812 36116 20864 36125
rect 22560 36116 22612 36168
rect 22652 36159 22704 36168
rect 22652 36125 22661 36159
rect 22661 36125 22695 36159
rect 22695 36125 22704 36159
rect 22652 36116 22704 36125
rect 23480 36116 23532 36168
rect 24952 36184 25004 36236
rect 25780 36227 25832 36236
rect 25780 36193 25789 36227
rect 25789 36193 25823 36227
rect 25823 36193 25832 36227
rect 25780 36184 25832 36193
rect 26792 36184 26844 36236
rect 28908 36329 28917 36363
rect 28917 36329 28951 36363
rect 28951 36329 28960 36363
rect 28908 36320 28960 36329
rect 29552 36227 29604 36236
rect 29552 36193 29561 36227
rect 29561 36193 29595 36227
rect 29595 36193 29604 36227
rect 29552 36184 29604 36193
rect 24860 36159 24912 36168
rect 21916 36048 21968 36100
rect 22284 36048 22336 36100
rect 23204 36048 23256 36100
rect 24860 36125 24869 36159
rect 24869 36125 24903 36159
rect 24903 36125 24912 36159
rect 24860 36116 24912 36125
rect 25136 36048 25188 36100
rect 12072 35980 12124 36032
rect 15844 35980 15896 36032
rect 16028 35980 16080 36032
rect 19156 35980 19208 36032
rect 19524 35980 19576 36032
rect 21548 35980 21600 36032
rect 23848 35980 23900 36032
rect 27160 36116 27212 36168
rect 26056 36091 26108 36100
rect 26056 36057 26090 36091
rect 26090 36057 26108 36091
rect 26056 36048 26108 36057
rect 27436 36048 27488 36100
rect 26516 35980 26568 36032
rect 28540 36116 28592 36168
rect 28632 36116 28684 36168
rect 28264 35980 28316 36032
rect 30840 35980 30892 36032
rect 7288 35878 7340 35930
rect 17592 35878 17644 35930
rect 27896 35878 27948 35930
rect 3240 35776 3292 35828
rect 2228 35708 2280 35760
rect 3332 35708 3384 35760
rect 10600 35776 10652 35828
rect 11520 35776 11572 35828
rect 6460 35708 6512 35760
rect 1400 35683 1452 35692
rect 1400 35649 1409 35683
rect 1409 35649 1443 35683
rect 1443 35649 1452 35683
rect 1400 35640 1452 35649
rect 1676 35683 1728 35692
rect 1676 35649 1710 35683
rect 1710 35649 1728 35683
rect 1676 35640 1728 35649
rect 7012 35683 7064 35692
rect 7012 35649 7021 35683
rect 7021 35649 7055 35683
rect 7055 35649 7064 35683
rect 7012 35640 7064 35649
rect 9864 35708 9916 35760
rect 9956 35708 10008 35760
rect 13360 35751 13412 35760
rect 8944 35640 8996 35692
rect 9680 35640 9732 35692
rect 10876 35640 10928 35692
rect 11060 35640 11112 35692
rect 11612 35640 11664 35692
rect 13360 35717 13369 35751
rect 13369 35717 13403 35751
rect 13403 35717 13412 35751
rect 13360 35708 13412 35717
rect 13452 35708 13504 35760
rect 14648 35708 14700 35760
rect 13544 35683 13596 35692
rect 6920 35572 6972 35624
rect 9036 35572 9088 35624
rect 9588 35572 9640 35624
rect 11520 35615 11572 35624
rect 11520 35581 11529 35615
rect 11529 35581 11563 35615
rect 11563 35581 11572 35615
rect 11520 35572 11572 35581
rect 7012 35504 7064 35556
rect 10048 35504 10100 35556
rect 13544 35649 13553 35683
rect 13553 35649 13587 35683
rect 13587 35649 13596 35683
rect 13544 35640 13596 35649
rect 13728 35683 13780 35692
rect 13728 35649 13737 35683
rect 13737 35649 13771 35683
rect 13771 35649 13780 35683
rect 13728 35640 13780 35649
rect 15108 35708 15160 35760
rect 20812 35776 20864 35828
rect 15844 35751 15896 35760
rect 15844 35717 15853 35751
rect 15853 35717 15887 35751
rect 15887 35717 15896 35751
rect 15844 35708 15896 35717
rect 15568 35640 15620 35692
rect 16856 35683 16908 35692
rect 16856 35649 16865 35683
rect 16865 35649 16899 35683
rect 16899 35649 16908 35683
rect 16856 35640 16908 35649
rect 17408 35640 17460 35692
rect 15660 35572 15712 35624
rect 15936 35615 15988 35624
rect 15936 35581 15945 35615
rect 15945 35581 15979 35615
rect 15979 35581 15988 35615
rect 15936 35572 15988 35581
rect 19248 35640 19300 35692
rect 20904 35683 20956 35692
rect 20904 35649 20913 35683
rect 20913 35649 20947 35683
rect 20947 35649 20956 35683
rect 20904 35640 20956 35649
rect 21548 35640 21600 35692
rect 21732 35640 21784 35692
rect 23020 35640 23072 35692
rect 24952 35708 25004 35760
rect 25044 35708 25096 35760
rect 24676 35683 24728 35692
rect 24676 35649 24710 35683
rect 24710 35649 24728 35683
rect 24676 35640 24728 35649
rect 26608 35640 26660 35692
rect 27160 35683 27212 35692
rect 27160 35649 27169 35683
rect 27169 35649 27203 35683
rect 27203 35649 27212 35683
rect 27160 35640 27212 35649
rect 3792 35436 3844 35488
rect 9220 35436 9272 35488
rect 12900 35479 12952 35488
rect 12900 35445 12909 35479
rect 12909 35445 12943 35479
rect 12943 35445 12952 35479
rect 12900 35436 12952 35445
rect 15200 35436 15252 35488
rect 15292 35436 15344 35488
rect 21180 35572 21232 35624
rect 21640 35572 21692 35624
rect 21548 35504 21600 35556
rect 23848 35547 23900 35556
rect 23848 35513 23857 35547
rect 23857 35513 23891 35547
rect 23891 35513 23900 35547
rect 23848 35504 23900 35513
rect 18236 35479 18288 35488
rect 18236 35445 18245 35479
rect 18245 35445 18279 35479
rect 18279 35445 18288 35479
rect 18236 35436 18288 35445
rect 18696 35436 18748 35488
rect 19984 35436 20036 35488
rect 21640 35436 21692 35488
rect 22376 35436 22428 35488
rect 25044 35436 25096 35488
rect 25136 35436 25188 35488
rect 27344 35708 27396 35760
rect 27436 35683 27488 35692
rect 27436 35649 27445 35683
rect 27445 35649 27479 35683
rect 27479 35649 27488 35683
rect 27436 35640 27488 35649
rect 28540 35708 28592 35760
rect 28172 35683 28224 35692
rect 28172 35649 28181 35683
rect 28181 35649 28215 35683
rect 28215 35649 28224 35683
rect 28172 35640 28224 35649
rect 29276 35683 29328 35692
rect 28448 35572 28500 35624
rect 29276 35649 29285 35683
rect 29285 35649 29319 35683
rect 29319 35649 29328 35683
rect 29276 35640 29328 35649
rect 29460 35683 29512 35692
rect 29460 35649 29469 35683
rect 29469 35649 29503 35683
rect 29503 35649 29512 35683
rect 29460 35640 29512 35649
rect 29736 35572 29788 35624
rect 27252 35504 27304 35556
rect 25780 35479 25832 35488
rect 25780 35445 25789 35479
rect 25789 35445 25823 35479
rect 25823 35445 25832 35479
rect 25780 35436 25832 35445
rect 26332 35436 26384 35488
rect 28080 35436 28132 35488
rect 28264 35479 28316 35488
rect 28264 35445 28273 35479
rect 28273 35445 28307 35479
rect 28307 35445 28316 35479
rect 28264 35436 28316 35445
rect 29000 35504 29052 35556
rect 29552 35504 29604 35556
rect 31300 35479 31352 35488
rect 31300 35445 31309 35479
rect 31309 35445 31343 35479
rect 31343 35445 31352 35479
rect 31300 35436 31352 35445
rect 2136 35334 2188 35386
rect 12440 35334 12492 35386
rect 22744 35334 22796 35386
rect 1676 35232 1728 35284
rect 2228 35275 2280 35284
rect 2228 35241 2237 35275
rect 2237 35241 2271 35275
rect 2271 35241 2280 35275
rect 2228 35232 2280 35241
rect 5080 35232 5132 35284
rect 6552 35232 6604 35284
rect 8944 35275 8996 35284
rect 8944 35241 8953 35275
rect 8953 35241 8987 35275
rect 8987 35241 8996 35275
rect 8944 35232 8996 35241
rect 12900 35232 12952 35284
rect 14924 35275 14976 35284
rect 14924 35241 14933 35275
rect 14933 35241 14967 35275
rect 14967 35241 14976 35275
rect 14924 35232 14976 35241
rect 15568 35275 15620 35284
rect 15568 35241 15577 35275
rect 15577 35241 15611 35275
rect 15611 35241 15620 35275
rect 15568 35232 15620 35241
rect 16948 35232 17000 35284
rect 17868 35232 17920 35284
rect 19248 35275 19300 35284
rect 2688 35096 2740 35148
rect 3792 35139 3844 35148
rect 3792 35105 3801 35139
rect 3801 35105 3835 35139
rect 3835 35105 3844 35139
rect 3792 35096 3844 35105
rect 2044 35071 2096 35080
rect 2044 35037 2053 35071
rect 2053 35037 2087 35071
rect 2087 35037 2096 35071
rect 2044 35028 2096 35037
rect 2964 35071 3016 35080
rect 2964 35037 2973 35071
rect 2973 35037 3007 35071
rect 3007 35037 3016 35071
rect 2964 35028 3016 35037
rect 4344 35028 4396 35080
rect 8116 35164 8168 35216
rect 10968 35164 11020 35216
rect 13544 35207 13596 35216
rect 13544 35173 13553 35207
rect 13553 35173 13587 35207
rect 13587 35173 13596 35207
rect 13544 35164 13596 35173
rect 16028 35164 16080 35216
rect 18696 35164 18748 35216
rect 19248 35241 19257 35275
rect 19257 35241 19291 35275
rect 19291 35241 19300 35275
rect 19248 35232 19300 35241
rect 19340 35232 19392 35284
rect 19432 35164 19484 35216
rect 20812 35164 20864 35216
rect 21456 35164 21508 35216
rect 22008 35232 22060 35284
rect 22100 35232 22152 35284
rect 23020 35275 23072 35284
rect 23020 35241 23029 35275
rect 23029 35241 23063 35275
rect 23063 35241 23072 35275
rect 23020 35232 23072 35241
rect 25228 35232 25280 35284
rect 26056 35275 26108 35284
rect 26056 35241 26065 35275
rect 26065 35241 26099 35275
rect 26099 35241 26108 35275
rect 26056 35232 26108 35241
rect 26148 35232 26200 35284
rect 7012 35096 7064 35148
rect 6920 35071 6972 35080
rect 6920 35037 6929 35071
rect 6929 35037 6963 35071
rect 6963 35037 6972 35071
rect 6920 35028 6972 35037
rect 7104 35071 7156 35080
rect 7104 35037 7113 35071
rect 7113 35037 7147 35071
rect 7147 35037 7156 35071
rect 7104 35028 7156 35037
rect 7932 35028 7984 35080
rect 1952 34960 2004 35012
rect 8300 35028 8352 35080
rect 9128 35071 9180 35080
rect 9128 35037 9137 35071
rect 9137 35037 9171 35071
rect 9171 35037 9180 35071
rect 9128 35028 9180 35037
rect 9864 35071 9916 35080
rect 9864 35037 9873 35071
rect 9873 35037 9907 35071
rect 9907 35037 9916 35071
rect 11888 35096 11940 35148
rect 14556 35139 14608 35148
rect 14556 35105 14565 35139
rect 14565 35105 14599 35139
rect 14599 35105 14608 35139
rect 14556 35096 14608 35105
rect 9864 35028 9916 35037
rect 9404 34960 9456 35012
rect 9588 34960 9640 35012
rect 10508 34960 10560 35012
rect 10784 34960 10836 35012
rect 15384 35071 15436 35080
rect 13360 35003 13412 35012
rect 13360 34969 13369 35003
rect 13369 34969 13403 35003
rect 13403 34969 13412 35003
rect 13360 34960 13412 34969
rect 14648 34960 14700 35012
rect 15384 35037 15393 35071
rect 15393 35037 15427 35071
rect 15427 35037 15436 35071
rect 15384 35028 15436 35037
rect 2780 34935 2832 34944
rect 2780 34901 2789 34935
rect 2789 34901 2823 34935
rect 2823 34901 2832 34935
rect 2780 34892 2832 34901
rect 6920 34892 6972 34944
rect 7472 34892 7524 34944
rect 7748 34892 7800 34944
rect 11060 34892 11112 34944
rect 12256 34935 12308 34944
rect 12256 34901 12265 34935
rect 12265 34901 12299 34935
rect 12299 34901 12308 34935
rect 12256 34892 12308 34901
rect 13084 34892 13136 34944
rect 16396 34960 16448 35012
rect 15384 34892 15436 34944
rect 16488 34892 16540 34944
rect 16672 35028 16724 35080
rect 17132 35028 17184 35080
rect 17960 35028 18012 35080
rect 18880 35028 18932 35080
rect 20904 35096 20956 35148
rect 22652 35164 22704 35216
rect 23112 35164 23164 35216
rect 26240 35164 26292 35216
rect 27252 35164 27304 35216
rect 29184 35232 29236 35284
rect 29460 35232 29512 35284
rect 29276 35164 29328 35216
rect 25964 35096 26016 35148
rect 19524 35028 19576 35080
rect 20168 35071 20220 35080
rect 17500 34960 17552 35012
rect 20168 35037 20177 35071
rect 20177 35037 20211 35071
rect 20211 35037 20220 35071
rect 20168 35028 20220 35037
rect 18236 34892 18288 34944
rect 19156 34892 19208 34944
rect 20076 34892 20128 34944
rect 21180 35071 21232 35080
rect 21180 35037 21189 35071
rect 21189 35037 21223 35071
rect 21223 35037 21232 35071
rect 21180 35028 21232 35037
rect 21364 35028 21416 35080
rect 21640 35028 21692 35080
rect 23204 35071 23256 35080
rect 23204 35037 23213 35071
rect 23213 35037 23247 35071
rect 23247 35037 23256 35071
rect 23204 35028 23256 35037
rect 23664 35028 23716 35080
rect 25136 35071 25188 35080
rect 25136 35037 25145 35071
rect 25145 35037 25179 35071
rect 25179 35037 25188 35071
rect 25136 35028 25188 35037
rect 22284 34960 22336 35012
rect 24860 34960 24912 35012
rect 25228 34960 25280 35012
rect 25504 35028 25556 35080
rect 25780 35028 25832 35080
rect 26332 35028 26384 35080
rect 26516 35071 26568 35080
rect 26516 35037 26525 35071
rect 26525 35037 26559 35071
rect 26559 35037 26568 35071
rect 26516 35028 26568 35037
rect 26792 35028 26844 35080
rect 27436 34960 27488 35012
rect 28724 35096 28776 35148
rect 29000 35028 29052 35080
rect 30196 35028 30248 35080
rect 30932 35071 30984 35080
rect 30932 35037 30941 35071
rect 30941 35037 30975 35071
rect 30975 35037 30984 35071
rect 30932 35028 30984 35037
rect 31300 35028 31352 35080
rect 28080 34960 28132 35012
rect 20352 34892 20404 34944
rect 25320 34892 25372 34944
rect 27160 34892 27212 34944
rect 7288 34790 7340 34842
rect 17592 34790 17644 34842
rect 27896 34790 27948 34842
rect 5172 34731 5224 34740
rect 2780 34620 2832 34672
rect 5172 34697 5181 34731
rect 5181 34697 5215 34731
rect 5215 34697 5224 34731
rect 5172 34688 5224 34697
rect 7012 34688 7064 34740
rect 7104 34688 7156 34740
rect 8024 34688 8076 34740
rect 10416 34688 10468 34740
rect 10784 34688 10836 34740
rect 10968 34688 11020 34740
rect 11888 34731 11940 34740
rect 11888 34697 11897 34731
rect 11897 34697 11931 34731
rect 11931 34697 11940 34731
rect 11888 34688 11940 34697
rect 14556 34688 14608 34740
rect 15384 34688 15436 34740
rect 15568 34688 15620 34740
rect 20076 34688 20128 34740
rect 21640 34688 21692 34740
rect 6368 34620 6420 34672
rect 8208 34620 8260 34672
rect 8576 34620 8628 34672
rect 5080 34552 5132 34604
rect 5632 34552 5684 34604
rect 5816 34595 5868 34604
rect 5816 34561 5825 34595
rect 5825 34561 5859 34595
rect 5859 34561 5868 34595
rect 5816 34552 5868 34561
rect 9864 34620 9916 34672
rect 11704 34663 11756 34672
rect 11704 34629 11713 34663
rect 11713 34629 11747 34663
rect 11747 34629 11756 34663
rect 11704 34620 11756 34629
rect 12256 34620 12308 34672
rect 15292 34620 15344 34672
rect 10048 34552 10100 34604
rect 13544 34552 13596 34604
rect 14188 34595 14240 34604
rect 6368 34527 6420 34536
rect 2688 34416 2740 34468
rect 6368 34493 6377 34527
rect 6377 34493 6411 34527
rect 6411 34493 6420 34527
rect 6368 34484 6420 34493
rect 12348 34484 12400 34536
rect 13268 34484 13320 34536
rect 13452 34527 13504 34536
rect 13452 34493 13461 34527
rect 13461 34493 13495 34527
rect 13495 34493 13504 34527
rect 14188 34561 14197 34595
rect 14197 34561 14231 34595
rect 14231 34561 14240 34595
rect 14188 34552 14240 34561
rect 14648 34595 14700 34604
rect 14648 34561 14657 34595
rect 14657 34561 14691 34595
rect 14691 34561 14700 34595
rect 14648 34552 14700 34561
rect 15200 34552 15252 34604
rect 15476 34595 15528 34604
rect 15476 34561 15485 34595
rect 15485 34561 15519 34595
rect 15519 34561 15528 34595
rect 15476 34552 15528 34561
rect 15660 34620 15712 34672
rect 13452 34484 13504 34493
rect 14924 34484 14976 34536
rect 16304 34484 16356 34536
rect 16396 34484 16448 34536
rect 17500 34552 17552 34604
rect 17960 34552 18012 34604
rect 18328 34552 18380 34604
rect 18512 34595 18564 34604
rect 18512 34561 18521 34595
rect 18521 34561 18555 34595
rect 18555 34561 18564 34595
rect 18512 34552 18564 34561
rect 19984 34620 20036 34672
rect 20628 34620 20680 34672
rect 20904 34552 20956 34604
rect 22468 34552 22520 34604
rect 15936 34416 15988 34468
rect 21180 34484 21232 34536
rect 28172 34688 28224 34740
rect 25964 34663 26016 34672
rect 23112 34595 23164 34604
rect 23112 34561 23121 34595
rect 23121 34561 23155 34595
rect 23155 34561 23164 34595
rect 23112 34552 23164 34561
rect 23204 34527 23256 34536
rect 17316 34416 17368 34468
rect 23204 34493 23213 34527
rect 23213 34493 23247 34527
rect 23247 34493 23256 34527
rect 23664 34595 23716 34604
rect 23664 34561 23673 34595
rect 23673 34561 23707 34595
rect 23707 34561 23716 34595
rect 23664 34552 23716 34561
rect 25044 34552 25096 34604
rect 25228 34552 25280 34604
rect 25964 34629 25973 34663
rect 25973 34629 26007 34663
rect 26007 34629 26016 34663
rect 25964 34620 26016 34629
rect 25780 34552 25832 34604
rect 26240 34552 26292 34604
rect 28908 34620 28960 34672
rect 27344 34552 27396 34604
rect 23204 34484 23256 34493
rect 28448 34552 28500 34604
rect 30380 34688 30432 34740
rect 30840 34688 30892 34740
rect 29276 34552 29328 34604
rect 29736 34552 29788 34604
rect 30196 34552 30248 34604
rect 1584 34391 1636 34400
rect 1584 34357 1593 34391
rect 1593 34357 1627 34391
rect 1627 34357 1636 34391
rect 1584 34348 1636 34357
rect 2872 34391 2924 34400
rect 2872 34357 2881 34391
rect 2881 34357 2915 34391
rect 2915 34357 2924 34391
rect 2872 34348 2924 34357
rect 3148 34348 3200 34400
rect 10416 34348 10468 34400
rect 15384 34348 15436 34400
rect 18420 34348 18472 34400
rect 19340 34348 19392 34400
rect 20536 34348 20588 34400
rect 22192 34416 22244 34468
rect 23848 34416 23900 34468
rect 29552 34484 29604 34536
rect 29828 34416 29880 34468
rect 30748 34416 30800 34468
rect 22376 34348 22428 34400
rect 23572 34348 23624 34400
rect 24768 34348 24820 34400
rect 2136 34246 2188 34298
rect 12440 34246 12492 34298
rect 22744 34246 22796 34298
rect 1952 34144 2004 34196
rect 2228 34187 2280 34196
rect 2228 34153 2237 34187
rect 2237 34153 2271 34187
rect 2271 34153 2280 34187
rect 2228 34144 2280 34153
rect 5724 34144 5776 34196
rect 6828 34144 6880 34196
rect 9128 34144 9180 34196
rect 10048 34187 10100 34196
rect 10048 34153 10057 34187
rect 10057 34153 10091 34187
rect 10091 34153 10100 34187
rect 10048 34144 10100 34153
rect 10692 34144 10744 34196
rect 14924 34144 14976 34196
rect 15476 34144 15528 34196
rect 2504 34008 2556 34060
rect 2780 34008 2832 34060
rect 3148 34051 3200 34060
rect 3148 34017 3157 34051
rect 3157 34017 3191 34051
rect 3191 34017 3200 34051
rect 3148 34008 3200 34017
rect 6368 34008 6420 34060
rect 8116 34008 8168 34060
rect 2964 33983 3016 33992
rect 2964 33949 2973 33983
rect 2973 33949 3007 33983
rect 3007 33949 3016 33983
rect 2964 33940 3016 33949
rect 3240 33983 3292 33992
rect 3240 33949 3249 33983
rect 3249 33949 3283 33983
rect 3283 33949 3292 33983
rect 3240 33940 3292 33949
rect 4436 33940 4488 33992
rect 18512 34076 18564 34128
rect 21732 34144 21784 34196
rect 23664 34144 23716 34196
rect 25780 34187 25832 34196
rect 25780 34153 25789 34187
rect 25789 34153 25823 34187
rect 25823 34153 25832 34187
rect 25780 34144 25832 34153
rect 20812 34076 20864 34128
rect 16304 34051 16356 34060
rect 7932 33940 7984 33992
rect 9128 33983 9180 33992
rect 9128 33949 9137 33983
rect 9137 33949 9171 33983
rect 9171 33949 9180 33983
rect 9128 33940 9180 33949
rect 9404 33983 9456 33992
rect 9404 33949 9413 33983
rect 9413 33949 9447 33983
rect 9447 33949 9456 33983
rect 9404 33940 9456 33949
rect 10232 33983 10284 33992
rect 2412 33872 2464 33924
rect 2872 33872 2924 33924
rect 7564 33872 7616 33924
rect 9220 33872 9272 33924
rect 10232 33949 10241 33983
rect 10241 33949 10275 33983
rect 10275 33949 10284 33983
rect 10232 33940 10284 33949
rect 11060 33983 11112 33992
rect 11060 33949 11069 33983
rect 11069 33949 11103 33983
rect 11103 33949 11112 33983
rect 11060 33940 11112 33949
rect 11888 33983 11940 33992
rect 11888 33949 11897 33983
rect 11897 33949 11931 33983
rect 11931 33949 11940 33983
rect 11888 33940 11940 33949
rect 11980 33983 12032 33992
rect 11980 33949 11989 33983
rect 11989 33949 12023 33983
rect 12023 33949 12032 33983
rect 12992 33983 13044 33992
rect 11980 33940 12032 33949
rect 12992 33949 13001 33983
rect 13001 33949 13035 33983
rect 13035 33949 13044 33983
rect 12992 33940 13044 33949
rect 14188 33940 14240 33992
rect 14464 33983 14516 33992
rect 14464 33949 14473 33983
rect 14473 33949 14507 33983
rect 14507 33949 14516 33983
rect 14464 33940 14516 33949
rect 15476 33940 15528 33992
rect 15660 33983 15712 33992
rect 15660 33949 15669 33983
rect 15669 33949 15703 33983
rect 15703 33949 15712 33983
rect 15660 33940 15712 33949
rect 16304 34017 16313 34051
rect 16313 34017 16347 34051
rect 16347 34017 16356 34051
rect 16304 34008 16356 34017
rect 18696 34051 18748 34060
rect 18696 34017 18705 34051
rect 18705 34017 18739 34051
rect 18739 34017 18748 34051
rect 18696 34008 18748 34017
rect 29000 34144 29052 34196
rect 28540 34119 28592 34128
rect 28540 34085 28549 34119
rect 28549 34085 28583 34119
rect 28583 34085 28592 34119
rect 28540 34076 28592 34085
rect 28908 34119 28960 34128
rect 28908 34085 28917 34119
rect 28917 34085 28951 34119
rect 28951 34085 28960 34119
rect 28908 34076 28960 34085
rect 15936 33940 15988 33992
rect 16488 33983 16540 33992
rect 16488 33949 16497 33983
rect 16497 33949 16531 33983
rect 16531 33949 16540 33983
rect 16488 33940 16540 33949
rect 18420 33983 18472 33992
rect 18420 33949 18429 33983
rect 18429 33949 18463 33983
rect 18463 33949 18472 33983
rect 18420 33940 18472 33949
rect 19340 33983 19392 33992
rect 19340 33949 19349 33983
rect 19349 33949 19383 33983
rect 19383 33949 19392 33983
rect 19340 33940 19392 33949
rect 20168 33940 20220 33992
rect 29276 34008 29328 34060
rect 21364 33983 21416 33992
rect 21364 33949 21373 33983
rect 21373 33949 21407 33983
rect 21407 33949 21416 33983
rect 21364 33940 21416 33949
rect 22192 33940 22244 33992
rect 22376 33983 22428 33992
rect 22376 33949 22410 33983
rect 22410 33949 22428 33983
rect 22376 33940 22428 33949
rect 24952 33940 25004 33992
rect 25780 33940 25832 33992
rect 28724 33983 28776 33992
rect 28724 33949 28733 33983
rect 28733 33949 28767 33983
rect 28767 33949 28776 33983
rect 28724 33940 28776 33949
rect 29460 33940 29512 33992
rect 29736 33983 29788 33992
rect 29736 33949 29745 33983
rect 29745 33949 29779 33983
rect 29779 33949 29788 33983
rect 29736 33940 29788 33949
rect 30104 33940 30156 33992
rect 30196 33983 30248 33992
rect 30196 33949 30205 33983
rect 30205 33949 30239 33983
rect 30239 33949 30248 33983
rect 30840 33983 30892 33992
rect 30196 33940 30248 33949
rect 30840 33949 30849 33983
rect 30849 33949 30883 33983
rect 30883 33949 30892 33983
rect 30840 33940 30892 33949
rect 31116 33983 31168 33992
rect 31116 33949 31125 33983
rect 31125 33949 31159 33983
rect 31159 33949 31168 33983
rect 31116 33940 31168 33949
rect 11704 33915 11756 33924
rect 11704 33881 11713 33915
rect 11713 33881 11747 33915
rect 11747 33881 11756 33915
rect 11704 33872 11756 33881
rect 13360 33872 13412 33924
rect 16580 33872 16632 33924
rect 22008 33872 22060 33924
rect 3332 33804 3384 33856
rect 8300 33847 8352 33856
rect 8300 33813 8309 33847
rect 8309 33813 8343 33847
rect 8343 33813 8352 33847
rect 8300 33804 8352 33813
rect 8944 33804 8996 33856
rect 12164 33804 12216 33856
rect 13452 33804 13504 33856
rect 14280 33847 14332 33856
rect 14280 33813 14289 33847
rect 14289 33813 14323 33847
rect 14323 33813 14332 33847
rect 14280 33804 14332 33813
rect 15752 33804 15804 33856
rect 18788 33804 18840 33856
rect 22100 33804 22152 33856
rect 22376 33804 22428 33856
rect 24676 33915 24728 33924
rect 24676 33881 24710 33915
rect 24710 33881 24728 33915
rect 24676 33872 24728 33881
rect 27804 33804 27856 33856
rect 28724 33804 28776 33856
rect 30196 33804 30248 33856
rect 7288 33702 7340 33754
rect 17592 33702 17644 33754
rect 27896 33702 27948 33754
rect 5080 33643 5132 33652
rect 5080 33609 5089 33643
rect 5089 33609 5123 33643
rect 5123 33609 5132 33643
rect 5080 33600 5132 33609
rect 7564 33643 7616 33652
rect 7564 33609 7573 33643
rect 7573 33609 7607 33643
rect 7607 33609 7616 33643
rect 7564 33600 7616 33609
rect 10232 33600 10284 33652
rect 11704 33600 11756 33652
rect 2688 33532 2740 33584
rect 1400 33507 1452 33516
rect 1400 33473 1409 33507
rect 1409 33473 1443 33507
rect 1443 33473 1452 33507
rect 1400 33464 1452 33473
rect 1676 33507 1728 33516
rect 1676 33473 1710 33507
rect 1710 33473 1728 33507
rect 4436 33532 4488 33584
rect 5448 33532 5500 33584
rect 1676 33464 1728 33473
rect 3332 33464 3384 33516
rect 5356 33464 5408 33516
rect 4712 33328 4764 33380
rect 5724 33507 5776 33516
rect 5724 33473 5733 33507
rect 5733 33473 5767 33507
rect 5767 33473 5776 33507
rect 5724 33464 5776 33473
rect 6736 33464 6788 33516
rect 7472 33464 7524 33516
rect 7748 33507 7800 33516
rect 7748 33473 7757 33507
rect 7757 33473 7791 33507
rect 7791 33473 7800 33507
rect 7748 33464 7800 33473
rect 8024 33507 8076 33516
rect 8024 33473 8033 33507
rect 8033 33473 8067 33507
rect 8067 33473 8076 33507
rect 8024 33464 8076 33473
rect 9128 33464 9180 33516
rect 9312 33464 9364 33516
rect 10416 33532 10468 33584
rect 10692 33464 10744 33516
rect 11704 33507 11756 33516
rect 7840 33396 7892 33448
rect 8116 33396 8168 33448
rect 9956 33396 10008 33448
rect 11704 33473 11713 33507
rect 11713 33473 11747 33507
rect 11747 33473 11756 33507
rect 11704 33464 11756 33473
rect 11980 33464 12032 33516
rect 14280 33532 14332 33584
rect 15200 33600 15252 33652
rect 15752 33643 15804 33652
rect 15752 33609 15761 33643
rect 15761 33609 15795 33643
rect 15795 33609 15804 33643
rect 15752 33600 15804 33609
rect 18420 33600 18472 33652
rect 18512 33600 18564 33652
rect 13728 33464 13780 33516
rect 16672 33464 16724 33516
rect 16856 33507 16908 33516
rect 16856 33473 16865 33507
rect 16865 33473 16899 33507
rect 16899 33473 16908 33507
rect 16856 33464 16908 33473
rect 17868 33464 17920 33516
rect 19340 33532 19392 33584
rect 20168 33600 20220 33652
rect 21916 33643 21968 33652
rect 21916 33609 21925 33643
rect 21925 33609 21959 33643
rect 21959 33609 21968 33643
rect 21916 33600 21968 33609
rect 24676 33600 24728 33652
rect 25688 33643 25740 33652
rect 25688 33609 25713 33643
rect 25713 33609 25740 33643
rect 25688 33600 25740 33609
rect 29092 33600 29144 33652
rect 30012 33600 30064 33652
rect 30840 33600 30892 33652
rect 18788 33464 18840 33516
rect 21548 33532 21600 33584
rect 22928 33532 22980 33584
rect 25504 33575 25556 33584
rect 13176 33439 13228 33448
rect 13176 33405 13185 33439
rect 13185 33405 13219 33439
rect 13219 33405 13228 33439
rect 13176 33396 13228 33405
rect 15936 33439 15988 33448
rect 15936 33405 15945 33439
rect 15945 33405 15979 33439
rect 15979 33405 15988 33439
rect 15936 33396 15988 33405
rect 20628 33396 20680 33448
rect 21180 33464 21232 33516
rect 22836 33507 22888 33516
rect 22836 33473 22845 33507
rect 22845 33473 22879 33507
rect 22879 33473 22888 33507
rect 22836 33464 22888 33473
rect 23848 33464 23900 33516
rect 22100 33396 22152 33448
rect 22560 33396 22612 33448
rect 24768 33507 24820 33516
rect 24768 33473 24777 33507
rect 24777 33473 24811 33507
rect 24811 33473 24820 33507
rect 24768 33464 24820 33473
rect 25504 33541 25513 33575
rect 25513 33541 25547 33575
rect 25547 33541 25556 33575
rect 25504 33532 25556 33541
rect 27160 33507 27212 33516
rect 27160 33473 27169 33507
rect 27169 33473 27203 33507
rect 27203 33473 27212 33507
rect 27160 33464 27212 33473
rect 27620 33507 27672 33516
rect 6552 33328 6604 33380
rect 10232 33328 10284 33380
rect 21364 33328 21416 33380
rect 21548 33328 21600 33380
rect 23480 33328 23532 33380
rect 24124 33328 24176 33380
rect 27068 33396 27120 33448
rect 27620 33473 27629 33507
rect 27629 33473 27663 33507
rect 27663 33473 27672 33507
rect 27620 33464 27672 33473
rect 29000 33532 29052 33584
rect 29276 33532 29328 33584
rect 30104 33532 30156 33584
rect 28540 33507 28592 33516
rect 28540 33473 28574 33507
rect 28574 33473 28592 33507
rect 28540 33464 28592 33473
rect 29736 33464 29788 33516
rect 29460 33396 29512 33448
rect 31300 33396 31352 33448
rect 2872 33260 2924 33312
rect 4620 33303 4672 33312
rect 4620 33269 4629 33303
rect 4629 33269 4663 33303
rect 4663 33269 4672 33303
rect 4620 33260 4672 33269
rect 7748 33260 7800 33312
rect 10140 33303 10192 33312
rect 10140 33269 10149 33303
rect 10149 33269 10183 33303
rect 10183 33269 10192 33303
rect 10140 33260 10192 33269
rect 10784 33303 10836 33312
rect 10784 33269 10793 33303
rect 10793 33269 10827 33303
rect 10827 33269 10836 33303
rect 10784 33260 10836 33269
rect 12532 33303 12584 33312
rect 12532 33269 12541 33303
rect 12541 33269 12575 33303
rect 12575 33269 12584 33303
rect 12532 33260 12584 33269
rect 14556 33303 14608 33312
rect 14556 33269 14565 33303
rect 14565 33269 14599 33303
rect 14599 33269 14608 33303
rect 14556 33260 14608 33269
rect 18236 33303 18288 33312
rect 18236 33269 18245 33303
rect 18245 33269 18279 33303
rect 18279 33269 18288 33303
rect 18236 33260 18288 33269
rect 20168 33260 20220 33312
rect 20720 33260 20772 33312
rect 22008 33303 22060 33312
rect 22008 33269 22017 33303
rect 22017 33269 22051 33303
rect 22051 33269 22060 33303
rect 22008 33260 22060 33269
rect 22284 33260 22336 33312
rect 23296 33260 23348 33312
rect 23664 33303 23716 33312
rect 23664 33269 23673 33303
rect 23673 33269 23707 33303
rect 23707 33269 23716 33303
rect 23664 33260 23716 33269
rect 23848 33303 23900 33312
rect 23848 33269 23857 33303
rect 23857 33269 23891 33303
rect 23891 33269 23900 33303
rect 23848 33260 23900 33269
rect 25136 33260 25188 33312
rect 26148 33260 26200 33312
rect 28172 33260 28224 33312
rect 2136 33158 2188 33210
rect 12440 33158 12492 33210
rect 22744 33158 22796 33210
rect 1676 33099 1728 33108
rect 1676 33065 1685 33099
rect 1685 33065 1719 33099
rect 1719 33065 1728 33099
rect 1676 33056 1728 33065
rect 2872 33056 2924 33108
rect 3240 33056 3292 33108
rect 2780 32988 2832 33040
rect 2504 32852 2556 32904
rect 3424 32920 3476 32972
rect 4160 32988 4212 33040
rect 5356 32988 5408 33040
rect 7564 32988 7616 33040
rect 4620 32920 4672 32972
rect 5448 32920 5500 32972
rect 11612 33056 11664 33108
rect 8300 32988 8352 33040
rect 10416 32963 10468 32972
rect 3056 32895 3108 32904
rect 3056 32861 3065 32895
rect 3065 32861 3099 32895
rect 3099 32861 3108 32895
rect 3056 32852 3108 32861
rect 3976 32895 4028 32904
rect 3976 32861 3985 32895
rect 3985 32861 4019 32895
rect 4019 32861 4028 32895
rect 3976 32852 4028 32861
rect 4528 32852 4580 32904
rect 4712 32895 4764 32904
rect 4712 32861 4721 32895
rect 4721 32861 4755 32895
rect 4755 32861 4764 32895
rect 4712 32852 4764 32861
rect 5908 32895 5960 32904
rect 5908 32861 5917 32895
rect 5917 32861 5951 32895
rect 5951 32861 5960 32895
rect 5908 32852 5960 32861
rect 6092 32895 6144 32904
rect 6092 32861 6101 32895
rect 6101 32861 6135 32895
rect 6135 32861 6144 32895
rect 6092 32852 6144 32861
rect 6828 32852 6880 32904
rect 7012 32895 7064 32904
rect 7012 32861 7021 32895
rect 7021 32861 7055 32895
rect 7055 32861 7064 32895
rect 7012 32852 7064 32861
rect 7104 32895 7156 32904
rect 7104 32861 7113 32895
rect 7113 32861 7147 32895
rect 7147 32861 7156 32895
rect 7104 32852 7156 32861
rect 8116 32852 8168 32904
rect 3976 32716 4028 32768
rect 5816 32784 5868 32836
rect 6368 32784 6420 32836
rect 5724 32759 5776 32768
rect 5724 32725 5733 32759
rect 5733 32725 5767 32759
rect 5767 32725 5776 32759
rect 5724 32716 5776 32725
rect 7656 32716 7708 32768
rect 8024 32716 8076 32768
rect 10416 32929 10425 32963
rect 10425 32929 10459 32963
rect 10459 32929 10468 32963
rect 10416 32920 10468 32929
rect 11888 32920 11940 32972
rect 14924 33056 14976 33108
rect 16028 33056 16080 33108
rect 22836 33099 22888 33108
rect 17040 32988 17092 33040
rect 21732 32988 21784 33040
rect 22836 33065 22845 33099
rect 22845 33065 22879 33099
rect 22879 33065 22888 33099
rect 22836 33056 22888 33065
rect 25412 33056 25464 33108
rect 25780 33056 25832 33108
rect 28632 33056 28684 33108
rect 24400 32988 24452 33040
rect 13176 32920 13228 32972
rect 10232 32852 10284 32904
rect 12624 32852 12676 32904
rect 13084 32852 13136 32904
rect 8944 32827 8996 32836
rect 8944 32793 8953 32827
rect 8953 32793 8987 32827
rect 8987 32793 8996 32827
rect 8944 32784 8996 32793
rect 9864 32784 9916 32836
rect 11704 32784 11756 32836
rect 11888 32784 11940 32836
rect 14188 32852 14240 32904
rect 14556 32895 14608 32904
rect 14556 32861 14565 32895
rect 14565 32861 14599 32895
rect 14599 32861 14608 32895
rect 14556 32852 14608 32861
rect 14924 32852 14976 32904
rect 15384 32895 15436 32904
rect 15384 32861 15418 32895
rect 15418 32861 15436 32895
rect 15384 32852 15436 32861
rect 15752 32852 15804 32904
rect 16212 32852 16264 32904
rect 18788 32920 18840 32972
rect 20352 32920 20404 32972
rect 20536 32920 20588 32972
rect 21824 32920 21876 32972
rect 23204 32920 23256 32972
rect 23572 32963 23624 32972
rect 23572 32929 23581 32963
rect 23581 32929 23615 32963
rect 23615 32929 23624 32963
rect 23572 32920 23624 32929
rect 23664 32963 23716 32972
rect 23664 32929 23673 32963
rect 23673 32929 23707 32963
rect 23707 32929 23716 32963
rect 27620 32988 27672 33040
rect 23664 32920 23716 32929
rect 9312 32759 9364 32768
rect 9312 32725 9321 32759
rect 9321 32725 9355 32759
rect 9355 32725 9364 32759
rect 9312 32716 9364 32725
rect 12256 32759 12308 32768
rect 12256 32725 12265 32759
rect 12265 32725 12299 32759
rect 12299 32725 12308 32759
rect 12256 32716 12308 32725
rect 13176 32716 13228 32768
rect 14096 32759 14148 32768
rect 14096 32725 14105 32759
rect 14105 32725 14139 32759
rect 14139 32725 14148 32759
rect 14096 32716 14148 32725
rect 16120 32784 16172 32836
rect 18236 32784 18288 32836
rect 19616 32852 19668 32904
rect 21732 32852 21784 32904
rect 20444 32784 20496 32836
rect 22928 32852 22980 32904
rect 21916 32784 21968 32836
rect 23848 32852 23900 32904
rect 24952 32895 25004 32904
rect 24952 32861 24961 32895
rect 24961 32861 24995 32895
rect 24995 32861 25004 32895
rect 24952 32852 25004 32861
rect 26056 32895 26108 32904
rect 23940 32784 23992 32836
rect 26056 32861 26065 32895
rect 26065 32861 26099 32895
rect 26099 32861 26108 32895
rect 26056 32852 26108 32861
rect 16396 32716 16448 32768
rect 17224 32716 17276 32768
rect 19708 32716 19760 32768
rect 21180 32716 21232 32768
rect 22836 32716 22888 32768
rect 23388 32716 23440 32768
rect 24676 32716 24728 32768
rect 26700 32852 26752 32904
rect 27160 32920 27212 32972
rect 27528 32920 27580 32972
rect 29092 33056 29144 33108
rect 31300 33099 31352 33108
rect 31300 33065 31309 33099
rect 31309 33065 31343 33099
rect 31343 33065 31352 33099
rect 31300 33056 31352 33065
rect 28908 33031 28960 33040
rect 28908 32997 28917 33031
rect 28917 32997 28951 33031
rect 28951 32997 28960 33031
rect 28908 32988 28960 32997
rect 29276 32920 29328 32972
rect 27068 32895 27120 32904
rect 27068 32861 27077 32895
rect 27077 32861 27111 32895
rect 27111 32861 27120 32895
rect 27068 32852 27120 32861
rect 27804 32852 27856 32904
rect 28264 32852 28316 32904
rect 28632 32852 28684 32904
rect 30196 32895 30248 32904
rect 26332 32784 26384 32836
rect 28080 32784 28132 32836
rect 29552 32784 29604 32836
rect 30196 32861 30230 32895
rect 30230 32861 30248 32895
rect 30196 32852 30248 32861
rect 30472 32784 30524 32836
rect 30932 32784 30984 32836
rect 27528 32716 27580 32768
rect 28908 32716 28960 32768
rect 29644 32716 29696 32768
rect 31116 32716 31168 32768
rect 7288 32614 7340 32666
rect 17592 32614 17644 32666
rect 27896 32614 27948 32666
rect 5632 32512 5684 32564
rect 5908 32512 5960 32564
rect 9312 32512 9364 32564
rect 12256 32512 12308 32564
rect 3056 32444 3108 32496
rect 1400 32419 1452 32428
rect 1400 32385 1409 32419
rect 1409 32385 1443 32419
rect 1443 32385 1452 32419
rect 1400 32376 1452 32385
rect 2412 32376 2464 32428
rect 3424 32419 3476 32428
rect 3424 32385 3433 32419
rect 3433 32385 3467 32419
rect 3467 32385 3476 32419
rect 3424 32376 3476 32385
rect 4252 32444 4304 32496
rect 4528 32444 4580 32496
rect 5724 32444 5776 32496
rect 4436 32419 4488 32428
rect 2504 32240 2556 32292
rect 4436 32385 4445 32419
rect 4445 32385 4479 32419
rect 4479 32385 4488 32419
rect 4436 32376 4488 32385
rect 4988 32376 5040 32428
rect 7840 32487 7892 32496
rect 7840 32453 7849 32487
rect 7849 32453 7883 32487
rect 7883 32453 7892 32487
rect 7840 32444 7892 32453
rect 8208 32444 8260 32496
rect 5448 32308 5500 32360
rect 6644 32376 6696 32428
rect 2688 32172 2740 32224
rect 6552 32240 6604 32292
rect 5632 32172 5684 32224
rect 6644 32172 6696 32224
rect 9220 32376 9272 32428
rect 11520 32444 11572 32496
rect 11612 32444 11664 32496
rect 13360 32512 13412 32564
rect 14464 32555 14516 32564
rect 12716 32444 12768 32496
rect 14096 32444 14148 32496
rect 14464 32521 14473 32555
rect 14473 32521 14507 32555
rect 14507 32521 14516 32555
rect 14464 32512 14516 32521
rect 15384 32512 15436 32564
rect 16120 32555 16172 32564
rect 16120 32521 16129 32555
rect 16129 32521 16163 32555
rect 16163 32521 16172 32555
rect 16120 32512 16172 32521
rect 16672 32555 16724 32564
rect 16672 32521 16681 32555
rect 16681 32521 16715 32555
rect 16715 32521 16724 32555
rect 16672 32512 16724 32521
rect 17868 32555 17920 32564
rect 17868 32521 17877 32555
rect 17877 32521 17911 32555
rect 17911 32521 17920 32555
rect 17868 32512 17920 32521
rect 19340 32512 19392 32564
rect 9404 32308 9456 32360
rect 12256 32376 12308 32428
rect 15200 32444 15252 32496
rect 15660 32444 15712 32496
rect 12624 32351 12676 32360
rect 12624 32317 12633 32351
rect 12633 32317 12667 32351
rect 12667 32317 12676 32351
rect 12624 32308 12676 32317
rect 10508 32240 10560 32292
rect 8944 32215 8996 32224
rect 8944 32181 8953 32215
rect 8953 32181 8987 32215
rect 8987 32181 8996 32215
rect 8944 32172 8996 32181
rect 12072 32215 12124 32224
rect 12072 32181 12081 32215
rect 12081 32181 12115 32215
rect 12115 32181 12124 32215
rect 12072 32172 12124 32181
rect 14372 32308 14424 32360
rect 15016 32376 15068 32428
rect 15568 32376 15620 32428
rect 17040 32419 17092 32428
rect 17040 32385 17049 32419
rect 17049 32385 17083 32419
rect 17083 32385 17092 32419
rect 17040 32376 17092 32385
rect 15292 32308 15344 32360
rect 15476 32308 15528 32360
rect 16948 32308 17000 32360
rect 17132 32351 17184 32360
rect 17132 32317 17141 32351
rect 17141 32317 17175 32351
rect 17175 32317 17184 32351
rect 17132 32308 17184 32317
rect 17684 32376 17736 32428
rect 18144 32376 18196 32428
rect 19524 32444 19576 32496
rect 19984 32512 20036 32564
rect 27712 32512 27764 32564
rect 28080 32512 28132 32564
rect 28356 32512 28408 32564
rect 28448 32512 28500 32564
rect 18972 32376 19024 32428
rect 19616 32419 19668 32428
rect 19616 32385 19625 32419
rect 19625 32385 19659 32419
rect 19659 32385 19668 32419
rect 19616 32376 19668 32385
rect 20352 32419 20404 32428
rect 20352 32385 20361 32419
rect 20361 32385 20395 32419
rect 20395 32385 20404 32419
rect 20352 32376 20404 32385
rect 21180 32487 21232 32496
rect 21180 32453 21189 32487
rect 21189 32453 21223 32487
rect 21223 32453 21232 32487
rect 21180 32444 21232 32453
rect 14832 32240 14884 32292
rect 16304 32240 16356 32292
rect 20168 32308 20220 32360
rect 20628 32308 20680 32360
rect 17776 32240 17828 32292
rect 21180 32308 21232 32360
rect 21364 32308 21416 32360
rect 21916 32308 21968 32360
rect 22100 32419 22152 32428
rect 22100 32385 22109 32419
rect 22109 32385 22143 32419
rect 22143 32385 22152 32419
rect 22560 32419 22612 32428
rect 22100 32376 22152 32385
rect 22560 32385 22569 32419
rect 22569 32385 22603 32419
rect 22603 32385 22612 32419
rect 22560 32376 22612 32385
rect 23296 32444 23348 32496
rect 23572 32376 23624 32428
rect 26516 32444 26568 32496
rect 24676 32419 24728 32428
rect 24676 32385 24710 32419
rect 24710 32385 24728 32419
rect 24676 32376 24728 32385
rect 26792 32376 26844 32428
rect 27528 32376 27580 32428
rect 28264 32376 28316 32428
rect 29460 32419 29512 32428
rect 29460 32385 29469 32419
rect 29469 32385 29503 32419
rect 29503 32385 29512 32419
rect 29460 32376 29512 32385
rect 12900 32172 12952 32224
rect 14464 32172 14516 32224
rect 17960 32172 18012 32224
rect 19432 32172 19484 32224
rect 19708 32172 19760 32224
rect 20720 32172 20772 32224
rect 20996 32215 21048 32224
rect 20996 32181 21005 32215
rect 21005 32181 21039 32215
rect 21039 32181 21048 32215
rect 20996 32172 21048 32181
rect 22468 32240 22520 32292
rect 23940 32283 23992 32292
rect 23940 32249 23949 32283
rect 23949 32249 23983 32283
rect 23983 32249 23992 32283
rect 23940 32240 23992 32249
rect 29644 32351 29696 32360
rect 29644 32317 29653 32351
rect 29653 32317 29687 32351
rect 29687 32317 29696 32351
rect 30380 32351 30432 32360
rect 29644 32308 29696 32317
rect 27528 32240 27580 32292
rect 27620 32240 27672 32292
rect 21916 32172 21968 32224
rect 23480 32172 23532 32224
rect 25872 32172 25924 32224
rect 26240 32215 26292 32224
rect 26240 32181 26249 32215
rect 26249 32181 26283 32215
rect 26283 32181 26292 32215
rect 26240 32172 26292 32181
rect 29828 32240 29880 32292
rect 29092 32172 29144 32224
rect 30380 32317 30389 32351
rect 30389 32317 30423 32351
rect 30423 32317 30432 32351
rect 30380 32308 30432 32317
rect 30472 32351 30524 32360
rect 30472 32317 30506 32351
rect 30506 32317 30524 32351
rect 30472 32308 30524 32317
rect 30656 32351 30708 32360
rect 30656 32317 30665 32351
rect 30665 32317 30699 32351
rect 30699 32317 30708 32351
rect 30656 32308 30708 32317
rect 30380 32172 30432 32224
rect 30656 32172 30708 32224
rect 2136 32070 2188 32122
rect 12440 32070 12492 32122
rect 22744 32070 22796 32122
rect 2412 32011 2464 32020
rect 2412 31977 2421 32011
rect 2421 31977 2455 32011
rect 2455 31977 2464 32011
rect 2412 31968 2464 31977
rect 2964 31968 3016 32020
rect 8944 31968 8996 32020
rect 11704 31968 11756 32020
rect 11980 31968 12032 32020
rect 20352 31968 20404 32020
rect 21180 31968 21232 32020
rect 2780 31943 2832 31952
rect 2780 31909 2789 31943
rect 2789 31909 2823 31943
rect 2823 31909 2832 31943
rect 2780 31900 2832 31909
rect 2044 31764 2096 31816
rect 2688 31764 2740 31816
rect 2872 31807 2924 31816
rect 2872 31773 2881 31807
rect 2881 31773 2915 31807
rect 2915 31773 2924 31807
rect 2872 31764 2924 31773
rect 4068 31900 4120 31952
rect 6828 31900 6880 31952
rect 4988 31875 5040 31884
rect 4988 31841 4997 31875
rect 4997 31841 5031 31875
rect 5031 31841 5040 31875
rect 4988 31832 5040 31841
rect 4160 31764 4212 31816
rect 4252 31807 4304 31816
rect 4252 31773 4261 31807
rect 4261 31773 4295 31807
rect 4295 31773 4304 31807
rect 4252 31764 4304 31773
rect 4620 31764 4672 31816
rect 6092 31832 6144 31884
rect 6368 31832 6420 31884
rect 6460 31807 6512 31816
rect 6460 31773 6469 31807
rect 6469 31773 6503 31807
rect 6503 31773 6512 31807
rect 6460 31764 6512 31773
rect 6552 31807 6604 31816
rect 6552 31773 6562 31807
rect 6562 31773 6596 31807
rect 6596 31773 6604 31807
rect 6552 31764 6604 31773
rect 6828 31807 6880 31816
rect 6828 31773 6837 31807
rect 6837 31773 6871 31807
rect 6871 31773 6880 31807
rect 6828 31764 6880 31773
rect 7472 31696 7524 31748
rect 7656 31832 7708 31884
rect 8024 31875 8076 31884
rect 8024 31841 8033 31875
rect 8033 31841 8067 31875
rect 8067 31841 8076 31875
rect 8024 31832 8076 31841
rect 7748 31807 7800 31816
rect 7748 31773 7757 31807
rect 7757 31773 7791 31807
rect 7791 31773 7800 31807
rect 7748 31764 7800 31773
rect 7932 31807 7984 31816
rect 7932 31773 7941 31807
rect 7941 31773 7975 31807
rect 7975 31773 7984 31807
rect 7932 31764 7984 31773
rect 8300 31764 8352 31816
rect 8024 31696 8076 31748
rect 9312 31739 9364 31748
rect 9312 31705 9321 31739
rect 9321 31705 9355 31739
rect 9355 31705 9364 31739
rect 9312 31696 9364 31705
rect 9404 31696 9456 31748
rect 10508 31807 10560 31816
rect 10508 31773 10517 31807
rect 10517 31773 10551 31807
rect 10551 31773 10560 31807
rect 10508 31764 10560 31773
rect 12716 31900 12768 31952
rect 12808 31900 12860 31952
rect 14188 31943 14240 31952
rect 12164 31875 12216 31884
rect 12164 31841 12173 31875
rect 12173 31841 12207 31875
rect 12207 31841 12216 31875
rect 12164 31832 12216 31841
rect 12072 31764 12124 31816
rect 11888 31696 11940 31748
rect 12716 31764 12768 31816
rect 14188 31909 14197 31943
rect 14197 31909 14231 31943
rect 14231 31909 14240 31943
rect 14188 31900 14240 31909
rect 13360 31807 13412 31816
rect 13360 31773 13369 31807
rect 13369 31773 13403 31807
rect 13403 31773 13412 31807
rect 13360 31764 13412 31773
rect 14372 31807 14424 31816
rect 14372 31773 14381 31807
rect 14381 31773 14415 31807
rect 14415 31773 14424 31807
rect 14372 31764 14424 31773
rect 15200 31900 15252 31952
rect 17224 31943 17276 31952
rect 17224 31909 17233 31943
rect 17233 31909 17267 31943
rect 17267 31909 17276 31943
rect 17224 31900 17276 31909
rect 17868 31900 17920 31952
rect 21548 31900 21600 31952
rect 22376 31900 22428 31952
rect 22928 31968 22980 32020
rect 24952 31968 25004 32020
rect 26240 31968 26292 32020
rect 15108 31832 15160 31884
rect 16028 31832 16080 31884
rect 16948 31832 17000 31884
rect 18144 31832 18196 31884
rect 14832 31807 14884 31816
rect 14832 31773 14841 31807
rect 14841 31773 14875 31807
rect 14875 31773 14884 31807
rect 14832 31764 14884 31773
rect 15660 31807 15712 31816
rect 15660 31773 15669 31807
rect 15669 31773 15703 31807
rect 15703 31773 15712 31807
rect 15660 31764 15712 31773
rect 16580 31807 16632 31816
rect 7564 31628 7616 31680
rect 9036 31628 9088 31680
rect 11428 31671 11480 31680
rect 11428 31637 11437 31671
rect 11437 31637 11471 31671
rect 11471 31637 11480 31671
rect 16120 31696 16172 31748
rect 15476 31671 15528 31680
rect 11428 31628 11480 31637
rect 15476 31637 15485 31671
rect 15485 31637 15519 31671
rect 15519 31637 15528 31671
rect 15476 31628 15528 31637
rect 16580 31773 16589 31807
rect 16589 31773 16623 31807
rect 16623 31773 16632 31807
rect 16580 31764 16632 31773
rect 18328 31764 18380 31816
rect 19248 31807 19300 31816
rect 17040 31628 17092 31680
rect 17776 31696 17828 31748
rect 19248 31773 19257 31807
rect 19257 31773 19291 31807
rect 19291 31773 19300 31807
rect 19248 31764 19300 31773
rect 19340 31696 19392 31748
rect 19524 31807 19576 31816
rect 19524 31773 19558 31807
rect 19558 31773 19576 31807
rect 19524 31764 19576 31773
rect 20720 31764 20772 31816
rect 17408 31628 17460 31680
rect 17960 31628 18012 31680
rect 18512 31628 18564 31680
rect 19064 31628 19116 31680
rect 20260 31628 20312 31680
rect 21088 31628 21140 31680
rect 21364 31628 21416 31680
rect 21548 31807 21600 31816
rect 21548 31773 21557 31807
rect 21557 31773 21591 31807
rect 21591 31773 21600 31807
rect 21548 31764 21600 31773
rect 21732 31807 21784 31816
rect 21732 31773 21741 31807
rect 21741 31773 21775 31807
rect 21775 31773 21784 31807
rect 22376 31807 22428 31816
rect 21732 31764 21784 31773
rect 22376 31773 22385 31807
rect 22385 31773 22419 31807
rect 22419 31773 22428 31807
rect 22376 31764 22428 31773
rect 22652 31875 22704 31884
rect 22652 31841 22661 31875
rect 22661 31841 22695 31875
rect 22695 31841 22704 31875
rect 22652 31832 22704 31841
rect 22836 31764 22888 31816
rect 25688 31900 25740 31952
rect 27620 31968 27672 32020
rect 28540 32011 28592 32020
rect 28540 31977 28549 32011
rect 28549 31977 28583 32011
rect 28583 31977 28592 32011
rect 28540 31968 28592 31977
rect 29736 31968 29788 32020
rect 28908 31900 28960 31952
rect 23480 31807 23532 31816
rect 23480 31773 23489 31807
rect 23489 31773 23523 31807
rect 23523 31773 23532 31807
rect 23480 31764 23532 31773
rect 25504 31832 25556 31884
rect 26332 31832 26384 31884
rect 26516 31875 26568 31884
rect 26516 31841 26525 31875
rect 26525 31841 26559 31875
rect 26559 31841 26568 31875
rect 26516 31832 26568 31841
rect 27528 31832 27580 31884
rect 29184 31832 29236 31884
rect 30104 31832 30156 31884
rect 22468 31696 22520 31748
rect 25964 31764 26016 31816
rect 28356 31764 28408 31816
rect 28724 31807 28776 31816
rect 28724 31773 28733 31807
rect 28733 31773 28767 31807
rect 28767 31773 28776 31807
rect 28724 31764 28776 31773
rect 28816 31764 28868 31816
rect 30288 31807 30340 31816
rect 30288 31773 30297 31807
rect 30297 31773 30331 31807
rect 30331 31773 30340 31807
rect 30288 31764 30340 31773
rect 30748 31764 30800 31816
rect 26424 31696 26476 31748
rect 26700 31696 26752 31748
rect 23020 31628 23072 31680
rect 24032 31628 24084 31680
rect 24492 31628 24544 31680
rect 30196 31628 30248 31680
rect 31208 31671 31260 31680
rect 31208 31637 31217 31671
rect 31217 31637 31251 31671
rect 31251 31637 31260 31671
rect 31208 31628 31260 31637
rect 7288 31526 7340 31578
rect 17592 31526 17644 31578
rect 27896 31526 27948 31578
rect 3884 31424 3936 31476
rect 2044 31356 2096 31408
rect 2504 31356 2556 31408
rect 2596 31331 2648 31340
rect 2596 31297 2605 31331
rect 2605 31297 2639 31331
rect 2639 31297 2648 31331
rect 2596 31288 2648 31297
rect 3976 31288 4028 31340
rect 4252 31288 4304 31340
rect 7932 31424 7984 31476
rect 8024 31424 8076 31476
rect 6644 31356 6696 31408
rect 1768 31220 1820 31272
rect 2044 31220 2096 31272
rect 3608 31220 3660 31272
rect 4068 31220 4120 31272
rect 4804 31263 4856 31272
rect 4804 31229 4813 31263
rect 4813 31229 4847 31263
rect 4847 31229 4856 31263
rect 4804 31220 4856 31229
rect 7012 31331 7064 31340
rect 7012 31297 7021 31331
rect 7021 31297 7055 31331
rect 7055 31297 7064 31331
rect 7012 31288 7064 31297
rect 7380 31220 7432 31272
rect 7656 31220 7708 31272
rect 8116 31220 8168 31272
rect 5172 31152 5224 31204
rect 7012 31152 7064 31204
rect 8668 31263 8720 31272
rect 8668 31229 8677 31263
rect 8677 31229 8711 31263
rect 8711 31229 8720 31263
rect 9588 31356 9640 31408
rect 9864 31424 9916 31476
rect 11888 31424 11940 31476
rect 13268 31467 13320 31476
rect 11704 31356 11756 31408
rect 11980 31399 12032 31408
rect 11980 31365 11989 31399
rect 11989 31365 12023 31399
rect 12023 31365 12032 31399
rect 11980 31356 12032 31365
rect 8668 31220 8720 31229
rect 10048 31288 10100 31340
rect 11060 31288 11112 31340
rect 11152 31220 11204 31272
rect 11796 31220 11848 31272
rect 10600 31152 10652 31204
rect 11888 31152 11940 31204
rect 12808 31220 12860 31272
rect 13268 31433 13277 31467
rect 13277 31433 13311 31467
rect 13311 31433 13320 31467
rect 13268 31424 13320 31433
rect 14648 31424 14700 31476
rect 15660 31424 15712 31476
rect 16120 31424 16172 31476
rect 15200 31356 15252 31408
rect 13176 31288 13228 31340
rect 13268 31288 13320 31340
rect 14280 31288 14332 31340
rect 15292 31288 15344 31340
rect 15660 31288 15712 31340
rect 15936 31331 15988 31340
rect 15936 31297 15945 31331
rect 15945 31297 15979 31331
rect 15979 31297 15988 31331
rect 15936 31288 15988 31297
rect 16304 31288 16356 31340
rect 16856 31331 16908 31340
rect 16856 31297 16865 31331
rect 16865 31297 16899 31331
rect 16899 31297 16908 31331
rect 16856 31288 16908 31297
rect 17316 31288 17368 31340
rect 18972 31467 19024 31476
rect 18972 31433 18981 31467
rect 18981 31433 19015 31467
rect 19015 31433 19024 31467
rect 18972 31424 19024 31433
rect 19064 31424 19116 31476
rect 19340 31424 19392 31476
rect 21548 31424 21600 31476
rect 21824 31467 21876 31476
rect 21824 31433 21833 31467
rect 21833 31433 21867 31467
rect 21867 31433 21876 31467
rect 21824 31424 21876 31433
rect 22100 31424 22152 31476
rect 23848 31424 23900 31476
rect 28356 31467 28408 31476
rect 28356 31433 28365 31467
rect 28365 31433 28399 31467
rect 28399 31433 28408 31467
rect 28356 31424 28408 31433
rect 31116 31424 31168 31476
rect 31300 31467 31352 31476
rect 31300 31433 31309 31467
rect 31309 31433 31343 31467
rect 31343 31433 31352 31467
rect 31300 31424 31352 31433
rect 17960 31288 18012 31340
rect 18236 31331 18288 31340
rect 18236 31297 18245 31331
rect 18245 31297 18279 31331
rect 18279 31297 18288 31331
rect 18236 31288 18288 31297
rect 19156 31331 19208 31340
rect 19156 31297 19165 31331
rect 19165 31297 19199 31331
rect 19199 31297 19208 31331
rect 19156 31288 19208 31297
rect 20444 31356 20496 31408
rect 21732 31356 21784 31408
rect 19616 31331 19668 31340
rect 19616 31297 19625 31331
rect 19625 31297 19659 31331
rect 19659 31297 19668 31331
rect 19616 31288 19668 31297
rect 20260 31288 20312 31340
rect 20536 31331 20588 31340
rect 20536 31297 20545 31331
rect 20545 31297 20579 31331
rect 20579 31297 20588 31331
rect 20536 31288 20588 31297
rect 20996 31288 21048 31340
rect 22468 31356 22520 31408
rect 14096 31263 14148 31272
rect 1768 31084 1820 31136
rect 3700 31127 3752 31136
rect 3700 31093 3709 31127
rect 3709 31093 3743 31127
rect 3743 31093 3752 31127
rect 3700 31084 3752 31093
rect 4344 31127 4396 31136
rect 4344 31093 4353 31127
rect 4353 31093 4387 31127
rect 4387 31093 4396 31127
rect 4344 31084 4396 31093
rect 5816 31084 5868 31136
rect 8668 31084 8720 31136
rect 8852 31084 8904 31136
rect 10416 31127 10468 31136
rect 10416 31093 10425 31127
rect 10425 31093 10459 31127
rect 10459 31093 10468 31127
rect 10416 31084 10468 31093
rect 10508 31084 10560 31136
rect 10968 31084 11020 31136
rect 12256 31084 12308 31136
rect 12532 31084 12584 31136
rect 13636 31152 13688 31204
rect 14096 31229 14105 31263
rect 14105 31229 14139 31263
rect 14139 31229 14148 31263
rect 14096 31220 14148 31229
rect 19800 31220 19852 31272
rect 23388 31288 23440 31340
rect 23940 31288 23992 31340
rect 25136 31288 25188 31340
rect 25964 31288 26016 31340
rect 26148 31288 26200 31340
rect 27988 31288 28040 31340
rect 28172 31288 28224 31340
rect 28632 31288 28684 31340
rect 24032 31220 24084 31272
rect 25872 31220 25924 31272
rect 13084 31127 13136 31136
rect 13084 31093 13093 31127
rect 13093 31093 13127 31127
rect 13127 31093 13136 31127
rect 13084 31084 13136 31093
rect 14464 31127 14516 31136
rect 14464 31093 14473 31127
rect 14473 31093 14507 31127
rect 14507 31093 14516 31127
rect 14464 31084 14516 31093
rect 16672 31127 16724 31136
rect 16672 31093 16681 31127
rect 16681 31093 16715 31127
rect 16715 31093 16724 31127
rect 16672 31084 16724 31093
rect 17040 31127 17092 31136
rect 17040 31093 17049 31127
rect 17049 31093 17083 31127
rect 17083 31093 17092 31127
rect 17040 31084 17092 31093
rect 25136 31152 25188 31204
rect 25228 31152 25280 31204
rect 26056 31152 26108 31204
rect 26792 31152 26844 31204
rect 22100 31084 22152 31136
rect 22468 31084 22520 31136
rect 23664 31127 23716 31136
rect 23664 31093 23673 31127
rect 23673 31093 23707 31127
rect 23707 31093 23716 31127
rect 23664 31084 23716 31093
rect 25044 31127 25096 31136
rect 25044 31093 25053 31127
rect 25053 31093 25087 31127
rect 25087 31093 25096 31127
rect 25044 31084 25096 31093
rect 26608 31084 26660 31136
rect 30196 31331 30248 31340
rect 30196 31297 30230 31331
rect 30230 31297 30248 31331
rect 30196 31288 30248 31297
rect 29920 31263 29972 31272
rect 29920 31229 29929 31263
rect 29929 31229 29963 31263
rect 29963 31229 29972 31263
rect 29920 31220 29972 31229
rect 30656 31084 30708 31136
rect 2136 30982 2188 31034
rect 12440 30982 12492 31034
rect 22744 30982 22796 31034
rect 4252 30923 4304 30932
rect 4252 30889 4261 30923
rect 4261 30889 4295 30923
rect 4295 30889 4304 30923
rect 4252 30880 4304 30889
rect 6460 30880 6512 30932
rect 8208 30880 8260 30932
rect 9404 30880 9456 30932
rect 2872 30855 2924 30864
rect 2872 30821 2881 30855
rect 2881 30821 2915 30855
rect 2915 30821 2924 30855
rect 2872 30812 2924 30821
rect 7748 30812 7800 30864
rect 10968 30880 11020 30932
rect 11152 30923 11204 30932
rect 11152 30889 11161 30923
rect 11161 30889 11195 30923
rect 11195 30889 11204 30923
rect 11152 30880 11204 30889
rect 11704 30880 11756 30932
rect 7932 30744 7984 30796
rect 1400 30676 1452 30728
rect 1768 30719 1820 30728
rect 1768 30685 1802 30719
rect 1802 30685 1820 30719
rect 1768 30676 1820 30685
rect 3700 30676 3752 30728
rect 4896 30719 4948 30728
rect 4160 30608 4212 30660
rect 4896 30685 4905 30719
rect 4905 30685 4939 30719
rect 4939 30685 4948 30719
rect 4896 30676 4948 30685
rect 5908 30676 5960 30728
rect 7564 30676 7616 30728
rect 7012 30608 7064 30660
rect 8116 30719 8168 30728
rect 8116 30685 8125 30719
rect 8125 30685 8159 30719
rect 8159 30685 8168 30719
rect 8300 30719 8352 30728
rect 8116 30676 8168 30685
rect 8300 30685 8309 30719
rect 8309 30685 8343 30719
rect 8343 30685 8352 30719
rect 8300 30676 8352 30685
rect 8852 30676 8904 30728
rect 9772 30719 9824 30728
rect 9772 30685 9781 30719
rect 9781 30685 9815 30719
rect 9815 30685 9824 30719
rect 9772 30676 9824 30685
rect 9864 30676 9916 30728
rect 10416 30676 10468 30728
rect 12716 30880 12768 30932
rect 14096 30923 14148 30932
rect 14096 30889 14105 30923
rect 14105 30889 14139 30923
rect 14139 30889 14148 30923
rect 14096 30880 14148 30889
rect 15936 30880 15988 30932
rect 17316 30880 17368 30932
rect 17776 30880 17828 30932
rect 22100 30880 22152 30932
rect 23572 30923 23624 30932
rect 14280 30812 14332 30864
rect 15108 30812 15160 30864
rect 19432 30812 19484 30864
rect 19984 30812 20036 30864
rect 21732 30855 21784 30864
rect 21732 30821 21741 30855
rect 21741 30821 21775 30855
rect 21775 30821 21784 30855
rect 21732 30812 21784 30821
rect 23572 30889 23581 30923
rect 23581 30889 23615 30923
rect 23615 30889 23624 30923
rect 23572 30880 23624 30889
rect 25964 30880 26016 30932
rect 30288 30880 30340 30932
rect 12164 30676 12216 30728
rect 13084 30676 13136 30728
rect 8944 30608 8996 30660
rect 12532 30651 12584 30660
rect 12532 30617 12541 30651
rect 12541 30617 12575 30651
rect 12575 30617 12584 30651
rect 12532 30608 12584 30617
rect 12624 30608 12676 30660
rect 14372 30719 14424 30728
rect 14372 30685 14381 30719
rect 14381 30685 14415 30719
rect 14415 30685 14424 30719
rect 14924 30744 14976 30796
rect 19248 30744 19300 30796
rect 14372 30676 14424 30685
rect 15200 30719 15252 30728
rect 15200 30685 15209 30719
rect 15209 30685 15243 30719
rect 15243 30685 15252 30719
rect 15200 30676 15252 30685
rect 15476 30719 15528 30728
rect 15476 30685 15510 30719
rect 15510 30685 15528 30719
rect 15476 30676 15528 30685
rect 18052 30676 18104 30728
rect 19156 30676 19208 30728
rect 22192 30787 22244 30796
rect 22192 30753 22201 30787
rect 22201 30753 22235 30787
rect 22235 30753 22244 30787
rect 22192 30744 22244 30753
rect 26332 30744 26384 30796
rect 16672 30608 16724 30660
rect 19248 30608 19300 30660
rect 20628 30651 20680 30660
rect 20628 30617 20662 30651
rect 20662 30617 20680 30651
rect 25044 30676 25096 30728
rect 25136 30676 25188 30728
rect 26240 30676 26292 30728
rect 26424 30719 26476 30728
rect 26424 30685 26433 30719
rect 26433 30685 26467 30719
rect 26467 30685 26476 30719
rect 26424 30676 26476 30685
rect 20628 30608 20680 30617
rect 22192 30608 22244 30660
rect 6092 30540 6144 30592
rect 6368 30583 6420 30592
rect 6368 30549 6377 30583
rect 6377 30549 6411 30583
rect 6411 30549 6420 30583
rect 6368 30540 6420 30549
rect 6736 30540 6788 30592
rect 7196 30583 7248 30592
rect 7196 30549 7205 30583
rect 7205 30549 7239 30583
rect 7239 30549 7248 30583
rect 7196 30540 7248 30549
rect 7380 30540 7432 30592
rect 12072 30540 12124 30592
rect 13912 30540 13964 30592
rect 16948 30540 17000 30592
rect 17408 30540 17460 30592
rect 18144 30540 18196 30592
rect 21824 30540 21876 30592
rect 25320 30540 25372 30592
rect 27988 30676 28040 30728
rect 28908 30719 28960 30728
rect 28908 30685 28917 30719
rect 28917 30685 28951 30719
rect 28951 30685 28960 30719
rect 28908 30676 28960 30685
rect 29000 30719 29052 30728
rect 29000 30685 29009 30719
rect 29009 30685 29043 30719
rect 29043 30685 29052 30719
rect 30748 30744 30800 30796
rect 29000 30676 29052 30685
rect 30104 30676 30156 30728
rect 31208 30744 31260 30796
rect 31300 30719 31352 30728
rect 31300 30685 31309 30719
rect 31309 30685 31343 30719
rect 31343 30685 31352 30719
rect 31300 30676 31352 30685
rect 30656 30608 30708 30660
rect 30012 30540 30064 30592
rect 7288 30438 7340 30490
rect 17592 30438 17644 30490
rect 27896 30438 27948 30490
rect 2596 30336 2648 30388
rect 2872 30200 2924 30252
rect 3700 30268 3752 30320
rect 4344 30268 4396 30320
rect 6644 30268 6696 30320
rect 8484 30336 8536 30388
rect 8668 30336 8720 30388
rect 9680 30336 9732 30388
rect 12532 30336 12584 30388
rect 12808 30336 12860 30388
rect 12900 30336 12952 30388
rect 14556 30336 14608 30388
rect 15200 30336 15252 30388
rect 16856 30336 16908 30388
rect 3608 30243 3660 30252
rect 3608 30209 3617 30243
rect 3617 30209 3651 30243
rect 3651 30209 3660 30243
rect 3608 30200 3660 30209
rect 6736 30200 6788 30252
rect 8300 30268 8352 30320
rect 12256 30268 12308 30320
rect 14924 30268 14976 30320
rect 7380 30243 7432 30252
rect 7380 30209 7389 30243
rect 7389 30209 7423 30243
rect 7423 30209 7432 30243
rect 7380 30200 7432 30209
rect 8208 30200 8260 30252
rect 8484 30243 8536 30252
rect 8484 30209 8493 30243
rect 8493 30209 8527 30243
rect 8527 30209 8536 30243
rect 9496 30243 9548 30252
rect 8484 30200 8536 30209
rect 9496 30209 9505 30243
rect 9505 30209 9539 30243
rect 9539 30209 9548 30243
rect 9496 30200 9548 30209
rect 9588 30200 9640 30252
rect 12532 30243 12584 30252
rect 12532 30209 12541 30243
rect 12541 30209 12575 30243
rect 12575 30209 12584 30243
rect 12532 30200 12584 30209
rect 4252 30175 4304 30184
rect 4252 30141 4261 30175
rect 4261 30141 4295 30175
rect 4295 30141 4304 30175
rect 4252 30132 4304 30141
rect 7472 30132 7524 30184
rect 9864 30132 9916 30184
rect 10508 30132 10560 30184
rect 11980 30175 12032 30184
rect 11980 30141 11989 30175
rect 11989 30141 12023 30175
rect 12023 30141 12032 30175
rect 11980 30132 12032 30141
rect 12072 30132 12124 30184
rect 12992 30200 13044 30252
rect 4160 30064 4212 30116
rect 9496 30064 9548 30116
rect 15476 30200 15528 30252
rect 16580 30200 16632 30252
rect 17500 30200 17552 30252
rect 18236 30336 18288 30388
rect 19156 30336 19208 30388
rect 19524 30336 19576 30388
rect 20444 30336 20496 30388
rect 20628 30379 20680 30388
rect 20628 30345 20637 30379
rect 20637 30345 20671 30379
rect 20671 30345 20680 30379
rect 20628 30336 20680 30345
rect 22192 30336 22244 30388
rect 17960 30243 18012 30252
rect 17960 30209 17969 30243
rect 17969 30209 18003 30243
rect 18003 30209 18012 30243
rect 17960 30200 18012 30209
rect 18144 30243 18196 30252
rect 18144 30209 18153 30243
rect 18153 30209 18187 30243
rect 18187 30209 18196 30243
rect 18144 30200 18196 30209
rect 18512 30200 18564 30252
rect 19248 30268 19300 30320
rect 19340 30268 19392 30320
rect 26424 30336 26476 30388
rect 16120 30132 16172 30184
rect 14372 30064 14424 30116
rect 15016 30064 15068 30116
rect 18604 30175 18656 30184
rect 18604 30141 18613 30175
rect 18613 30141 18647 30175
rect 18647 30141 18656 30175
rect 18604 30132 18656 30141
rect 20812 30243 20864 30252
rect 20812 30209 20821 30243
rect 20821 30209 20855 30243
rect 20855 30209 20864 30243
rect 20812 30200 20864 30209
rect 22100 30200 22152 30252
rect 22468 30243 22520 30252
rect 22468 30209 22477 30243
rect 22477 30209 22511 30243
rect 22511 30209 22520 30243
rect 22468 30200 22520 30209
rect 23664 30243 23716 30252
rect 20996 30132 21048 30184
rect 22836 30132 22888 30184
rect 19800 30107 19852 30116
rect 19800 30073 19809 30107
rect 19809 30073 19843 30107
rect 19843 30073 19852 30107
rect 19800 30064 19852 30073
rect 20076 30064 20128 30116
rect 2780 29996 2832 30048
rect 4896 29996 4948 30048
rect 8392 29996 8444 30048
rect 8760 30039 8812 30048
rect 8760 30005 8769 30039
rect 8769 30005 8803 30039
rect 8803 30005 8812 30039
rect 8760 29996 8812 30005
rect 11704 29996 11756 30048
rect 16304 29996 16356 30048
rect 18696 29996 18748 30048
rect 20628 29996 20680 30048
rect 22100 30064 22152 30116
rect 23664 30209 23673 30243
rect 23673 30209 23707 30243
rect 23707 30209 23716 30243
rect 23664 30200 23716 30209
rect 26332 30200 26384 30252
rect 26424 30243 26476 30252
rect 26424 30209 26433 30243
rect 26433 30209 26467 30243
rect 26467 30209 26476 30243
rect 27712 30268 27764 30320
rect 28264 30311 28316 30320
rect 28264 30277 28273 30311
rect 28273 30277 28307 30311
rect 28307 30277 28316 30311
rect 28264 30268 28316 30277
rect 26424 30200 26476 30209
rect 30656 30243 30708 30252
rect 30656 30209 30665 30243
rect 30665 30209 30699 30243
rect 30699 30209 30708 30243
rect 30656 30200 30708 30209
rect 30748 30200 30800 30252
rect 31116 30243 31168 30252
rect 31116 30209 31125 30243
rect 31125 30209 31159 30243
rect 31159 30209 31168 30243
rect 31116 30200 31168 30209
rect 25320 30175 25372 30184
rect 23664 30064 23716 30116
rect 25320 30141 25329 30175
rect 25329 30141 25363 30175
rect 25363 30141 25372 30175
rect 25320 30132 25372 30141
rect 27344 30132 27396 30184
rect 26608 30064 26660 30116
rect 25228 30039 25280 30048
rect 25228 30005 25237 30039
rect 25237 30005 25271 30039
rect 25271 30005 25280 30039
rect 25228 29996 25280 30005
rect 25780 29996 25832 30048
rect 29828 30132 29880 30184
rect 28724 30064 28776 30116
rect 27528 29996 27580 30048
rect 29920 29996 29972 30048
rect 2136 29894 2188 29946
rect 12440 29894 12492 29946
rect 22744 29894 22796 29946
rect 3608 29792 3660 29844
rect 6552 29792 6604 29844
rect 7104 29792 7156 29844
rect 7196 29792 7248 29844
rect 12900 29792 12952 29844
rect 13084 29792 13136 29844
rect 13452 29792 13504 29844
rect 16580 29792 16632 29844
rect 1400 29631 1452 29640
rect 1400 29597 1409 29631
rect 1409 29597 1443 29631
rect 1443 29597 1452 29631
rect 4252 29724 4304 29776
rect 3148 29656 3200 29708
rect 6000 29724 6052 29776
rect 6368 29724 6420 29776
rect 8208 29724 8260 29776
rect 8300 29724 8352 29776
rect 8484 29724 8536 29776
rect 8668 29724 8720 29776
rect 5172 29699 5224 29708
rect 5172 29665 5181 29699
rect 5181 29665 5215 29699
rect 5215 29665 5224 29699
rect 5172 29656 5224 29665
rect 6184 29656 6236 29708
rect 6736 29656 6788 29708
rect 7380 29699 7432 29708
rect 1400 29588 1452 29597
rect 3700 29588 3752 29640
rect 2596 29520 2648 29572
rect 4160 29520 4212 29572
rect 4804 29588 4856 29640
rect 4988 29588 5040 29640
rect 7380 29665 7389 29699
rect 7389 29665 7423 29699
rect 7423 29665 7432 29699
rect 11888 29724 11940 29776
rect 14188 29724 14240 29776
rect 17040 29792 17092 29844
rect 20628 29792 20680 29844
rect 20812 29835 20864 29844
rect 20812 29801 20821 29835
rect 20821 29801 20855 29835
rect 20855 29801 20864 29835
rect 20812 29792 20864 29801
rect 20996 29792 21048 29844
rect 23664 29792 23716 29844
rect 26700 29792 26752 29844
rect 30104 29792 30156 29844
rect 7380 29656 7432 29665
rect 5356 29520 5408 29572
rect 6368 29520 6420 29572
rect 4344 29452 4396 29504
rect 6184 29452 6236 29504
rect 7656 29588 7708 29640
rect 18604 29724 18656 29776
rect 19524 29724 19576 29776
rect 20904 29724 20956 29776
rect 21364 29724 21416 29776
rect 22836 29724 22888 29776
rect 25320 29724 25372 29776
rect 6828 29520 6880 29572
rect 8668 29520 8720 29572
rect 9220 29554 9272 29606
rect 10232 29588 10284 29640
rect 12992 29588 13044 29640
rect 14096 29588 14148 29640
rect 11520 29520 11572 29572
rect 15200 29588 15252 29640
rect 15660 29631 15712 29640
rect 15660 29597 15669 29631
rect 15669 29597 15703 29631
rect 15703 29597 15712 29631
rect 15660 29588 15712 29597
rect 18236 29656 18288 29708
rect 19248 29656 19300 29708
rect 24584 29656 24636 29708
rect 25688 29699 25740 29708
rect 25688 29665 25697 29699
rect 25697 29665 25731 29699
rect 25731 29665 25740 29699
rect 25688 29656 25740 29665
rect 26516 29699 26568 29708
rect 26516 29665 26525 29699
rect 26525 29665 26559 29699
rect 26559 29665 26568 29699
rect 26516 29656 26568 29665
rect 29920 29699 29972 29708
rect 29920 29665 29929 29699
rect 29929 29665 29963 29699
rect 29963 29665 29972 29699
rect 29920 29656 29972 29665
rect 17960 29631 18012 29640
rect 17960 29597 17969 29631
rect 17969 29597 18003 29631
rect 18003 29597 18012 29631
rect 17960 29588 18012 29597
rect 18328 29588 18380 29640
rect 16120 29520 16172 29572
rect 16304 29520 16356 29572
rect 18696 29520 18748 29572
rect 20720 29588 20772 29640
rect 20904 29520 20956 29572
rect 21548 29588 21600 29640
rect 25780 29631 25832 29640
rect 25780 29597 25789 29631
rect 25789 29597 25823 29631
rect 25823 29597 25832 29631
rect 25780 29588 25832 29597
rect 25964 29631 26016 29640
rect 25964 29597 25973 29631
rect 25973 29597 26007 29631
rect 26007 29597 26016 29631
rect 25964 29588 26016 29597
rect 27528 29588 27580 29640
rect 28724 29631 28776 29640
rect 28724 29597 28733 29631
rect 28733 29597 28767 29631
rect 28767 29597 28776 29631
rect 28724 29588 28776 29597
rect 28908 29631 28960 29640
rect 28908 29597 28917 29631
rect 28917 29597 28951 29631
rect 28951 29597 28960 29631
rect 28908 29588 28960 29597
rect 29276 29588 29328 29640
rect 30012 29588 30064 29640
rect 7932 29452 7984 29504
rect 8208 29452 8260 29504
rect 9220 29452 9272 29504
rect 9496 29495 9548 29504
rect 9496 29461 9505 29495
rect 9505 29461 9539 29495
rect 9539 29461 9548 29495
rect 9496 29452 9548 29461
rect 9864 29452 9916 29504
rect 12256 29452 12308 29504
rect 13176 29452 13228 29504
rect 17316 29452 17368 29504
rect 17684 29452 17736 29504
rect 20444 29452 20496 29504
rect 21916 29520 21968 29572
rect 23112 29520 23164 29572
rect 23480 29520 23532 29572
rect 26056 29520 26108 29572
rect 26608 29520 26660 29572
rect 29736 29520 29788 29572
rect 30380 29520 30432 29572
rect 22192 29452 22244 29504
rect 22928 29452 22980 29504
rect 23756 29495 23808 29504
rect 23756 29461 23765 29495
rect 23765 29461 23799 29495
rect 23799 29461 23808 29495
rect 23756 29452 23808 29461
rect 24400 29452 24452 29504
rect 24676 29452 24728 29504
rect 26424 29452 26476 29504
rect 30012 29452 30064 29504
rect 7288 29350 7340 29402
rect 17592 29350 17644 29402
rect 27896 29350 27948 29402
rect 3148 29248 3200 29300
rect 3700 29180 3752 29232
rect 4804 29248 4856 29300
rect 4896 29180 4948 29232
rect 3792 29155 3844 29164
rect 3792 29121 3801 29155
rect 3801 29121 3835 29155
rect 3835 29121 3844 29155
rect 3792 29112 3844 29121
rect 4252 29112 4304 29164
rect 4528 29112 4580 29164
rect 7472 29248 7524 29300
rect 9220 29248 9272 29300
rect 4160 29044 4212 29096
rect 7380 29112 7432 29164
rect 7932 29155 7984 29164
rect 7932 29121 7941 29155
rect 7941 29121 7975 29155
rect 7975 29121 7984 29155
rect 7932 29112 7984 29121
rect 9772 29180 9824 29232
rect 10232 29248 10284 29300
rect 11520 29248 11572 29300
rect 6828 29087 6880 29096
rect 6828 29053 6837 29087
rect 6837 29053 6871 29087
rect 6871 29053 6880 29087
rect 6828 29044 6880 29053
rect 7012 29044 7064 29096
rect 7472 29044 7524 29096
rect 11152 29112 11204 29164
rect 12900 29180 12952 29232
rect 13636 29180 13688 29232
rect 14832 29180 14884 29232
rect 12072 29112 12124 29164
rect 13452 29155 13504 29164
rect 13452 29121 13461 29155
rect 13461 29121 13495 29155
rect 13495 29121 13504 29155
rect 13452 29112 13504 29121
rect 15292 29112 15344 29164
rect 15660 29180 15712 29232
rect 17132 29248 17184 29300
rect 17776 29248 17828 29300
rect 20996 29248 21048 29300
rect 21916 29248 21968 29300
rect 12532 29044 12584 29096
rect 12992 29044 13044 29096
rect 2228 28951 2280 28960
rect 2228 28917 2237 28951
rect 2237 28917 2271 28951
rect 2271 28917 2280 28951
rect 2228 28908 2280 28917
rect 8208 28976 8260 29028
rect 10600 28976 10652 29028
rect 14096 29044 14148 29096
rect 14372 29087 14424 29096
rect 14372 29053 14381 29087
rect 14381 29053 14415 29087
rect 14415 29053 14424 29087
rect 14372 29044 14424 29053
rect 14648 29044 14700 29096
rect 15200 29044 15252 29096
rect 16672 29112 16724 29164
rect 17316 29155 17368 29164
rect 17316 29121 17325 29155
rect 17325 29121 17359 29155
rect 17359 29121 17368 29155
rect 17316 29112 17368 29121
rect 17408 29112 17460 29164
rect 17684 29112 17736 29164
rect 19432 29112 19484 29164
rect 17040 29044 17092 29096
rect 17960 29044 18012 29096
rect 18144 29044 18196 29096
rect 18696 29044 18748 29096
rect 22192 29248 22244 29300
rect 22928 29248 22980 29300
rect 24124 29248 24176 29300
rect 13912 28976 13964 29028
rect 14740 28976 14792 29028
rect 17132 28976 17184 29028
rect 18788 28976 18840 29028
rect 19248 28976 19300 29028
rect 20996 28976 21048 29028
rect 22468 29112 22520 29164
rect 22560 29112 22612 29164
rect 23112 29155 23164 29164
rect 22652 29044 22704 29096
rect 23112 29121 23121 29155
rect 23121 29121 23155 29155
rect 23155 29121 23164 29155
rect 23112 29112 23164 29121
rect 24124 29155 24176 29164
rect 24124 29121 24133 29155
rect 24133 29121 24167 29155
rect 24167 29121 24176 29155
rect 24124 29112 24176 29121
rect 23020 29044 23072 29096
rect 24216 29044 24268 29096
rect 24676 29112 24728 29164
rect 25872 29180 25924 29232
rect 24676 28976 24728 29028
rect 24952 29044 25004 29096
rect 25136 29044 25188 29096
rect 28080 29112 28132 29164
rect 28356 29155 28408 29164
rect 28356 29121 28365 29155
rect 28365 29121 28399 29155
rect 28399 29121 28408 29155
rect 28356 29112 28408 29121
rect 29276 29112 29328 29164
rect 26516 28976 26568 29028
rect 27160 29044 27212 29096
rect 27344 29087 27396 29096
rect 27344 29053 27353 29087
rect 27353 29053 27387 29087
rect 27387 29053 27396 29087
rect 27344 29044 27396 29053
rect 29184 29087 29236 29096
rect 29184 29053 29193 29087
rect 29193 29053 29227 29087
rect 29227 29053 29236 29087
rect 29184 29044 29236 29053
rect 30104 29155 30156 29164
rect 30104 29121 30113 29155
rect 30113 29121 30147 29155
rect 30147 29121 30156 29155
rect 30380 29155 30432 29164
rect 30104 29112 30156 29121
rect 30380 29121 30389 29155
rect 30389 29121 30423 29155
rect 30423 29121 30432 29155
rect 30380 29112 30432 29121
rect 27804 28976 27856 29028
rect 29828 29019 29880 29028
rect 29828 28985 29837 29019
rect 29837 28985 29871 29019
rect 29871 28985 29880 29019
rect 29828 28976 29880 28985
rect 4436 28908 4488 28960
rect 5172 28908 5224 28960
rect 8116 28908 8168 28960
rect 9128 28908 9180 28960
rect 9496 28908 9548 28960
rect 10508 28908 10560 28960
rect 11520 28908 11572 28960
rect 12716 28908 12768 28960
rect 20260 28908 20312 28960
rect 21180 28908 21232 28960
rect 22192 28908 22244 28960
rect 22468 28951 22520 28960
rect 22468 28917 22477 28951
rect 22477 28917 22511 28951
rect 22511 28917 22520 28951
rect 22468 28908 22520 28917
rect 24216 28908 24268 28960
rect 24584 28908 24636 28960
rect 25688 28908 25740 28960
rect 25964 28951 26016 28960
rect 25964 28917 25973 28951
rect 25973 28917 26007 28951
rect 26007 28917 26016 28951
rect 25964 28908 26016 28917
rect 26884 28908 26936 28960
rect 29736 28908 29788 28960
rect 30196 29087 30248 29096
rect 30196 29053 30230 29087
rect 30230 29053 30248 29087
rect 30196 29044 30248 29053
rect 30840 28908 30892 28960
rect 31024 28951 31076 28960
rect 31024 28917 31033 28951
rect 31033 28917 31067 28951
rect 31067 28917 31076 28951
rect 31024 28908 31076 28917
rect 2136 28806 2188 28858
rect 12440 28806 12492 28858
rect 22744 28806 22796 28858
rect 4528 28704 4580 28756
rect 8208 28704 8260 28756
rect 8944 28747 8996 28756
rect 8944 28713 8953 28747
rect 8953 28713 8987 28747
rect 8987 28713 8996 28747
rect 8944 28704 8996 28713
rect 10048 28747 10100 28756
rect 10048 28713 10057 28747
rect 10057 28713 10091 28747
rect 10091 28713 10100 28747
rect 10048 28704 10100 28713
rect 11152 28747 11204 28756
rect 11152 28713 11161 28747
rect 11161 28713 11195 28747
rect 11195 28713 11204 28747
rect 11152 28704 11204 28713
rect 11520 28747 11572 28756
rect 11520 28713 11529 28747
rect 11529 28713 11563 28747
rect 11563 28713 11572 28747
rect 11520 28704 11572 28713
rect 12072 28747 12124 28756
rect 12072 28713 12081 28747
rect 12081 28713 12115 28747
rect 12115 28713 12124 28747
rect 12072 28704 12124 28713
rect 12348 28704 12400 28756
rect 12624 28704 12676 28756
rect 14464 28704 14516 28756
rect 14832 28704 14884 28756
rect 3056 28636 3108 28688
rect 3792 28636 3844 28688
rect 7932 28636 7984 28688
rect 4436 28568 4488 28620
rect 5356 28611 5408 28620
rect 1400 28500 1452 28552
rect 2688 28500 2740 28552
rect 4344 28543 4396 28552
rect 4344 28509 4353 28543
rect 4353 28509 4387 28543
rect 4387 28509 4396 28543
rect 4344 28500 4396 28509
rect 5356 28577 5365 28611
rect 5365 28577 5399 28611
rect 5399 28577 5408 28611
rect 5356 28568 5408 28577
rect 8116 28568 8168 28620
rect 2228 28432 2280 28484
rect 6368 28500 6420 28552
rect 6644 28543 6696 28552
rect 6644 28509 6653 28543
rect 6653 28509 6687 28543
rect 6687 28509 6696 28543
rect 7932 28543 7984 28552
rect 6644 28500 6696 28509
rect 7932 28509 7941 28543
rect 7941 28509 7975 28543
rect 7975 28509 7984 28543
rect 7932 28500 7984 28509
rect 8208 28543 8260 28552
rect 8208 28509 8217 28543
rect 8217 28509 8251 28543
rect 8251 28509 8260 28543
rect 8208 28500 8260 28509
rect 9588 28636 9640 28688
rect 9772 28636 9824 28688
rect 10968 28636 11020 28688
rect 15200 28636 15252 28688
rect 15752 28704 15804 28756
rect 8760 28568 8812 28620
rect 6184 28432 6236 28484
rect 9220 28543 9272 28552
rect 9220 28509 9229 28543
rect 9229 28509 9263 28543
rect 9263 28509 9272 28543
rect 9404 28543 9456 28552
rect 9220 28500 9272 28509
rect 9404 28509 9413 28543
rect 9413 28509 9447 28543
rect 9447 28509 9456 28543
rect 9404 28500 9456 28509
rect 9680 28500 9732 28552
rect 10508 28543 10560 28552
rect 10508 28509 10517 28543
rect 10517 28509 10551 28543
rect 10551 28509 10560 28543
rect 10508 28500 10560 28509
rect 11152 28568 11204 28620
rect 11980 28500 12032 28552
rect 12072 28500 12124 28552
rect 12532 28543 12584 28552
rect 12532 28509 12541 28543
rect 12541 28509 12575 28543
rect 12575 28509 12584 28543
rect 12532 28500 12584 28509
rect 7380 28364 7432 28416
rect 11888 28432 11940 28484
rect 12808 28500 12860 28552
rect 13176 28432 13228 28484
rect 9496 28364 9548 28416
rect 9680 28364 9732 28416
rect 11060 28364 11112 28416
rect 11704 28364 11756 28416
rect 12164 28364 12216 28416
rect 13912 28432 13964 28484
rect 13728 28364 13780 28416
rect 14372 28500 14424 28552
rect 14648 28500 14700 28552
rect 18328 28704 18380 28756
rect 20720 28704 20772 28756
rect 21548 28704 21600 28756
rect 22376 28704 22428 28756
rect 23112 28704 23164 28756
rect 25504 28704 25556 28756
rect 26884 28747 26936 28756
rect 26884 28713 26893 28747
rect 26893 28713 26927 28747
rect 26927 28713 26936 28747
rect 26884 28704 26936 28713
rect 29000 28747 29052 28756
rect 18696 28679 18748 28688
rect 18696 28645 18705 28679
rect 18705 28645 18739 28679
rect 18739 28645 18748 28679
rect 18696 28636 18748 28645
rect 20260 28636 20312 28688
rect 15752 28543 15804 28552
rect 15752 28509 15761 28543
rect 15761 28509 15795 28543
rect 15795 28509 15804 28543
rect 15752 28500 15804 28509
rect 16304 28500 16356 28552
rect 17316 28500 17368 28552
rect 18052 28500 18104 28552
rect 19248 28543 19300 28552
rect 19248 28509 19257 28543
rect 19257 28509 19291 28543
rect 19291 28509 19300 28543
rect 19248 28500 19300 28509
rect 21916 28568 21968 28620
rect 22468 28568 22520 28620
rect 22928 28636 22980 28688
rect 21180 28500 21232 28552
rect 16764 28475 16816 28484
rect 16764 28441 16798 28475
rect 16798 28441 16816 28475
rect 16764 28432 16816 28441
rect 18512 28475 18564 28484
rect 18512 28441 18521 28475
rect 18521 28441 18555 28475
rect 18555 28441 18564 28475
rect 18512 28432 18564 28441
rect 20168 28432 20220 28484
rect 22652 28500 22704 28552
rect 24308 28636 24360 28688
rect 25320 28636 25372 28688
rect 25688 28636 25740 28688
rect 29000 28713 29009 28747
rect 29009 28713 29043 28747
rect 29043 28713 29052 28747
rect 29000 28704 29052 28713
rect 29736 28704 29788 28756
rect 30196 28704 30248 28756
rect 29092 28636 29144 28688
rect 24216 28568 24268 28620
rect 24768 28611 24820 28620
rect 14832 28364 14884 28416
rect 22836 28432 22888 28484
rect 23848 28500 23900 28552
rect 24768 28577 24777 28611
rect 24777 28577 24811 28611
rect 24811 28577 24820 28611
rect 24768 28568 24820 28577
rect 27620 28611 27672 28620
rect 27620 28577 27629 28611
rect 27629 28577 27663 28611
rect 27663 28577 27672 28611
rect 27620 28568 27672 28577
rect 25044 28500 25096 28552
rect 25412 28500 25464 28552
rect 25596 28543 25648 28552
rect 25596 28509 25605 28543
rect 25605 28509 25639 28543
rect 25639 28509 25648 28543
rect 25596 28500 25648 28509
rect 25780 28543 25832 28552
rect 25780 28509 25789 28543
rect 25789 28509 25823 28543
rect 25823 28509 25832 28543
rect 25780 28500 25832 28509
rect 26148 28500 26200 28552
rect 29920 28543 29972 28552
rect 29920 28509 29929 28543
rect 29929 28509 29963 28543
rect 29963 28509 29972 28543
rect 29920 28500 29972 28509
rect 30012 28500 30064 28552
rect 25228 28432 25280 28484
rect 25964 28432 26016 28484
rect 22008 28364 22060 28416
rect 22468 28364 22520 28416
rect 24492 28364 24544 28416
rect 24768 28364 24820 28416
rect 24860 28364 24912 28416
rect 26424 28364 26476 28416
rect 27068 28407 27120 28416
rect 27068 28373 27077 28407
rect 27077 28373 27111 28407
rect 27111 28373 27120 28407
rect 27068 28364 27120 28373
rect 28540 28432 28592 28484
rect 29184 28364 29236 28416
rect 31116 28364 31168 28416
rect 7288 28262 7340 28314
rect 17592 28262 17644 28314
rect 27896 28262 27948 28314
rect 1952 28160 2004 28212
rect 2412 28160 2464 28212
rect 8208 28160 8260 28212
rect 7748 28092 7800 28144
rect 2412 28024 2464 28076
rect 5540 28024 5592 28076
rect 7196 28024 7248 28076
rect 7932 28024 7984 28076
rect 9680 28203 9732 28212
rect 9680 28169 9689 28203
rect 9689 28169 9723 28203
rect 9723 28169 9732 28203
rect 9680 28160 9732 28169
rect 8760 28092 8812 28144
rect 11060 28160 11112 28212
rect 11612 28160 11664 28212
rect 11980 28160 12032 28212
rect 12348 28160 12400 28212
rect 12716 28160 12768 28212
rect 2320 27956 2372 28008
rect 5448 27956 5500 28008
rect 5724 27956 5776 28008
rect 6368 27999 6420 28008
rect 6368 27965 6377 27999
rect 6377 27965 6411 27999
rect 6411 27965 6420 27999
rect 6368 27956 6420 27965
rect 7472 27956 7524 28008
rect 8484 27956 8536 28008
rect 4344 27888 4396 27940
rect 5356 27888 5408 27940
rect 8116 27888 8168 27940
rect 9772 28024 9824 28076
rect 10508 28092 10560 28144
rect 14648 28160 14700 28212
rect 10232 28024 10284 28076
rect 10968 28067 11020 28076
rect 10968 28033 10977 28067
rect 10977 28033 11011 28067
rect 11011 28033 11020 28067
rect 10968 28024 11020 28033
rect 11612 28024 11664 28076
rect 11520 27956 11572 28008
rect 9772 27888 9824 27940
rect 1400 27820 1452 27872
rect 2320 27863 2372 27872
rect 2320 27829 2329 27863
rect 2329 27829 2363 27863
rect 2363 27829 2372 27863
rect 2320 27820 2372 27829
rect 2688 27820 2740 27872
rect 4252 27863 4304 27872
rect 4252 27829 4261 27863
rect 4261 27829 4295 27863
rect 4295 27829 4304 27863
rect 4252 27820 4304 27829
rect 5172 27863 5224 27872
rect 5172 27829 5181 27863
rect 5181 27829 5215 27863
rect 5215 27829 5224 27863
rect 5172 27820 5224 27829
rect 7840 27820 7892 27872
rect 8392 27820 8444 27872
rect 13636 28024 13688 28076
rect 14096 28024 14148 28076
rect 15384 28067 15436 28076
rect 12808 27888 12860 27940
rect 13452 27888 13504 27940
rect 13084 27863 13136 27872
rect 13084 27829 13093 27863
rect 13093 27829 13127 27863
rect 13127 27829 13136 27863
rect 13084 27820 13136 27829
rect 15384 28033 15393 28067
rect 15393 28033 15427 28067
rect 15427 28033 15436 28067
rect 15384 28024 15436 28033
rect 16212 28160 16264 28212
rect 17132 28160 17184 28212
rect 17960 28160 18012 28212
rect 18328 28135 18380 28144
rect 18328 28101 18337 28135
rect 18337 28101 18371 28135
rect 18371 28101 18380 28135
rect 18328 28092 18380 28101
rect 19340 28160 19392 28212
rect 18696 28092 18748 28144
rect 19524 28092 19576 28144
rect 22468 28160 22520 28212
rect 24216 28203 24268 28212
rect 24216 28169 24225 28203
rect 24225 28169 24259 28203
rect 24259 28169 24268 28203
rect 24216 28160 24268 28169
rect 24308 28160 24360 28212
rect 24584 28160 24636 28212
rect 24768 28160 24820 28212
rect 24400 28092 24452 28144
rect 25044 28160 25096 28212
rect 25228 28160 25280 28212
rect 15292 27956 15344 28008
rect 16948 28024 17000 28076
rect 16120 27956 16172 28008
rect 18236 28024 18288 28076
rect 18972 28024 19024 28076
rect 19800 27999 19852 28008
rect 19800 27965 19809 27999
rect 19809 27965 19843 27999
rect 19843 27965 19852 27999
rect 19800 27956 19852 27965
rect 21088 28067 21140 28076
rect 21088 28033 21097 28067
rect 21097 28033 21131 28067
rect 21131 28033 21140 28067
rect 21088 28024 21140 28033
rect 21180 27956 21232 28008
rect 21548 27956 21600 28008
rect 22560 28024 22612 28076
rect 23204 28067 23256 28076
rect 23204 28033 23213 28067
rect 23213 28033 23247 28067
rect 23247 28033 23256 28067
rect 23204 28024 23256 28033
rect 24584 28067 24636 28076
rect 24584 28033 24593 28067
rect 24593 28033 24627 28067
rect 24627 28033 24636 28067
rect 24584 28024 24636 28033
rect 24676 28067 24728 28076
rect 24676 28033 24685 28067
rect 24685 28033 24719 28067
rect 24719 28033 24728 28067
rect 24676 28024 24728 28033
rect 25688 28024 25740 28076
rect 25872 28024 25924 28076
rect 27068 28024 27120 28076
rect 27804 28160 27856 28212
rect 28448 28160 28500 28212
rect 31208 28160 31260 28212
rect 27344 28092 27396 28144
rect 28172 28092 28224 28144
rect 31024 28092 31076 28144
rect 22652 27956 22704 28008
rect 23388 27956 23440 28008
rect 24124 27956 24176 28008
rect 25780 27956 25832 28008
rect 14556 27820 14608 27872
rect 16304 27820 16356 27872
rect 18972 27820 19024 27872
rect 19064 27820 19116 27872
rect 20076 27820 20128 27872
rect 21272 27888 21324 27940
rect 22468 27888 22520 27940
rect 24952 27888 25004 27940
rect 25596 27888 25648 27940
rect 26240 27999 26292 28008
rect 26240 27965 26249 27999
rect 26249 27965 26283 27999
rect 26283 27965 26292 27999
rect 26240 27956 26292 27965
rect 29736 28067 29788 28076
rect 28448 27999 28500 28008
rect 28448 27965 28457 27999
rect 28457 27965 28491 27999
rect 28491 27965 28500 27999
rect 28448 27956 28500 27965
rect 26884 27888 26936 27940
rect 29276 27888 29328 27940
rect 23756 27820 23808 27872
rect 24584 27820 24636 27872
rect 24676 27820 24728 27872
rect 24860 27820 24912 27872
rect 27344 27863 27396 27872
rect 27344 27829 27353 27863
rect 27353 27829 27387 27863
rect 27387 27829 27396 27863
rect 27344 27820 27396 27829
rect 28632 27820 28684 27872
rect 28724 27820 28776 27872
rect 29736 28033 29745 28067
rect 29745 28033 29779 28067
rect 29779 28033 29788 28067
rect 29736 28024 29788 28033
rect 30656 28024 30708 28076
rect 30748 28067 30800 28076
rect 30748 28033 30757 28067
rect 30757 28033 30791 28067
rect 30791 28033 30800 28067
rect 30748 28024 30800 28033
rect 30932 28067 30984 28076
rect 30932 28033 30941 28067
rect 30941 28033 30975 28067
rect 30975 28033 30984 28067
rect 30932 28024 30984 28033
rect 31300 28024 31352 28076
rect 30564 27820 30616 27872
rect 2136 27718 2188 27770
rect 12440 27718 12492 27770
rect 22744 27718 22796 27770
rect 2596 27591 2648 27600
rect 2596 27557 2605 27591
rect 2605 27557 2639 27591
rect 2639 27557 2648 27591
rect 2596 27548 2648 27557
rect 4436 27616 4488 27668
rect 4344 27591 4396 27600
rect 4344 27557 4353 27591
rect 4353 27557 4387 27591
rect 4387 27557 4396 27591
rect 4344 27548 4396 27557
rect 6920 27548 6972 27600
rect 7472 27548 7524 27600
rect 8484 27616 8536 27668
rect 9128 27616 9180 27668
rect 11612 27616 11664 27668
rect 11796 27616 11848 27668
rect 10416 27548 10468 27600
rect 13912 27548 13964 27600
rect 14188 27548 14240 27600
rect 15752 27616 15804 27668
rect 21088 27616 21140 27668
rect 23020 27616 23072 27668
rect 23296 27616 23348 27668
rect 23572 27616 23624 27668
rect 24492 27659 24544 27668
rect 24492 27625 24501 27659
rect 24501 27625 24535 27659
rect 24535 27625 24544 27659
rect 24492 27616 24544 27625
rect 25872 27616 25924 27668
rect 26240 27616 26292 27668
rect 27436 27616 27488 27668
rect 28540 27659 28592 27668
rect 1584 27480 1636 27532
rect 2872 27480 2924 27532
rect 3056 27523 3108 27532
rect 3056 27489 3065 27523
rect 3065 27489 3099 27523
rect 3099 27489 3108 27523
rect 3056 27480 3108 27489
rect 4252 27480 4304 27532
rect 2780 27455 2832 27464
rect 2780 27421 2789 27455
rect 2789 27421 2823 27455
rect 2823 27421 2832 27455
rect 4160 27455 4212 27464
rect 2780 27412 2832 27421
rect 4160 27421 4169 27455
rect 4169 27421 4203 27455
rect 4203 27421 4212 27455
rect 4160 27412 4212 27421
rect 5172 27455 5224 27464
rect 5172 27421 5206 27455
rect 5206 27421 5224 27455
rect 4344 27344 4396 27396
rect 5172 27412 5224 27421
rect 7840 27480 7892 27532
rect 5080 27344 5132 27396
rect 2780 27276 2832 27328
rect 4068 27276 4120 27328
rect 7012 27276 7064 27328
rect 7932 27455 7984 27464
rect 7932 27421 7941 27455
rect 7941 27421 7975 27455
rect 7975 27421 7984 27455
rect 8208 27455 8260 27464
rect 7932 27412 7984 27421
rect 8208 27421 8217 27455
rect 8217 27421 8251 27455
rect 8251 27421 8260 27455
rect 8208 27412 8260 27421
rect 9220 27480 9272 27532
rect 10232 27480 10284 27532
rect 9496 27412 9548 27464
rect 10508 27412 10560 27464
rect 12808 27480 12860 27532
rect 14372 27480 14424 27532
rect 11888 27412 11940 27464
rect 12072 27412 12124 27464
rect 12900 27455 12952 27464
rect 12900 27421 12909 27455
rect 12909 27421 12943 27455
rect 12943 27421 12952 27455
rect 12900 27412 12952 27421
rect 13084 27455 13136 27464
rect 13084 27421 13093 27455
rect 13093 27421 13127 27455
rect 13127 27421 13136 27455
rect 13084 27412 13136 27421
rect 13176 27412 13228 27464
rect 14004 27412 14056 27464
rect 14556 27412 14608 27464
rect 14740 27412 14792 27464
rect 15200 27412 15252 27464
rect 17316 27455 17368 27464
rect 17316 27421 17325 27455
rect 17325 27421 17359 27455
rect 17359 27421 17368 27455
rect 17316 27412 17368 27421
rect 19064 27480 19116 27532
rect 12808 27344 12860 27396
rect 15108 27344 15160 27396
rect 18604 27412 18656 27464
rect 21272 27548 21324 27600
rect 22560 27548 22612 27600
rect 23204 27548 23256 27600
rect 24308 27548 24360 27600
rect 25596 27548 25648 27600
rect 28540 27625 28549 27659
rect 28549 27625 28583 27659
rect 28583 27625 28592 27659
rect 28540 27616 28592 27625
rect 28632 27616 28684 27668
rect 29828 27616 29880 27668
rect 31300 27659 31352 27668
rect 31300 27625 31309 27659
rect 31309 27625 31343 27659
rect 31343 27625 31352 27659
rect 31300 27616 31352 27625
rect 22652 27480 22704 27532
rect 23848 27480 23900 27532
rect 25688 27480 25740 27532
rect 29184 27480 29236 27532
rect 29920 27523 29972 27532
rect 29920 27489 29929 27523
rect 29929 27489 29963 27523
rect 29963 27489 29972 27523
rect 29920 27480 29972 27489
rect 17684 27344 17736 27396
rect 18788 27344 18840 27396
rect 20076 27412 20128 27464
rect 20720 27455 20772 27464
rect 20720 27421 20729 27455
rect 20729 27421 20763 27455
rect 20763 27421 20772 27455
rect 20720 27412 20772 27421
rect 21916 27412 21968 27464
rect 22376 27412 22428 27464
rect 22928 27412 22980 27464
rect 23388 27412 23440 27464
rect 24124 27412 24176 27464
rect 24400 27455 24452 27464
rect 24400 27421 24409 27455
rect 24409 27421 24443 27455
rect 24443 27421 24452 27455
rect 24400 27412 24452 27421
rect 25504 27412 25556 27464
rect 26700 27455 26752 27464
rect 26700 27421 26709 27455
rect 26709 27421 26743 27455
rect 26743 27421 26752 27455
rect 26700 27412 26752 27421
rect 28724 27455 28776 27464
rect 28724 27421 28733 27455
rect 28733 27421 28767 27455
rect 28767 27421 28776 27455
rect 28724 27412 28776 27421
rect 28908 27455 28960 27464
rect 28908 27421 28917 27455
rect 28917 27421 28951 27455
rect 28951 27421 28960 27455
rect 28908 27412 28960 27421
rect 19984 27344 20036 27396
rect 20904 27344 20956 27396
rect 21732 27344 21784 27396
rect 25136 27344 25188 27396
rect 26148 27344 26200 27396
rect 26792 27344 26844 27396
rect 30380 27344 30432 27396
rect 8944 27319 8996 27328
rect 8944 27285 8953 27319
rect 8953 27285 8987 27319
rect 8987 27285 8996 27319
rect 8944 27276 8996 27285
rect 9496 27276 9548 27328
rect 18420 27276 18472 27328
rect 19064 27276 19116 27328
rect 23572 27276 23624 27328
rect 24768 27276 24820 27328
rect 28448 27276 28500 27328
rect 29368 27276 29420 27328
rect 30104 27276 30156 27328
rect 7288 27174 7340 27226
rect 17592 27174 17644 27226
rect 27896 27174 27948 27226
rect 1860 27072 1912 27124
rect 2596 27072 2648 27124
rect 7196 27115 7248 27124
rect 7196 27081 7205 27115
rect 7205 27081 7239 27115
rect 7239 27081 7248 27115
rect 7196 27072 7248 27081
rect 2688 27004 2740 27056
rect 9496 27072 9548 27124
rect 10324 27072 10376 27124
rect 11244 27072 11296 27124
rect 11612 27072 11664 27124
rect 12532 27072 12584 27124
rect 12900 27072 12952 27124
rect 13176 27072 13228 27124
rect 13636 27072 13688 27124
rect 17040 27072 17092 27124
rect 17684 27115 17736 27124
rect 17684 27081 17693 27115
rect 17693 27081 17727 27115
rect 17727 27081 17736 27115
rect 17684 27072 17736 27081
rect 1676 26979 1728 26988
rect 1676 26945 1710 26979
rect 1710 26945 1728 26979
rect 1676 26936 1728 26945
rect 4068 26979 4120 26988
rect 4068 26945 4102 26979
rect 4102 26945 4120 26979
rect 4068 26936 4120 26945
rect 8944 27004 8996 27056
rect 7380 26979 7432 26988
rect 1400 26911 1452 26920
rect 1400 26877 1409 26911
rect 1409 26877 1443 26911
rect 1443 26877 1452 26911
rect 1400 26868 1452 26877
rect 1768 26732 1820 26784
rect 2688 26732 2740 26784
rect 2872 26732 2924 26784
rect 3148 26732 3200 26784
rect 5724 26800 5776 26852
rect 7380 26945 7389 26979
rect 7389 26945 7423 26979
rect 7423 26945 7432 26979
rect 7380 26936 7432 26945
rect 7472 26936 7524 26988
rect 7840 26936 7892 26988
rect 8760 26936 8812 26988
rect 11428 26936 11480 26988
rect 11704 26936 11756 26988
rect 11888 26945 11897 26972
rect 11897 26945 11931 26972
rect 11931 26945 11940 26972
rect 11888 26920 11940 26945
rect 8116 26911 8168 26920
rect 8116 26877 8125 26911
rect 8125 26877 8159 26911
rect 8159 26877 8168 26911
rect 8116 26868 8168 26877
rect 10876 26868 10928 26920
rect 5632 26775 5684 26784
rect 5632 26741 5641 26775
rect 5641 26741 5675 26775
rect 5675 26741 5684 26775
rect 5632 26732 5684 26741
rect 6460 26732 6512 26784
rect 7380 26732 7432 26784
rect 7656 26732 7708 26784
rect 9220 26800 9272 26852
rect 9772 26800 9824 26852
rect 10600 26800 10652 26852
rect 11244 26800 11296 26852
rect 11888 26800 11940 26852
rect 12256 26936 12308 26988
rect 12716 26936 12768 26988
rect 12900 26936 12952 26988
rect 13452 27004 13504 27056
rect 15292 27004 15344 27056
rect 19984 27004 20036 27056
rect 22928 27072 22980 27124
rect 23480 27072 23532 27124
rect 25044 27072 25096 27124
rect 26792 27072 26844 27124
rect 27344 27072 27396 27124
rect 30380 27115 30432 27124
rect 23388 27004 23440 27056
rect 25872 27004 25924 27056
rect 26332 27004 26384 27056
rect 13728 26979 13780 26988
rect 13728 26945 13737 26979
rect 13737 26945 13771 26979
rect 13771 26945 13780 26979
rect 13728 26936 13780 26945
rect 14004 26979 14056 26988
rect 14004 26945 14013 26979
rect 14013 26945 14047 26979
rect 14047 26945 14056 26979
rect 14004 26936 14056 26945
rect 14372 26936 14424 26988
rect 14188 26868 14240 26920
rect 15384 26936 15436 26988
rect 16212 26936 16264 26988
rect 16948 26979 17000 26988
rect 16948 26945 16957 26979
rect 16957 26945 16991 26979
rect 16991 26945 17000 26979
rect 16948 26936 17000 26945
rect 17868 26979 17920 26988
rect 17868 26945 17877 26979
rect 17877 26945 17911 26979
rect 17911 26945 17920 26979
rect 17868 26936 17920 26945
rect 18604 26936 18656 26988
rect 19064 26979 19116 26988
rect 19064 26945 19073 26979
rect 19073 26945 19107 26979
rect 19107 26945 19116 26979
rect 19064 26936 19116 26945
rect 20076 26979 20128 26988
rect 20076 26945 20085 26979
rect 20085 26945 20119 26979
rect 20119 26945 20128 26979
rect 20076 26936 20128 26945
rect 20720 26936 20772 26988
rect 20996 26979 21048 26988
rect 20996 26945 21005 26979
rect 21005 26945 21039 26979
rect 21039 26945 21048 26979
rect 20996 26936 21048 26945
rect 21824 26979 21876 26988
rect 21824 26945 21833 26979
rect 21833 26945 21867 26979
rect 21867 26945 21876 26979
rect 21824 26936 21876 26945
rect 22376 26936 22428 26988
rect 22836 26936 22888 26988
rect 23480 26936 23532 26988
rect 16488 26868 16540 26920
rect 16580 26800 16632 26852
rect 19340 26868 19392 26920
rect 19708 26868 19760 26920
rect 20812 26868 20864 26920
rect 21180 26868 21232 26920
rect 24124 26911 24176 26920
rect 24124 26877 24133 26911
rect 24133 26877 24167 26911
rect 24167 26877 24176 26911
rect 24124 26868 24176 26877
rect 26424 26911 26476 26920
rect 26424 26877 26433 26911
rect 26433 26877 26467 26911
rect 26467 26877 26476 26911
rect 26424 26868 26476 26877
rect 19064 26800 19116 26852
rect 11060 26732 11112 26784
rect 13912 26775 13964 26784
rect 13912 26741 13921 26775
rect 13921 26741 13955 26775
rect 13955 26741 13964 26775
rect 13912 26732 13964 26741
rect 14004 26732 14056 26784
rect 16672 26732 16724 26784
rect 17132 26775 17184 26784
rect 17132 26741 17141 26775
rect 17141 26741 17175 26775
rect 17175 26741 17184 26775
rect 17132 26732 17184 26741
rect 18420 26732 18472 26784
rect 19892 26775 19944 26784
rect 19892 26741 19901 26775
rect 19901 26741 19935 26775
rect 19935 26741 19944 26775
rect 19892 26732 19944 26741
rect 21088 26732 21140 26784
rect 22192 26732 22244 26784
rect 23756 26732 23808 26784
rect 24768 26732 24820 26784
rect 25228 26732 25280 26784
rect 27528 26936 27580 26988
rect 27988 26936 28040 26988
rect 29184 26979 29236 26988
rect 29184 26945 29193 26979
rect 29193 26945 29227 26979
rect 29227 26945 29236 26979
rect 29184 26936 29236 26945
rect 30380 27081 30389 27115
rect 30389 27081 30423 27115
rect 30423 27081 30432 27115
rect 30380 27072 30432 27081
rect 29920 26936 29972 26988
rect 30564 26979 30616 26988
rect 30564 26945 30573 26979
rect 30573 26945 30607 26979
rect 30607 26945 30616 26979
rect 30564 26936 30616 26945
rect 28540 26911 28592 26920
rect 28540 26877 28549 26911
rect 28549 26877 28583 26911
rect 28583 26877 28592 26911
rect 28540 26868 28592 26877
rect 29460 26911 29512 26920
rect 29460 26877 29469 26911
rect 29469 26877 29503 26911
rect 29503 26877 29512 26911
rect 29460 26868 29512 26877
rect 31024 26868 31076 26920
rect 28908 26800 28960 26852
rect 28080 26775 28132 26784
rect 28080 26741 28089 26775
rect 28089 26741 28123 26775
rect 28123 26741 28132 26775
rect 28080 26732 28132 26741
rect 28448 26775 28500 26784
rect 28448 26741 28457 26775
rect 28457 26741 28491 26775
rect 28491 26741 28500 26775
rect 28448 26732 28500 26741
rect 28632 26732 28684 26784
rect 2136 26630 2188 26682
rect 12440 26630 12492 26682
rect 22744 26630 22796 26682
rect 4160 26528 4212 26580
rect 5540 26571 5592 26580
rect 5540 26537 5549 26571
rect 5549 26537 5583 26571
rect 5583 26537 5592 26571
rect 5540 26528 5592 26537
rect 3332 26460 3384 26512
rect 2504 26392 2556 26444
rect 4528 26392 4580 26444
rect 1860 26324 1912 26376
rect 1492 26256 1544 26308
rect 2872 26324 2924 26376
rect 3240 26367 3292 26376
rect 3240 26333 3249 26367
rect 3249 26333 3283 26367
rect 3283 26333 3292 26367
rect 3240 26324 3292 26333
rect 4068 26324 4120 26376
rect 4712 26324 4764 26376
rect 4988 26324 5040 26376
rect 5724 26528 5776 26580
rect 7104 26528 7156 26580
rect 7840 26528 7892 26580
rect 8392 26528 8444 26580
rect 11612 26528 11664 26580
rect 16948 26528 17000 26580
rect 17132 26528 17184 26580
rect 11796 26460 11848 26512
rect 14004 26460 14056 26512
rect 14096 26460 14148 26512
rect 15476 26460 15528 26512
rect 18236 26460 18288 26512
rect 20996 26528 21048 26580
rect 23020 26528 23072 26580
rect 23480 26528 23532 26580
rect 23756 26503 23808 26512
rect 23756 26469 23765 26503
rect 23765 26469 23799 26503
rect 23799 26469 23808 26503
rect 23756 26460 23808 26469
rect 12532 26392 12584 26444
rect 12716 26392 12768 26444
rect 12900 26435 12952 26444
rect 12900 26401 12909 26435
rect 12909 26401 12943 26435
rect 12943 26401 12952 26435
rect 12900 26392 12952 26401
rect 13544 26392 13596 26444
rect 5816 26324 5868 26376
rect 4804 26256 4856 26308
rect 6368 26324 6420 26376
rect 6828 26324 6880 26376
rect 7012 26367 7064 26376
rect 7012 26333 7046 26367
rect 7046 26333 7064 26367
rect 7012 26324 7064 26333
rect 8116 26324 8168 26376
rect 11520 26324 11572 26376
rect 11796 26324 11848 26376
rect 11888 26324 11940 26376
rect 12256 26324 12308 26376
rect 6920 26256 6972 26308
rect 9772 26256 9824 26308
rect 13636 26324 13688 26376
rect 13820 26324 13872 26376
rect 15292 26367 15344 26376
rect 15292 26333 15301 26367
rect 15301 26333 15335 26367
rect 15335 26333 15344 26367
rect 15292 26324 15344 26333
rect 19708 26392 19760 26444
rect 21640 26392 21692 26444
rect 26700 26528 26752 26580
rect 29920 26571 29972 26580
rect 29920 26537 29929 26571
rect 29929 26537 29963 26571
rect 29963 26537 29972 26571
rect 29920 26528 29972 26537
rect 30932 26528 30984 26580
rect 29736 26460 29788 26512
rect 15660 26324 15712 26376
rect 15844 26324 15896 26376
rect 16672 26324 16724 26376
rect 17132 26324 17184 26376
rect 17408 26324 17460 26376
rect 17500 26324 17552 26376
rect 17960 26324 18012 26376
rect 18696 26367 18748 26376
rect 18696 26333 18705 26367
rect 18705 26333 18739 26367
rect 18739 26333 18748 26367
rect 18696 26324 18748 26333
rect 20812 26324 20864 26376
rect 21732 26324 21784 26376
rect 12716 26256 12768 26308
rect 14464 26299 14516 26308
rect 14464 26265 14473 26299
rect 14473 26265 14507 26299
rect 14507 26265 14516 26299
rect 14464 26256 14516 26265
rect 14924 26256 14976 26308
rect 15384 26256 15436 26308
rect 16580 26256 16632 26308
rect 18236 26256 18288 26308
rect 1768 26188 1820 26240
rect 3792 26231 3844 26240
rect 3792 26197 3801 26231
rect 3801 26197 3835 26231
rect 3835 26197 3844 26231
rect 3792 26188 3844 26197
rect 5080 26188 5132 26240
rect 9680 26188 9732 26240
rect 10876 26188 10928 26240
rect 11612 26188 11664 26240
rect 11704 26188 11756 26240
rect 14188 26188 14240 26240
rect 16672 26188 16724 26240
rect 19892 26256 19944 26308
rect 22652 26324 22704 26376
rect 22928 26367 22980 26376
rect 21180 26231 21232 26240
rect 21180 26197 21189 26231
rect 21189 26197 21223 26231
rect 21223 26197 21232 26231
rect 21180 26188 21232 26197
rect 22468 26256 22520 26308
rect 22928 26333 22937 26367
rect 22937 26333 22971 26367
rect 22971 26333 22980 26367
rect 22928 26324 22980 26333
rect 24124 26392 24176 26444
rect 24492 26324 24544 26376
rect 25044 26367 25096 26376
rect 22836 26188 22888 26240
rect 25044 26333 25053 26367
rect 25053 26333 25087 26367
rect 25087 26333 25096 26367
rect 25044 26324 25096 26333
rect 29000 26392 29052 26444
rect 30104 26392 30156 26444
rect 26792 26324 26844 26376
rect 27712 26324 27764 26376
rect 29092 26324 29144 26376
rect 30564 26324 30616 26376
rect 25228 26188 25280 26240
rect 26976 26256 27028 26308
rect 30104 26256 30156 26308
rect 26332 26188 26384 26240
rect 26516 26188 26568 26240
rect 29736 26188 29788 26240
rect 7288 26086 7340 26138
rect 17592 26086 17644 26138
rect 27896 26086 27948 26138
rect 1676 25984 1728 26036
rect 2228 25984 2280 26036
rect 1308 25916 1360 25968
rect 2780 25959 2832 25968
rect 2780 25925 2814 25959
rect 2814 25925 2832 25959
rect 2780 25916 2832 25925
rect 4344 25959 4396 25968
rect 4344 25925 4353 25959
rect 4353 25925 4387 25959
rect 4387 25925 4396 25959
rect 4344 25916 4396 25925
rect 9404 25984 9456 26036
rect 6920 25916 6972 25968
rect 9588 25916 9640 25968
rect 1768 25891 1820 25900
rect 1768 25857 1777 25891
rect 1777 25857 1811 25891
rect 1811 25857 1820 25891
rect 1768 25848 1820 25857
rect 1860 25848 1912 25900
rect 4804 25891 4856 25900
rect 4804 25857 4813 25891
rect 4813 25857 4847 25891
rect 4847 25857 4856 25891
rect 4804 25848 4856 25857
rect 7748 25891 7800 25900
rect 1676 25780 1728 25832
rect 1400 25712 1452 25764
rect 6276 25780 6328 25832
rect 7748 25857 7757 25891
rect 7757 25857 7791 25891
rect 7791 25857 7800 25891
rect 7748 25848 7800 25857
rect 9312 25848 9364 25900
rect 12808 25984 12860 26036
rect 12900 26027 12952 26036
rect 12900 25993 12909 26027
rect 12909 25993 12943 26027
rect 12943 25993 12952 26027
rect 12900 25984 12952 25993
rect 14832 25984 14884 26036
rect 16672 25984 16724 26036
rect 11060 25916 11112 25968
rect 10600 25848 10652 25900
rect 6000 25712 6052 25764
rect 1584 25644 1636 25696
rect 4436 25644 4488 25696
rect 6552 25644 6604 25696
rect 6736 25644 6788 25696
rect 10324 25780 10376 25832
rect 10876 25848 10928 25900
rect 11520 25891 11572 25900
rect 11520 25857 11529 25891
rect 11529 25857 11563 25891
rect 11563 25857 11572 25891
rect 11520 25848 11572 25857
rect 11612 25848 11664 25900
rect 12348 25916 12400 25968
rect 12716 25916 12768 25968
rect 13636 25916 13688 25968
rect 16120 25916 16172 25968
rect 13544 25891 13596 25900
rect 13544 25857 13553 25891
rect 13553 25857 13587 25891
rect 13587 25857 13596 25891
rect 13544 25848 13596 25857
rect 14556 25891 14608 25900
rect 14556 25857 14565 25891
rect 14565 25857 14599 25891
rect 14599 25857 14608 25891
rect 14556 25848 14608 25857
rect 15200 25848 15252 25900
rect 16304 25848 16356 25900
rect 18512 25984 18564 26036
rect 20076 25984 20128 26036
rect 21824 25984 21876 26036
rect 16948 25916 17000 25968
rect 19432 25916 19484 25968
rect 18052 25848 18104 25900
rect 19524 25891 19576 25900
rect 19524 25857 19533 25891
rect 19533 25857 19567 25891
rect 19567 25857 19576 25891
rect 19524 25848 19576 25857
rect 20628 25891 20680 25900
rect 12808 25780 12860 25832
rect 13636 25780 13688 25832
rect 16856 25780 16908 25832
rect 17316 25780 17368 25832
rect 19432 25780 19484 25832
rect 20628 25857 20637 25891
rect 20637 25857 20671 25891
rect 20671 25857 20680 25891
rect 20628 25848 20680 25857
rect 21180 25848 21232 25900
rect 24492 25984 24544 26036
rect 23756 25916 23808 25968
rect 27712 25848 27764 25900
rect 28632 25848 28684 25900
rect 30104 25916 30156 25968
rect 21640 25780 21692 25832
rect 22192 25780 22244 25832
rect 23204 25780 23256 25832
rect 8208 25712 8260 25764
rect 11060 25712 11112 25764
rect 9220 25644 9272 25696
rect 9312 25644 9364 25696
rect 10232 25644 10284 25696
rect 12624 25644 12676 25696
rect 13084 25644 13136 25696
rect 13912 25644 13964 25696
rect 14924 25644 14976 25696
rect 15844 25644 15896 25696
rect 17408 25644 17460 25696
rect 18696 25644 18748 25696
rect 23572 25644 23624 25696
rect 29000 25687 29052 25696
rect 29000 25653 29009 25687
rect 29009 25653 29043 25687
rect 29043 25653 29052 25687
rect 29000 25644 29052 25653
rect 31116 25644 31168 25696
rect 2136 25542 2188 25594
rect 12440 25542 12492 25594
rect 22744 25542 22796 25594
rect 3976 25440 4028 25492
rect 6552 25440 6604 25492
rect 11704 25440 11756 25492
rect 11980 25440 12032 25492
rect 13636 25440 13688 25492
rect 15200 25483 15252 25492
rect 15200 25449 15209 25483
rect 15209 25449 15243 25483
rect 15243 25449 15252 25483
rect 15200 25440 15252 25449
rect 18052 25483 18104 25492
rect 18052 25449 18061 25483
rect 18061 25449 18095 25483
rect 18095 25449 18104 25483
rect 18052 25440 18104 25449
rect 19524 25440 19576 25492
rect 2964 25372 3016 25424
rect 1492 25236 1544 25288
rect 2228 25304 2280 25356
rect 2872 25347 2924 25356
rect 2872 25313 2881 25347
rect 2881 25313 2915 25347
rect 2915 25313 2924 25347
rect 2872 25304 2924 25313
rect 6552 25304 6604 25356
rect 9404 25372 9456 25424
rect 9220 25347 9272 25356
rect 9220 25313 9229 25347
rect 9229 25313 9263 25347
rect 9263 25313 9272 25347
rect 9220 25304 9272 25313
rect 9772 25304 9824 25356
rect 10600 25304 10652 25356
rect 4712 25279 4764 25288
rect 2228 25168 2280 25220
rect 3976 25168 4028 25220
rect 4712 25245 4721 25279
rect 4721 25245 4755 25279
rect 4755 25245 4764 25279
rect 4712 25236 4764 25245
rect 4988 25279 5040 25288
rect 4988 25245 4997 25279
rect 4997 25245 5031 25279
rect 5031 25245 5040 25279
rect 4988 25236 5040 25245
rect 5080 25236 5132 25288
rect 7196 25279 7248 25288
rect 7196 25245 7205 25279
rect 7205 25245 7239 25279
rect 7239 25245 7248 25279
rect 7196 25236 7248 25245
rect 8208 25279 8260 25288
rect 8208 25245 8217 25279
rect 8217 25245 8251 25279
rect 8251 25245 8260 25279
rect 8208 25236 8260 25245
rect 9312 25279 9364 25288
rect 9312 25245 9321 25279
rect 9321 25245 9355 25279
rect 9355 25245 9364 25279
rect 9312 25236 9364 25245
rect 9404 25279 9456 25288
rect 9404 25245 9413 25279
rect 9413 25245 9447 25279
rect 9447 25245 9456 25279
rect 9404 25236 9456 25245
rect 9680 25236 9732 25288
rect 12716 25304 12768 25356
rect 12992 25304 13044 25356
rect 11428 25279 11480 25288
rect 1492 25100 1544 25152
rect 1768 25100 1820 25152
rect 3792 25100 3844 25152
rect 5172 25100 5224 25152
rect 10232 25100 10284 25152
rect 10600 25100 10652 25152
rect 10968 25100 11020 25152
rect 11428 25245 11437 25279
rect 11437 25245 11471 25279
rect 11471 25245 11480 25279
rect 11428 25236 11480 25245
rect 12072 25279 12124 25288
rect 12072 25245 12081 25279
rect 12081 25245 12115 25279
rect 12115 25245 12124 25279
rect 12072 25236 12124 25245
rect 12256 25236 12308 25288
rect 12532 25279 12584 25288
rect 11336 25168 11388 25220
rect 11980 25168 12032 25220
rect 12532 25245 12541 25279
rect 12541 25245 12575 25279
rect 12575 25245 12584 25279
rect 12532 25236 12584 25245
rect 12808 25236 12860 25288
rect 15108 25372 15160 25424
rect 16028 25372 16080 25424
rect 20904 25372 20956 25424
rect 23756 25440 23808 25492
rect 24492 25440 24544 25492
rect 31208 25440 31260 25492
rect 27160 25372 27212 25424
rect 15292 25304 15344 25356
rect 11612 25100 11664 25152
rect 12348 25100 12400 25152
rect 13636 25168 13688 25220
rect 13176 25100 13228 25152
rect 14740 25279 14792 25288
rect 14004 25168 14056 25220
rect 14740 25245 14749 25279
rect 14749 25245 14783 25279
rect 14783 25245 14792 25279
rect 14740 25236 14792 25245
rect 15384 25279 15436 25288
rect 15384 25245 15393 25279
rect 15393 25245 15427 25279
rect 15427 25245 15436 25279
rect 15384 25236 15436 25245
rect 16396 25304 16448 25356
rect 20628 25304 20680 25356
rect 18420 25279 18472 25288
rect 18420 25245 18429 25279
rect 18429 25245 18463 25279
rect 18463 25245 18472 25279
rect 18420 25236 18472 25245
rect 19432 25279 19484 25288
rect 15752 25168 15804 25220
rect 16304 25211 16356 25220
rect 16304 25177 16313 25211
rect 16313 25177 16347 25211
rect 16347 25177 16356 25211
rect 16304 25168 16356 25177
rect 16672 25168 16724 25220
rect 18328 25168 18380 25220
rect 19432 25245 19441 25279
rect 19441 25245 19475 25279
rect 19475 25245 19484 25279
rect 19432 25236 19484 25245
rect 19708 25279 19760 25288
rect 19708 25245 19717 25279
rect 19717 25245 19751 25279
rect 19751 25245 19760 25279
rect 19708 25236 19760 25245
rect 22468 25304 22520 25356
rect 24768 25304 24820 25356
rect 18696 25168 18748 25220
rect 22100 25236 22152 25288
rect 22560 25279 22612 25288
rect 22560 25245 22569 25279
rect 22569 25245 22603 25279
rect 22603 25245 22612 25279
rect 22560 25236 22612 25245
rect 23388 25236 23440 25288
rect 25228 25236 25280 25288
rect 26332 25236 26384 25288
rect 26516 25236 26568 25288
rect 28264 25236 28316 25288
rect 21640 25168 21692 25220
rect 24124 25168 24176 25220
rect 16488 25100 16540 25152
rect 20260 25100 20312 25152
rect 20996 25100 21048 25152
rect 22468 25100 22520 25152
rect 23572 25143 23624 25152
rect 23572 25109 23581 25143
rect 23581 25109 23615 25143
rect 23615 25109 23624 25143
rect 23572 25100 23624 25109
rect 24952 25168 25004 25220
rect 24308 25100 24360 25152
rect 25320 25100 25372 25152
rect 27160 25100 27212 25152
rect 27804 25100 27856 25152
rect 30288 25168 30340 25220
rect 7288 24998 7340 25050
rect 17592 24998 17644 25050
rect 27896 24998 27948 25050
rect 2228 24896 2280 24948
rect 5080 24896 5132 24948
rect 6368 24896 6420 24948
rect 7196 24896 7248 24948
rect 9404 24896 9456 24948
rect 1676 24871 1728 24880
rect 1676 24837 1685 24871
rect 1685 24837 1719 24871
rect 1719 24837 1728 24871
rect 1676 24828 1728 24837
rect 2596 24828 2648 24880
rect 2228 24760 2280 24812
rect 2964 24803 3016 24812
rect 2964 24769 2973 24803
rect 2973 24769 3007 24803
rect 3007 24769 3016 24803
rect 2964 24760 3016 24769
rect 4436 24828 4488 24880
rect 9588 24828 9640 24880
rect 10600 24896 10652 24948
rect 11796 24896 11848 24948
rect 12164 24896 12216 24948
rect 16488 24896 16540 24948
rect 18052 24896 18104 24948
rect 18420 24896 18472 24948
rect 19248 24896 19300 24948
rect 22192 24939 22244 24948
rect 22192 24905 22225 24939
rect 22225 24905 22244 24939
rect 22192 24896 22244 24905
rect 22560 24896 22612 24948
rect 4896 24760 4948 24812
rect 6368 24803 6420 24812
rect 6368 24769 6377 24803
rect 6377 24769 6411 24803
rect 6411 24769 6420 24803
rect 6368 24760 6420 24769
rect 2596 24692 2648 24744
rect 3516 24692 3568 24744
rect 6644 24803 6696 24812
rect 6644 24769 6653 24803
rect 6653 24769 6687 24803
rect 6687 24769 6696 24803
rect 6644 24760 6696 24769
rect 6828 24760 6880 24812
rect 8208 24760 8260 24812
rect 8668 24760 8720 24812
rect 9128 24760 9180 24812
rect 9404 24760 9456 24812
rect 10416 24828 10468 24880
rect 10784 24828 10836 24880
rect 11520 24828 11572 24880
rect 13084 24871 13136 24880
rect 11612 24760 11664 24812
rect 13084 24837 13118 24871
rect 13118 24837 13136 24871
rect 13084 24828 13136 24837
rect 14924 24871 14976 24880
rect 14924 24837 14933 24871
rect 14933 24837 14967 24871
rect 14967 24837 14976 24871
rect 14924 24828 14976 24837
rect 15476 24828 15528 24880
rect 15660 24828 15712 24880
rect 16212 24871 16264 24880
rect 16212 24837 16221 24871
rect 16221 24837 16255 24871
rect 16255 24837 16264 24871
rect 16212 24828 16264 24837
rect 22468 24828 22520 24880
rect 22652 24871 22704 24880
rect 22652 24837 22661 24871
rect 22661 24837 22695 24871
rect 22695 24837 22704 24871
rect 22652 24828 22704 24837
rect 13636 24760 13688 24812
rect 1952 24667 2004 24676
rect 1952 24633 1961 24667
rect 1961 24633 1995 24667
rect 1995 24633 2004 24667
rect 1952 24624 2004 24633
rect 6828 24624 6880 24676
rect 6552 24556 6604 24608
rect 9312 24624 9364 24676
rect 10324 24692 10376 24744
rect 10508 24692 10560 24744
rect 12808 24735 12860 24744
rect 12808 24701 12817 24735
rect 12817 24701 12851 24735
rect 12851 24701 12860 24735
rect 12808 24692 12860 24701
rect 14464 24760 14516 24812
rect 16948 24760 17000 24812
rect 18328 24760 18380 24812
rect 19432 24803 19484 24812
rect 16028 24692 16080 24744
rect 17316 24692 17368 24744
rect 19432 24769 19441 24803
rect 19441 24769 19475 24803
rect 19475 24769 19484 24803
rect 19432 24760 19484 24769
rect 19708 24803 19760 24812
rect 19708 24769 19717 24803
rect 19717 24769 19751 24803
rect 19751 24769 19760 24803
rect 19708 24760 19760 24769
rect 20996 24803 21048 24812
rect 19800 24692 19852 24744
rect 20996 24769 21005 24803
rect 21005 24769 21039 24803
rect 21039 24769 21048 24803
rect 20996 24760 21048 24769
rect 21088 24760 21140 24812
rect 22100 24760 22152 24812
rect 24676 24828 24728 24880
rect 23296 24803 23348 24812
rect 23296 24769 23305 24803
rect 23305 24769 23339 24803
rect 23339 24769 23348 24803
rect 23296 24760 23348 24769
rect 23480 24803 23532 24812
rect 23480 24769 23489 24803
rect 23489 24769 23523 24803
rect 23523 24769 23532 24803
rect 23480 24760 23532 24769
rect 25228 24803 25280 24812
rect 25228 24769 25237 24803
rect 25237 24769 25271 24803
rect 25271 24769 25280 24803
rect 25228 24760 25280 24769
rect 25504 24803 25556 24812
rect 25504 24769 25513 24803
rect 25513 24769 25547 24803
rect 25547 24769 25556 24803
rect 25504 24760 25556 24769
rect 22560 24692 22612 24744
rect 8484 24599 8536 24608
rect 8484 24565 8493 24599
rect 8493 24565 8527 24599
rect 8527 24565 8536 24599
rect 8484 24556 8536 24565
rect 9128 24556 9180 24608
rect 15936 24624 15988 24676
rect 17868 24624 17920 24676
rect 22008 24624 22060 24676
rect 23388 24692 23440 24744
rect 26516 24828 26568 24880
rect 26792 24760 26844 24812
rect 26976 24803 27028 24812
rect 26976 24769 26985 24803
rect 26985 24769 27019 24803
rect 27019 24769 27028 24803
rect 26976 24760 27028 24769
rect 27160 24803 27212 24812
rect 27160 24769 27169 24803
rect 27169 24769 27203 24803
rect 27203 24769 27212 24803
rect 27160 24760 27212 24769
rect 27436 24803 27488 24812
rect 27436 24769 27445 24803
rect 27445 24769 27479 24803
rect 27479 24769 27488 24803
rect 27436 24760 27488 24769
rect 28172 24760 28224 24812
rect 29092 24803 29144 24812
rect 29092 24769 29101 24803
rect 29101 24769 29135 24803
rect 29135 24769 29144 24803
rect 29092 24760 29144 24769
rect 25872 24624 25924 24676
rect 14096 24556 14148 24608
rect 14188 24599 14240 24608
rect 14188 24565 14197 24599
rect 14197 24565 14231 24599
rect 14231 24565 14240 24599
rect 14188 24556 14240 24565
rect 14924 24556 14976 24608
rect 18512 24556 18564 24608
rect 19156 24556 19208 24608
rect 20904 24556 20956 24608
rect 24768 24556 24820 24608
rect 27712 24692 27764 24744
rect 29736 24803 29788 24812
rect 29736 24769 29745 24803
rect 29745 24769 29779 24803
rect 29779 24769 29788 24803
rect 29736 24760 29788 24769
rect 30012 24760 30064 24812
rect 30656 24803 30708 24812
rect 30656 24769 30665 24803
rect 30665 24769 30699 24803
rect 30699 24769 30708 24803
rect 30656 24760 30708 24769
rect 31116 24760 31168 24812
rect 30564 24692 30616 24744
rect 27436 24556 27488 24608
rect 28448 24556 28500 24608
rect 2136 24454 2188 24506
rect 12440 24454 12492 24506
rect 22744 24454 22796 24506
rect 2688 24352 2740 24404
rect 3792 24395 3844 24404
rect 3792 24361 3801 24395
rect 3801 24361 3835 24395
rect 3835 24361 3844 24395
rect 3792 24352 3844 24361
rect 4896 24352 4948 24404
rect 5356 24395 5408 24404
rect 5356 24361 5365 24395
rect 5365 24361 5399 24395
rect 5399 24361 5408 24395
rect 5356 24352 5408 24361
rect 5540 24352 5592 24404
rect 8760 24352 8812 24404
rect 9404 24352 9456 24404
rect 9588 24352 9640 24404
rect 6368 24284 6420 24336
rect 1676 24216 1728 24268
rect 2780 24216 2832 24268
rect 4528 24216 4580 24268
rect 2688 24191 2740 24200
rect 2688 24157 2697 24191
rect 2697 24157 2731 24191
rect 2731 24157 2740 24191
rect 2688 24148 2740 24157
rect 5172 24191 5224 24200
rect 1584 24012 1636 24064
rect 5172 24157 5181 24191
rect 5181 24157 5215 24191
rect 5215 24157 5224 24191
rect 5172 24148 5224 24157
rect 6736 24216 6788 24268
rect 6920 24148 6972 24200
rect 7656 24148 7708 24200
rect 8484 24148 8536 24200
rect 8944 24148 8996 24200
rect 9128 24148 9180 24200
rect 9680 24148 9732 24200
rect 6092 24080 6144 24132
rect 7196 24080 7248 24132
rect 4528 24012 4580 24064
rect 5080 24012 5132 24064
rect 9864 24012 9916 24064
rect 11428 24352 11480 24404
rect 12624 24352 12676 24404
rect 13636 24352 13688 24404
rect 13820 24284 13872 24336
rect 14096 24352 14148 24404
rect 15108 24284 15160 24336
rect 15660 24284 15712 24336
rect 19156 24284 19208 24336
rect 19248 24284 19300 24336
rect 20260 24327 20312 24336
rect 10508 24216 10560 24268
rect 13084 24216 13136 24268
rect 14004 24216 14056 24268
rect 14188 24216 14240 24268
rect 14740 24216 14792 24268
rect 16856 24259 16908 24268
rect 10600 24148 10652 24200
rect 10968 24191 11020 24200
rect 10968 24157 10977 24191
rect 10977 24157 11011 24191
rect 11011 24157 11020 24191
rect 10968 24148 11020 24157
rect 11336 24148 11388 24200
rect 13728 24148 13780 24200
rect 14924 24148 14976 24200
rect 15108 24191 15160 24200
rect 15108 24157 15117 24191
rect 15117 24157 15151 24191
rect 15151 24157 15160 24191
rect 15108 24148 15160 24157
rect 15844 24191 15896 24200
rect 15844 24157 15853 24191
rect 15853 24157 15887 24191
rect 15887 24157 15896 24191
rect 15844 24148 15896 24157
rect 15936 24148 15988 24200
rect 16856 24225 16865 24259
rect 16865 24225 16899 24259
rect 16899 24225 16908 24259
rect 16856 24216 16908 24225
rect 20260 24293 20269 24327
rect 20269 24293 20303 24327
rect 20303 24293 20312 24327
rect 20260 24284 20312 24293
rect 20812 24259 20864 24268
rect 20812 24225 20821 24259
rect 20821 24225 20855 24259
rect 20855 24225 20864 24259
rect 20812 24216 20864 24225
rect 22192 24395 22244 24404
rect 22192 24361 22201 24395
rect 22201 24361 22235 24395
rect 22235 24361 22244 24395
rect 25872 24395 25924 24404
rect 22192 24352 22244 24361
rect 25872 24361 25881 24395
rect 25881 24361 25915 24395
rect 25915 24361 25924 24395
rect 25872 24352 25924 24361
rect 29184 24352 29236 24404
rect 22652 24327 22704 24336
rect 22652 24293 22661 24327
rect 22661 24293 22695 24327
rect 22695 24293 22704 24327
rect 22652 24284 22704 24293
rect 27620 24284 27672 24336
rect 28540 24284 28592 24336
rect 23296 24259 23348 24268
rect 11428 24080 11480 24132
rect 11796 24123 11848 24132
rect 11796 24089 11805 24123
rect 11805 24089 11839 24123
rect 11839 24089 11848 24123
rect 11796 24080 11848 24089
rect 12164 24080 12216 24132
rect 10784 24055 10836 24064
rect 10784 24021 10793 24055
rect 10793 24021 10827 24055
rect 10827 24021 10836 24055
rect 10784 24012 10836 24021
rect 12808 24012 12860 24064
rect 14004 24012 14056 24064
rect 14924 24055 14976 24064
rect 14924 24021 14933 24055
rect 14933 24021 14967 24055
rect 14967 24021 14976 24055
rect 14924 24012 14976 24021
rect 16212 24055 16264 24064
rect 16212 24021 16221 24055
rect 16221 24021 16255 24055
rect 16255 24021 16264 24055
rect 16212 24012 16264 24021
rect 17500 24080 17552 24132
rect 20076 24148 20128 24200
rect 20904 24148 20956 24200
rect 22652 24148 22704 24200
rect 22836 24148 22888 24200
rect 23296 24225 23305 24259
rect 23305 24225 23339 24259
rect 23339 24225 23348 24259
rect 23296 24216 23348 24225
rect 27344 24216 27396 24268
rect 23204 24148 23256 24200
rect 24216 24148 24268 24200
rect 17960 24012 18012 24064
rect 18328 24012 18380 24064
rect 19340 24012 19392 24064
rect 20260 24080 20312 24132
rect 21548 24080 21600 24132
rect 23112 24055 23164 24064
rect 23112 24021 23121 24055
rect 23121 24021 23155 24055
rect 23155 24021 23164 24055
rect 23112 24012 23164 24021
rect 24676 24080 24728 24132
rect 27436 24080 27488 24132
rect 27528 24080 27580 24132
rect 28724 24148 28776 24200
rect 29000 24148 29052 24200
rect 30012 24148 30064 24200
rect 30380 24148 30432 24200
rect 30656 24148 30708 24200
rect 30472 24080 30524 24132
rect 31208 24148 31260 24200
rect 27804 24012 27856 24064
rect 30840 24012 30892 24064
rect 7288 23910 7340 23962
rect 17592 23910 17644 23962
rect 27896 23910 27948 23962
rect 1308 23808 1360 23860
rect 1492 23808 1544 23860
rect 2780 23851 2832 23860
rect 2780 23817 2789 23851
rect 2789 23817 2823 23851
rect 2823 23817 2832 23851
rect 2780 23808 2832 23817
rect 3700 23740 3752 23792
rect 1400 23715 1452 23724
rect 1400 23681 1409 23715
rect 1409 23681 1443 23715
rect 1443 23681 1452 23715
rect 1400 23672 1452 23681
rect 1492 23672 1544 23724
rect 2228 23672 2280 23724
rect 5540 23808 5592 23860
rect 5724 23808 5776 23860
rect 6644 23808 6696 23860
rect 6920 23808 6972 23860
rect 8944 23851 8996 23860
rect 8944 23817 8953 23851
rect 8953 23817 8987 23851
rect 8987 23817 8996 23851
rect 8944 23808 8996 23817
rect 9588 23808 9640 23860
rect 10600 23808 10652 23860
rect 11060 23808 11112 23860
rect 12164 23851 12216 23860
rect 12164 23817 12173 23851
rect 12173 23817 12207 23851
rect 12207 23817 12216 23851
rect 12164 23808 12216 23817
rect 15384 23808 15436 23860
rect 16764 23808 16816 23860
rect 19524 23808 19576 23860
rect 4068 23740 4120 23792
rect 5724 23672 5776 23724
rect 6184 23672 6236 23724
rect 6368 23672 6420 23724
rect 8300 23740 8352 23792
rect 9680 23740 9732 23792
rect 4988 23604 5040 23656
rect 5264 23604 5316 23656
rect 6552 23604 6604 23656
rect 2964 23536 3016 23588
rect 4712 23536 4764 23588
rect 5448 23536 5500 23588
rect 6644 23536 6696 23588
rect 2688 23468 2740 23520
rect 3792 23511 3844 23520
rect 3792 23477 3801 23511
rect 3801 23477 3835 23511
rect 3835 23477 3844 23511
rect 3792 23468 3844 23477
rect 4160 23468 4212 23520
rect 4804 23468 4856 23520
rect 5172 23468 5224 23520
rect 6828 23468 6880 23520
rect 9864 23672 9916 23724
rect 10324 23715 10376 23724
rect 10324 23681 10333 23715
rect 10333 23681 10367 23715
rect 10367 23681 10376 23715
rect 10324 23672 10376 23681
rect 11428 23740 11480 23792
rect 14004 23740 14056 23792
rect 14924 23740 14976 23792
rect 15752 23740 15804 23792
rect 10508 23715 10560 23724
rect 10508 23681 10517 23715
rect 10517 23681 10551 23715
rect 10551 23681 10560 23715
rect 10508 23672 10560 23681
rect 12532 23604 12584 23656
rect 12900 23604 12952 23656
rect 15844 23672 15896 23724
rect 17868 23740 17920 23792
rect 19892 23740 19944 23792
rect 28356 23808 28408 23860
rect 30288 23808 30340 23860
rect 14280 23604 14332 23656
rect 18604 23672 18656 23724
rect 20260 23672 20312 23724
rect 20720 23740 20772 23792
rect 21272 23740 21324 23792
rect 21916 23740 21968 23792
rect 20628 23715 20680 23724
rect 20628 23681 20637 23715
rect 20637 23681 20671 23715
rect 20671 23681 20680 23715
rect 20628 23672 20680 23681
rect 10232 23468 10284 23520
rect 12808 23536 12860 23588
rect 23664 23672 23716 23724
rect 25228 23715 25280 23724
rect 25228 23681 25237 23715
rect 25237 23681 25271 23715
rect 25271 23681 25280 23715
rect 25504 23715 25556 23724
rect 25228 23672 25280 23681
rect 22468 23604 22520 23656
rect 22836 23647 22888 23656
rect 22836 23613 22845 23647
rect 22845 23613 22879 23647
rect 22879 23613 22888 23647
rect 22836 23604 22888 23613
rect 15752 23511 15804 23520
rect 15752 23477 15761 23511
rect 15761 23477 15795 23511
rect 15795 23477 15804 23511
rect 15752 23468 15804 23477
rect 15844 23468 15896 23520
rect 16948 23468 17000 23520
rect 17408 23468 17460 23520
rect 18604 23468 18656 23520
rect 20444 23511 20496 23520
rect 20444 23477 20453 23511
rect 20453 23477 20487 23511
rect 20487 23477 20496 23511
rect 20444 23468 20496 23477
rect 22100 23536 22152 23588
rect 24124 23536 24176 23588
rect 22008 23511 22060 23520
rect 22008 23477 22017 23511
rect 22017 23477 22051 23511
rect 22051 23477 22060 23511
rect 22008 23468 22060 23477
rect 25136 23536 25188 23588
rect 25504 23681 25513 23715
rect 25513 23681 25547 23715
rect 25547 23681 25556 23715
rect 25504 23672 25556 23681
rect 25596 23672 25648 23724
rect 26240 23715 26292 23724
rect 26240 23681 26249 23715
rect 26249 23681 26283 23715
rect 26283 23681 26292 23715
rect 26240 23672 26292 23681
rect 27160 23715 27212 23724
rect 27160 23681 27169 23715
rect 27169 23681 27203 23715
rect 27203 23681 27212 23715
rect 27160 23672 27212 23681
rect 27436 23715 27488 23724
rect 27436 23681 27445 23715
rect 27445 23681 27479 23715
rect 27479 23681 27488 23715
rect 27436 23672 27488 23681
rect 27620 23715 27672 23724
rect 27620 23681 27629 23715
rect 27629 23681 27663 23715
rect 27663 23681 27672 23715
rect 27620 23672 27672 23681
rect 28264 23672 28316 23724
rect 28908 23672 28960 23724
rect 30840 23715 30892 23724
rect 30840 23681 30849 23715
rect 30849 23681 30883 23715
rect 30883 23681 30892 23715
rect 30840 23672 30892 23681
rect 30932 23672 30984 23724
rect 26424 23604 26476 23656
rect 28172 23604 28224 23656
rect 25872 23536 25924 23588
rect 27436 23536 27488 23588
rect 30380 23604 30432 23656
rect 31116 23647 31168 23656
rect 31116 23613 31125 23647
rect 31125 23613 31159 23647
rect 31159 23613 31168 23647
rect 31116 23604 31168 23613
rect 24768 23468 24820 23520
rect 26240 23468 26292 23520
rect 2136 23366 2188 23418
rect 12440 23366 12492 23418
rect 22744 23366 22796 23418
rect 2596 23307 2648 23316
rect 2596 23273 2605 23307
rect 2605 23273 2639 23307
rect 2639 23273 2648 23307
rect 2596 23264 2648 23273
rect 4804 23264 4856 23316
rect 5356 23264 5408 23316
rect 8024 23307 8076 23316
rect 8024 23273 8033 23307
rect 8033 23273 8067 23307
rect 8067 23273 8076 23307
rect 8024 23264 8076 23273
rect 8208 23264 8260 23316
rect 12532 23264 12584 23316
rect 13360 23264 13412 23316
rect 14924 23264 14976 23316
rect 3976 23196 4028 23248
rect 8300 23196 8352 23248
rect 10784 23196 10836 23248
rect 13544 23196 13596 23248
rect 3792 23128 3844 23180
rect 4436 23171 4488 23180
rect 4436 23137 4445 23171
rect 4445 23137 4479 23171
rect 4479 23137 4488 23171
rect 4436 23128 4488 23137
rect 5264 23128 5316 23180
rect 3056 23103 3108 23112
rect 3056 23069 3065 23103
rect 3065 23069 3099 23103
rect 3099 23069 3108 23103
rect 3056 23060 3108 23069
rect 4160 23103 4212 23112
rect 4160 23069 4169 23103
rect 4169 23069 4203 23103
rect 4203 23069 4212 23103
rect 4160 23060 4212 23069
rect 5356 23060 5408 23112
rect 5816 23060 5868 23112
rect 6736 23128 6788 23180
rect 6644 23103 6696 23112
rect 6644 23069 6653 23103
rect 6653 23069 6687 23103
rect 6687 23069 6696 23103
rect 6644 23060 6696 23069
rect 7932 23103 7984 23112
rect 7932 23069 7941 23103
rect 7941 23069 7975 23103
rect 7975 23069 7984 23103
rect 7932 23060 7984 23069
rect 9312 23103 9364 23112
rect 9312 23069 9321 23103
rect 9321 23069 9355 23103
rect 9355 23069 9364 23103
rect 9312 23060 9364 23069
rect 9588 23103 9640 23112
rect 9588 23069 9597 23103
rect 9597 23069 9631 23103
rect 9631 23069 9640 23103
rect 9588 23060 9640 23069
rect 10232 23103 10284 23112
rect 10232 23069 10241 23103
rect 10241 23069 10275 23103
rect 10275 23069 10284 23103
rect 10232 23060 10284 23069
rect 10876 23128 10928 23180
rect 14648 23196 14700 23248
rect 17684 23264 17736 23316
rect 15200 23196 15252 23248
rect 17316 23196 17368 23248
rect 19432 23264 19484 23316
rect 19892 23264 19944 23316
rect 23480 23264 23532 23316
rect 24676 23264 24728 23316
rect 24952 23264 25004 23316
rect 27988 23307 28040 23316
rect 27988 23273 27997 23307
rect 27997 23273 28031 23307
rect 28031 23273 28040 23307
rect 27988 23264 28040 23273
rect 29184 23196 29236 23248
rect 10784 23060 10836 23112
rect 12808 23060 12860 23112
rect 2228 22992 2280 23044
rect 2964 23035 3016 23044
rect 2964 23001 2973 23035
rect 2973 23001 3007 23035
rect 3007 23001 3016 23035
rect 2964 22992 3016 23001
rect 4160 22924 4212 22976
rect 10968 22992 11020 23044
rect 12164 22992 12216 23044
rect 12256 22992 12308 23044
rect 13176 23060 13228 23112
rect 13728 23060 13780 23112
rect 16212 23128 16264 23180
rect 13820 22992 13872 23044
rect 14740 23060 14792 23112
rect 16672 23103 16724 23112
rect 16672 23069 16681 23103
rect 16681 23069 16715 23103
rect 16715 23069 16724 23103
rect 16672 23060 16724 23069
rect 18236 23128 18288 23180
rect 20904 23128 20956 23180
rect 21088 23171 21140 23180
rect 21088 23137 21097 23171
rect 21097 23137 21131 23171
rect 21131 23137 21140 23171
rect 21088 23128 21140 23137
rect 24124 23128 24176 23180
rect 27160 23128 27212 23180
rect 17040 23060 17092 23112
rect 18144 23103 18196 23112
rect 18144 23069 18153 23103
rect 18153 23069 18187 23103
rect 18187 23069 18196 23103
rect 18144 23060 18196 23069
rect 18328 23103 18380 23112
rect 18328 23069 18337 23103
rect 18337 23069 18371 23103
rect 18371 23069 18380 23103
rect 18328 23060 18380 23069
rect 19248 23103 19300 23112
rect 19248 23069 19257 23103
rect 19257 23069 19291 23103
rect 19291 23069 19300 23103
rect 19248 23060 19300 23069
rect 19340 23060 19392 23112
rect 25136 23060 25188 23112
rect 27252 23103 27304 23112
rect 5448 22924 5500 22976
rect 6460 22924 6512 22976
rect 7104 22924 7156 22976
rect 7840 22924 7892 22976
rect 9128 22967 9180 22976
rect 9128 22933 9137 22967
rect 9137 22933 9171 22967
rect 9171 22933 9180 22967
rect 9128 22924 9180 22933
rect 12900 22924 12952 22976
rect 13544 22924 13596 22976
rect 14096 22967 14148 22976
rect 14096 22933 14105 22967
rect 14105 22933 14139 22967
rect 14139 22933 14148 22967
rect 14096 22924 14148 22933
rect 14372 22924 14424 22976
rect 15752 22992 15804 23044
rect 19984 22992 20036 23044
rect 20720 22992 20772 23044
rect 23388 22992 23440 23044
rect 24308 22992 24360 23044
rect 25780 23035 25832 23044
rect 25780 23001 25789 23035
rect 25789 23001 25823 23035
rect 25823 23001 25832 23035
rect 25780 22992 25832 23001
rect 15844 22967 15896 22976
rect 15844 22933 15853 22967
rect 15853 22933 15887 22967
rect 15887 22933 15896 22967
rect 15844 22924 15896 22933
rect 16672 22924 16724 22976
rect 17868 22924 17920 22976
rect 18236 22924 18288 22976
rect 19800 22924 19852 22976
rect 22468 22967 22520 22976
rect 22468 22933 22477 22967
rect 22477 22933 22511 22967
rect 22511 22933 22520 22967
rect 22468 22924 22520 22933
rect 23940 22924 23992 22976
rect 25044 22967 25096 22976
rect 25044 22933 25069 22967
rect 25069 22933 25096 22967
rect 25044 22924 25096 22933
rect 26148 22924 26200 22976
rect 27252 23069 27261 23103
rect 27261 23069 27295 23103
rect 27295 23069 27304 23103
rect 27252 23060 27304 23069
rect 27804 23128 27856 23180
rect 27436 22992 27488 23044
rect 29460 23060 29512 23112
rect 29276 22992 29328 23044
rect 27160 22924 27212 22976
rect 30564 22924 30616 22976
rect 31300 22967 31352 22976
rect 31300 22933 31309 22967
rect 31309 22933 31343 22967
rect 31343 22933 31352 22967
rect 31300 22924 31352 22933
rect 7288 22822 7340 22874
rect 17592 22822 17644 22874
rect 27896 22822 27948 22874
rect 1492 22763 1544 22772
rect 1492 22729 1501 22763
rect 1501 22729 1535 22763
rect 1535 22729 1544 22763
rect 1492 22720 1544 22729
rect 1676 22720 1728 22772
rect 3056 22720 3108 22772
rect 6644 22720 6696 22772
rect 1676 22627 1728 22636
rect 1676 22593 1685 22627
rect 1685 22593 1719 22627
rect 1719 22593 1728 22627
rect 1676 22584 1728 22593
rect 4804 22695 4856 22704
rect 4804 22661 4813 22695
rect 4813 22661 4847 22695
rect 4847 22661 4856 22695
rect 4804 22652 4856 22661
rect 3424 22584 3476 22636
rect 3792 22627 3844 22636
rect 3792 22593 3801 22627
rect 3801 22593 3835 22627
rect 3835 22593 3844 22627
rect 3792 22584 3844 22593
rect 4068 22627 4120 22636
rect 4068 22593 4077 22627
rect 4077 22593 4111 22627
rect 4111 22593 4120 22627
rect 4068 22584 4120 22593
rect 4620 22627 4672 22636
rect 4620 22593 4629 22627
rect 4629 22593 4663 22627
rect 4663 22593 4672 22627
rect 4620 22584 4672 22593
rect 5448 22627 5500 22636
rect 5448 22593 5457 22627
rect 5457 22593 5491 22627
rect 5491 22593 5500 22627
rect 5448 22584 5500 22593
rect 6828 22652 6880 22704
rect 7656 22652 7708 22704
rect 9128 22652 9180 22704
rect 9312 22720 9364 22772
rect 10140 22720 10192 22772
rect 12072 22720 12124 22772
rect 13452 22720 13504 22772
rect 13544 22720 13596 22772
rect 15108 22763 15160 22772
rect 15108 22729 15117 22763
rect 15117 22729 15151 22763
rect 15151 22729 15160 22763
rect 15108 22720 15160 22729
rect 16580 22720 16632 22772
rect 17132 22720 17184 22772
rect 17500 22720 17552 22772
rect 18788 22763 18840 22772
rect 18788 22729 18797 22763
rect 18797 22729 18831 22763
rect 18831 22729 18840 22763
rect 18788 22720 18840 22729
rect 2596 22516 2648 22568
rect 2228 22448 2280 22500
rect 3056 22559 3108 22568
rect 3056 22525 3065 22559
rect 3065 22525 3099 22559
rect 3099 22525 3108 22559
rect 3056 22516 3108 22525
rect 4252 22516 4304 22568
rect 5908 22516 5960 22568
rect 8116 22584 8168 22636
rect 9772 22584 9824 22636
rect 9956 22584 10008 22636
rect 10324 22584 10376 22636
rect 4988 22448 5040 22500
rect 9680 22448 9732 22500
rect 14096 22652 14148 22704
rect 14280 22652 14332 22704
rect 17776 22652 17828 22704
rect 19892 22720 19944 22772
rect 20720 22763 20772 22772
rect 20720 22729 20729 22763
rect 20729 22729 20763 22763
rect 20763 22729 20772 22763
rect 20720 22720 20772 22729
rect 21180 22720 21232 22772
rect 21456 22720 21508 22772
rect 21916 22720 21968 22772
rect 24308 22720 24360 22772
rect 24584 22720 24636 22772
rect 26424 22720 26476 22772
rect 29460 22720 29512 22772
rect 29828 22720 29880 22772
rect 10968 22584 11020 22636
rect 15292 22627 15344 22636
rect 11152 22516 11204 22568
rect 12256 22516 12308 22568
rect 12808 22559 12860 22568
rect 12808 22525 12817 22559
rect 12817 22525 12851 22559
rect 12851 22525 12860 22559
rect 12808 22516 12860 22525
rect 15292 22593 15301 22627
rect 15301 22593 15335 22627
rect 15335 22593 15344 22627
rect 15292 22584 15344 22593
rect 15476 22584 15528 22636
rect 15752 22627 15804 22636
rect 15752 22593 15761 22627
rect 15761 22593 15795 22627
rect 15795 22593 15804 22627
rect 15752 22584 15804 22593
rect 16764 22627 16816 22636
rect 16764 22593 16773 22627
rect 16773 22593 16807 22627
rect 16807 22593 16816 22627
rect 16764 22584 16816 22593
rect 16948 22627 17000 22636
rect 16948 22593 16957 22627
rect 16957 22593 16991 22627
rect 16991 22593 17000 22627
rect 16948 22584 17000 22593
rect 17868 22627 17920 22636
rect 17040 22516 17092 22568
rect 11244 22448 11296 22500
rect 3608 22423 3660 22432
rect 3608 22389 3617 22423
rect 3617 22389 3651 22423
rect 3651 22389 3660 22423
rect 3608 22380 3660 22389
rect 5816 22380 5868 22432
rect 6736 22380 6788 22432
rect 10508 22380 10560 22432
rect 12624 22380 12676 22432
rect 14096 22448 14148 22500
rect 17868 22593 17877 22627
rect 17877 22593 17911 22627
rect 17911 22593 17920 22627
rect 17868 22584 17920 22593
rect 18236 22584 18288 22636
rect 18420 22584 18472 22636
rect 22376 22652 22428 22704
rect 23388 22652 23440 22704
rect 24676 22652 24728 22704
rect 28080 22695 28132 22704
rect 18788 22627 18840 22636
rect 18788 22593 18797 22627
rect 18797 22593 18831 22627
rect 18831 22593 18840 22627
rect 19432 22627 19484 22636
rect 18788 22584 18840 22593
rect 19432 22593 19441 22627
rect 19441 22593 19475 22627
rect 19475 22593 19484 22627
rect 19432 22584 19484 22593
rect 19524 22627 19576 22636
rect 19524 22593 19533 22627
rect 19533 22593 19567 22627
rect 19567 22593 19576 22627
rect 19800 22627 19852 22636
rect 19524 22584 19576 22593
rect 19800 22593 19809 22627
rect 19809 22593 19843 22627
rect 19843 22593 19852 22627
rect 19800 22584 19852 22593
rect 20904 22627 20956 22636
rect 20904 22593 20913 22627
rect 20913 22593 20947 22627
rect 20947 22593 20956 22627
rect 20904 22584 20956 22593
rect 21088 22584 21140 22636
rect 22008 22584 22060 22636
rect 24216 22627 24268 22636
rect 24216 22593 24225 22627
rect 24225 22593 24259 22627
rect 24259 22593 24268 22627
rect 24216 22584 24268 22593
rect 24492 22627 24544 22636
rect 24492 22593 24526 22627
rect 24526 22593 24544 22627
rect 24492 22584 24544 22593
rect 25780 22584 25832 22636
rect 27804 22627 27856 22636
rect 27804 22593 27813 22627
rect 27813 22593 27847 22627
rect 27847 22593 27856 22627
rect 27804 22584 27856 22593
rect 28080 22661 28114 22695
rect 28114 22661 28132 22695
rect 28080 22652 28132 22661
rect 28908 22652 28960 22704
rect 30012 22584 30064 22636
rect 30380 22627 30432 22636
rect 30380 22593 30389 22627
rect 30389 22593 30423 22627
rect 30423 22593 30432 22627
rect 30380 22584 30432 22593
rect 30564 22627 30616 22636
rect 30564 22593 30573 22627
rect 30573 22593 30607 22627
rect 30607 22593 30616 22627
rect 30564 22584 30616 22593
rect 19340 22516 19392 22568
rect 19708 22559 19760 22568
rect 19708 22525 19717 22559
rect 19717 22525 19751 22559
rect 19751 22525 19760 22559
rect 19708 22516 19760 22525
rect 20536 22516 20588 22568
rect 15108 22380 15160 22432
rect 15292 22380 15344 22432
rect 15568 22380 15620 22432
rect 17132 22380 17184 22432
rect 17408 22380 17460 22432
rect 18052 22423 18104 22432
rect 18052 22389 18061 22423
rect 18061 22389 18095 22423
rect 18095 22389 18104 22423
rect 18052 22380 18104 22389
rect 18696 22380 18748 22432
rect 18880 22380 18932 22432
rect 19524 22380 19576 22432
rect 19616 22380 19668 22432
rect 23756 22380 23808 22432
rect 25596 22423 25648 22432
rect 25596 22389 25605 22423
rect 25605 22389 25639 22423
rect 25639 22389 25648 22423
rect 25596 22380 25648 22389
rect 30656 22380 30708 22432
rect 2136 22278 2188 22330
rect 12440 22278 12492 22330
rect 22744 22278 22796 22330
rect 1676 22176 1728 22228
rect 3792 22219 3844 22228
rect 3792 22185 3801 22219
rect 3801 22185 3835 22219
rect 3835 22185 3844 22219
rect 3792 22176 3844 22185
rect 3884 22176 3936 22228
rect 4896 22151 4948 22160
rect 4896 22117 4905 22151
rect 4905 22117 4939 22151
rect 4939 22117 4948 22151
rect 4896 22108 4948 22117
rect 5264 22108 5316 22160
rect 5724 22176 5776 22228
rect 7932 22176 7984 22228
rect 9680 22176 9732 22228
rect 9772 22176 9824 22228
rect 12164 22219 12216 22228
rect 1860 21972 1912 22024
rect 2228 21972 2280 22024
rect 2688 21972 2740 22024
rect 3792 21972 3844 22024
rect 5172 22040 5224 22092
rect 9404 22108 9456 22160
rect 4436 22015 4488 22024
rect 4436 21981 4445 22015
rect 4445 21981 4479 22015
rect 4479 21981 4488 22015
rect 4436 21972 4488 21981
rect 4712 21972 4764 22024
rect 5080 22015 5132 22024
rect 5080 21981 5089 22015
rect 5089 21981 5123 22015
rect 5123 21981 5132 22015
rect 5080 21972 5132 21981
rect 5724 21972 5776 22024
rect 9036 22040 9088 22092
rect 6920 21947 6972 21956
rect 6920 21913 6929 21947
rect 6929 21913 6963 21947
rect 6963 21913 6972 21947
rect 6920 21904 6972 21913
rect 7748 21972 7800 22024
rect 8024 21972 8076 22024
rect 8300 21972 8352 22024
rect 8944 21972 8996 22024
rect 12164 22185 12173 22219
rect 12173 22185 12207 22219
rect 12207 22185 12216 22219
rect 12164 22176 12216 22185
rect 11244 22040 11296 22092
rect 12164 22040 12216 22092
rect 12716 22108 12768 22160
rect 13636 22108 13688 22160
rect 14372 22108 14424 22160
rect 14924 22108 14976 22160
rect 15292 22108 15344 22160
rect 15568 22176 15620 22228
rect 15936 22176 15988 22228
rect 17408 22176 17460 22228
rect 18236 22108 18288 22160
rect 19432 22176 19484 22228
rect 22560 22108 22612 22160
rect 27252 22108 27304 22160
rect 12532 22083 12584 22092
rect 12532 22049 12541 22083
rect 12541 22049 12575 22083
rect 12575 22049 12584 22083
rect 12532 22040 12584 22049
rect 12900 22040 12952 22092
rect 10876 21972 10928 22024
rect 3148 21836 3200 21888
rect 4252 21836 4304 21888
rect 6276 21836 6328 21888
rect 7472 21836 7524 21888
rect 7932 21836 7984 21888
rect 8392 21879 8444 21888
rect 8392 21845 8401 21879
rect 8401 21845 8435 21879
rect 8435 21845 8444 21879
rect 8392 21836 8444 21845
rect 10508 21836 10560 21888
rect 10784 21879 10836 21888
rect 10784 21845 10793 21879
rect 10793 21845 10827 21879
rect 10827 21845 10836 21879
rect 10784 21836 10836 21845
rect 10968 21836 11020 21888
rect 12348 22015 12400 22024
rect 12348 21981 12357 22015
rect 12357 21981 12391 22015
rect 12391 21981 12400 22015
rect 12348 21972 12400 21981
rect 13084 21972 13136 22024
rect 13452 22040 13504 22092
rect 16120 22040 16172 22092
rect 17408 22040 17460 22092
rect 12532 21904 12584 21956
rect 13820 21904 13872 21956
rect 14556 21972 14608 22024
rect 15108 22015 15160 22024
rect 15108 21981 15117 22015
rect 15117 21981 15151 22015
rect 15151 21981 15160 22015
rect 15108 21972 15160 21981
rect 15476 21972 15528 22024
rect 15568 22015 15620 22024
rect 15568 21981 15577 22015
rect 15577 21981 15611 22015
rect 15611 21981 15620 22015
rect 15568 21972 15620 21981
rect 14648 21904 14700 21956
rect 15292 21904 15344 21956
rect 16120 21904 16172 21956
rect 17132 21972 17184 22024
rect 18880 22040 18932 22092
rect 19616 22083 19668 22092
rect 19616 22049 19625 22083
rect 19625 22049 19659 22083
rect 19659 22049 19668 22083
rect 19616 22040 19668 22049
rect 20996 22040 21048 22092
rect 18052 21972 18104 22024
rect 19800 21972 19852 22024
rect 11612 21836 11664 21888
rect 14372 21836 14424 21888
rect 15476 21836 15528 21888
rect 18328 21904 18380 21956
rect 20904 21972 20956 22024
rect 22100 21972 22152 22024
rect 22928 22040 22980 22092
rect 27712 22083 27764 22092
rect 22376 21972 22428 22024
rect 21916 21904 21968 21956
rect 17684 21836 17736 21888
rect 18788 21836 18840 21888
rect 19156 21836 19208 21888
rect 20168 21836 20220 21888
rect 20904 21836 20956 21888
rect 21180 21879 21232 21888
rect 21180 21845 21189 21879
rect 21189 21845 21223 21879
rect 21223 21845 21232 21879
rect 21180 21836 21232 21845
rect 22376 21836 22428 21888
rect 22468 21836 22520 21888
rect 22928 21904 22980 21956
rect 23388 21972 23440 22024
rect 23756 22015 23808 22024
rect 23756 21981 23765 22015
rect 23765 21981 23799 22015
rect 23799 21981 23808 22015
rect 23756 21972 23808 21981
rect 24584 22015 24636 22024
rect 24584 21981 24593 22015
rect 24593 21981 24627 22015
rect 24627 21981 24636 22015
rect 24584 21972 24636 21981
rect 27712 22049 27721 22083
rect 27721 22049 27755 22083
rect 27755 22049 27764 22083
rect 27712 22040 27764 22049
rect 28448 22040 28500 22092
rect 24860 22015 24912 22024
rect 24860 21981 24869 22015
rect 24869 21981 24903 22015
rect 24903 21981 24912 22015
rect 24860 21972 24912 21981
rect 25688 21972 25740 22024
rect 26792 21972 26844 22024
rect 29276 21972 29328 22024
rect 29920 22015 29972 22024
rect 29920 21981 29929 22015
rect 29929 21981 29963 22015
rect 29963 21981 29972 22015
rect 29920 21972 29972 21981
rect 25964 21904 26016 21956
rect 30932 21972 30984 22024
rect 30748 21904 30800 21956
rect 24952 21836 25004 21888
rect 30564 21836 30616 21888
rect 7288 21734 7340 21786
rect 17592 21734 17644 21786
rect 27896 21734 27948 21786
rect 1400 21632 1452 21684
rect 2320 21632 2372 21684
rect 5080 21632 5132 21684
rect 6460 21632 6512 21684
rect 10876 21632 10928 21684
rect 3608 21564 3660 21616
rect 3792 21564 3844 21616
rect 2504 21496 2556 21548
rect 4896 21539 4948 21548
rect 4896 21505 4905 21539
rect 4905 21505 4939 21539
rect 4939 21505 4948 21539
rect 4896 21496 4948 21505
rect 2780 21428 2832 21480
rect 4436 21428 4488 21480
rect 5264 21428 5316 21480
rect 6460 21496 6512 21548
rect 7840 21539 7892 21548
rect 7840 21505 7849 21539
rect 7849 21505 7883 21539
rect 7883 21505 7892 21539
rect 7840 21496 7892 21505
rect 8392 21496 8444 21548
rect 9220 21539 9272 21548
rect 9220 21505 9229 21539
rect 9229 21505 9263 21539
rect 9263 21505 9272 21539
rect 9220 21496 9272 21505
rect 6920 21428 6972 21480
rect 8024 21471 8076 21480
rect 8024 21437 8033 21471
rect 8033 21437 8067 21471
rect 8067 21437 8076 21471
rect 13820 21632 13872 21684
rect 14648 21564 14700 21616
rect 15844 21564 15896 21616
rect 16304 21632 16356 21684
rect 16672 21564 16724 21616
rect 16764 21564 16816 21616
rect 9956 21496 10008 21548
rect 10324 21539 10376 21548
rect 10324 21505 10333 21539
rect 10333 21505 10367 21539
rect 10367 21505 10376 21539
rect 10324 21496 10376 21505
rect 10784 21496 10836 21548
rect 11244 21496 11296 21548
rect 11704 21496 11756 21548
rect 12164 21496 12216 21548
rect 12348 21496 12400 21548
rect 13452 21496 13504 21548
rect 14372 21539 14424 21548
rect 14372 21505 14381 21539
rect 14381 21505 14415 21539
rect 14415 21505 14424 21539
rect 14372 21496 14424 21505
rect 14832 21496 14884 21548
rect 15752 21496 15804 21548
rect 19156 21564 19208 21616
rect 19340 21564 19392 21616
rect 20444 21564 20496 21616
rect 20996 21632 21048 21684
rect 22008 21632 22060 21684
rect 22192 21632 22244 21684
rect 23204 21675 23256 21684
rect 23204 21641 23213 21675
rect 23213 21641 23247 21675
rect 23247 21641 23256 21675
rect 23204 21632 23256 21641
rect 24492 21632 24544 21684
rect 25964 21675 26016 21684
rect 25964 21641 25973 21675
rect 25973 21641 26007 21675
rect 26007 21641 26016 21675
rect 25964 21632 26016 21641
rect 26424 21632 26476 21684
rect 27344 21632 27396 21684
rect 21824 21564 21876 21616
rect 8024 21428 8076 21437
rect 14280 21428 14332 21480
rect 14924 21428 14976 21480
rect 15108 21471 15160 21480
rect 15108 21437 15117 21471
rect 15117 21437 15151 21471
rect 15151 21437 15160 21471
rect 15108 21428 15160 21437
rect 6736 21403 6788 21412
rect 1676 21292 1728 21344
rect 2320 21292 2372 21344
rect 3056 21292 3108 21344
rect 6736 21369 6745 21403
rect 6745 21369 6779 21403
rect 6779 21369 6788 21403
rect 6736 21360 6788 21369
rect 9588 21360 9640 21412
rect 10876 21360 10928 21412
rect 12348 21360 12400 21412
rect 14096 21360 14148 21412
rect 15660 21428 15712 21480
rect 4712 21335 4764 21344
rect 4712 21301 4721 21335
rect 4721 21301 4755 21335
rect 4755 21301 4764 21335
rect 4712 21292 4764 21301
rect 4988 21292 5040 21344
rect 11612 21292 11664 21344
rect 12532 21292 12584 21344
rect 12716 21292 12768 21344
rect 14188 21335 14240 21344
rect 14188 21301 14197 21335
rect 14197 21301 14231 21335
rect 14231 21301 14240 21335
rect 14188 21292 14240 21301
rect 15660 21292 15712 21344
rect 18696 21539 18748 21548
rect 18696 21505 18705 21539
rect 18705 21505 18739 21539
rect 18739 21505 18748 21539
rect 18696 21496 18748 21505
rect 18880 21496 18932 21548
rect 19892 21496 19944 21548
rect 22560 21496 22612 21548
rect 24860 21564 24912 21616
rect 24768 21539 24820 21548
rect 24768 21505 24777 21539
rect 24777 21505 24811 21539
rect 24811 21505 24820 21539
rect 24768 21496 24820 21505
rect 26148 21539 26200 21548
rect 26148 21505 26157 21539
rect 26157 21505 26191 21539
rect 26191 21505 26200 21539
rect 26148 21496 26200 21505
rect 26700 21564 26752 21616
rect 27712 21564 27764 21616
rect 27160 21539 27212 21548
rect 27160 21505 27169 21539
rect 27169 21505 27203 21539
rect 27203 21505 27212 21539
rect 27160 21496 27212 21505
rect 27436 21539 27488 21548
rect 27436 21505 27445 21539
rect 27445 21505 27479 21539
rect 27479 21505 27488 21539
rect 27436 21496 27488 21505
rect 27804 21496 27856 21548
rect 28264 21539 28316 21548
rect 28264 21505 28273 21539
rect 28273 21505 28307 21539
rect 28307 21505 28316 21539
rect 28264 21496 28316 21505
rect 16120 21292 16172 21344
rect 16396 21292 16448 21344
rect 19248 21428 19300 21480
rect 23388 21471 23440 21480
rect 23388 21437 23397 21471
rect 23397 21437 23431 21471
rect 23431 21437 23440 21471
rect 23388 21428 23440 21437
rect 25320 21428 25372 21480
rect 25596 21428 25648 21480
rect 27712 21428 27764 21480
rect 28540 21471 28592 21480
rect 28540 21437 28549 21471
rect 28549 21437 28583 21471
rect 28583 21437 28592 21471
rect 28540 21428 28592 21437
rect 31116 21632 31168 21684
rect 29184 21607 29236 21616
rect 29184 21573 29193 21607
rect 29193 21573 29227 21607
rect 29227 21573 29236 21607
rect 29184 21564 29236 21573
rect 29460 21564 29512 21616
rect 30012 21496 30064 21548
rect 30380 21496 30432 21548
rect 30564 21496 30616 21548
rect 30840 21496 30892 21548
rect 30104 21428 30156 21480
rect 17776 21360 17828 21412
rect 20904 21360 20956 21412
rect 24768 21360 24820 21412
rect 27528 21360 27580 21412
rect 28632 21360 28684 21412
rect 18328 21292 18380 21344
rect 18788 21292 18840 21344
rect 22192 21292 22244 21344
rect 22928 21292 22980 21344
rect 25044 21292 25096 21344
rect 26516 21292 26568 21344
rect 27988 21292 28040 21344
rect 28172 21292 28224 21344
rect 28908 21292 28960 21344
rect 30932 21292 30984 21344
rect 2136 21190 2188 21242
rect 12440 21190 12492 21242
rect 22744 21190 22796 21242
rect 2596 21088 2648 21140
rect 2872 21088 2924 21140
rect 3516 21088 3568 21140
rect 5632 21020 5684 21072
rect 5908 21020 5960 21072
rect 8668 21088 8720 21140
rect 9220 21088 9272 21140
rect 10784 21088 10836 21140
rect 11060 21088 11112 21140
rect 9404 21020 9456 21072
rect 9680 21020 9732 21072
rect 7196 20952 7248 21004
rect 12348 21020 12400 21072
rect 12900 21020 12952 21072
rect 2780 20884 2832 20936
rect 5632 20884 5684 20936
rect 6736 20927 6788 20936
rect 1860 20816 1912 20868
rect 4712 20816 4764 20868
rect 5080 20816 5132 20868
rect 6736 20893 6745 20927
rect 6745 20893 6779 20927
rect 6779 20893 6788 20927
rect 6736 20884 6788 20893
rect 6828 20927 6880 20936
rect 6828 20893 6837 20927
rect 6837 20893 6871 20927
rect 6871 20893 6880 20927
rect 6828 20884 6880 20893
rect 7472 20884 7524 20936
rect 7840 20884 7892 20936
rect 8576 20884 8628 20936
rect 9220 20884 9272 20936
rect 10692 20927 10744 20936
rect 7012 20816 7064 20868
rect 7564 20816 7616 20868
rect 9772 20859 9824 20868
rect 9772 20825 9781 20859
rect 9781 20825 9815 20859
rect 9815 20825 9824 20859
rect 9772 20816 9824 20825
rect 9956 20816 10008 20868
rect 10692 20893 10701 20927
rect 10701 20893 10735 20927
rect 10735 20893 10744 20927
rect 10692 20884 10744 20893
rect 12164 20952 12216 21004
rect 12808 20952 12860 21004
rect 18420 21088 18472 21140
rect 20628 21088 20680 21140
rect 20720 21088 20772 21140
rect 21272 21088 21324 21140
rect 24032 21088 24084 21140
rect 26700 21131 26752 21140
rect 26700 21097 26709 21131
rect 26709 21097 26743 21131
rect 26743 21097 26752 21131
rect 26700 21088 26752 21097
rect 27344 21020 27396 21072
rect 28540 21088 28592 21140
rect 30748 21131 30800 21140
rect 30748 21097 30757 21131
rect 30757 21097 30791 21131
rect 30791 21097 30800 21131
rect 30748 21088 30800 21097
rect 11244 20884 11296 20936
rect 11796 20884 11848 20936
rect 12072 20927 12124 20936
rect 12072 20893 12081 20927
rect 12081 20893 12115 20927
rect 12115 20893 12124 20927
rect 12072 20884 12124 20893
rect 12256 20927 12308 20936
rect 12256 20893 12265 20927
rect 12265 20893 12299 20927
rect 12299 20893 12308 20927
rect 12256 20884 12308 20893
rect 12348 20884 12400 20936
rect 12716 20927 12768 20936
rect 12716 20893 12725 20927
rect 12725 20893 12759 20927
rect 12759 20893 12768 20927
rect 12716 20884 12768 20893
rect 14096 20927 14148 20936
rect 14096 20893 14105 20927
rect 14105 20893 14139 20927
rect 14139 20893 14148 20927
rect 14096 20884 14148 20893
rect 14372 20884 14424 20936
rect 15016 20927 15068 20936
rect 15016 20893 15050 20927
rect 15050 20893 15068 20927
rect 15016 20884 15068 20893
rect 5724 20748 5776 20800
rect 8576 20748 8628 20800
rect 10048 20748 10100 20800
rect 11060 20748 11112 20800
rect 11980 20816 12032 20868
rect 15936 20884 15988 20936
rect 17132 20927 17184 20936
rect 17132 20893 17141 20927
rect 17141 20893 17175 20927
rect 17175 20893 17184 20927
rect 17132 20884 17184 20893
rect 15384 20816 15436 20868
rect 15752 20816 15804 20868
rect 16304 20816 16356 20868
rect 17684 20884 17736 20936
rect 17776 20884 17828 20936
rect 18052 20927 18104 20936
rect 18052 20893 18061 20927
rect 18061 20893 18095 20927
rect 18095 20893 18104 20927
rect 18052 20884 18104 20893
rect 18420 20884 18472 20936
rect 18696 20927 18748 20936
rect 18144 20816 18196 20868
rect 18696 20893 18705 20927
rect 18705 20893 18739 20927
rect 18739 20893 18748 20927
rect 18696 20884 18748 20893
rect 19432 20927 19484 20936
rect 19432 20893 19441 20927
rect 19441 20893 19475 20927
rect 19475 20893 19484 20927
rect 19432 20884 19484 20893
rect 21916 20952 21968 21004
rect 22376 20952 22428 21004
rect 23112 20995 23164 21004
rect 23112 20961 23121 20995
rect 23121 20961 23155 20995
rect 23155 20961 23164 20995
rect 23112 20952 23164 20961
rect 20996 20884 21048 20936
rect 21548 20884 21600 20936
rect 22468 20884 22520 20936
rect 26424 20952 26476 21004
rect 27252 20952 27304 21004
rect 28080 21020 28132 21072
rect 28172 21063 28224 21072
rect 28172 21029 28181 21063
rect 28181 21029 28215 21063
rect 28215 21029 28224 21063
rect 28172 21020 28224 21029
rect 24768 20927 24820 20936
rect 24768 20893 24777 20927
rect 24777 20893 24811 20927
rect 24811 20893 24820 20927
rect 24768 20884 24820 20893
rect 24952 20927 25004 20936
rect 24952 20893 24961 20927
rect 24961 20893 24995 20927
rect 24995 20893 25004 20927
rect 24952 20884 25004 20893
rect 26516 20927 26568 20936
rect 26516 20893 26525 20927
rect 26525 20893 26559 20927
rect 26559 20893 26568 20927
rect 26516 20884 26568 20893
rect 27528 20927 27580 20936
rect 27528 20893 27537 20927
rect 27537 20893 27571 20927
rect 27571 20893 27580 20927
rect 27528 20884 27580 20893
rect 27712 20884 27764 20936
rect 28540 20952 28592 21004
rect 18972 20816 19024 20868
rect 19156 20816 19208 20868
rect 19616 20816 19668 20868
rect 20444 20859 20496 20868
rect 20444 20825 20453 20859
rect 20453 20825 20487 20859
rect 20487 20825 20496 20859
rect 20444 20816 20496 20825
rect 12532 20748 12584 20800
rect 13728 20748 13780 20800
rect 14924 20748 14976 20800
rect 16948 20791 17000 20800
rect 16948 20757 16957 20791
rect 16957 20757 16991 20791
rect 16991 20757 17000 20791
rect 16948 20748 17000 20757
rect 17040 20748 17092 20800
rect 17224 20748 17276 20800
rect 17776 20791 17828 20800
rect 17776 20757 17785 20791
rect 17785 20757 17819 20791
rect 17819 20757 17828 20791
rect 17776 20748 17828 20757
rect 17868 20748 17920 20800
rect 19340 20748 19392 20800
rect 20260 20748 20312 20800
rect 22376 20816 22428 20868
rect 20812 20748 20864 20800
rect 21824 20748 21876 20800
rect 25136 20859 25188 20868
rect 25136 20825 25145 20859
rect 25145 20825 25179 20859
rect 25179 20825 25188 20859
rect 25136 20816 25188 20825
rect 27436 20816 27488 20868
rect 28448 20884 28500 20936
rect 28172 20816 28224 20868
rect 26148 20748 26200 20800
rect 27252 20748 27304 20800
rect 29644 20927 29696 20936
rect 29644 20893 29653 20927
rect 29653 20893 29687 20927
rect 29687 20893 29696 20927
rect 29644 20884 29696 20893
rect 31300 20952 31352 21004
rect 30104 20927 30156 20936
rect 30104 20893 30118 20927
rect 30118 20893 30152 20927
rect 30152 20893 30156 20927
rect 30932 20927 30984 20936
rect 30104 20884 30156 20893
rect 30932 20893 30941 20927
rect 30941 20893 30975 20927
rect 30975 20893 30984 20927
rect 30932 20884 30984 20893
rect 29460 20816 29512 20868
rect 30472 20816 30524 20868
rect 31208 20816 31260 20868
rect 7288 20646 7340 20698
rect 17592 20646 17644 20698
rect 27896 20646 27948 20698
rect 1860 20587 1912 20596
rect 1860 20553 1869 20587
rect 1869 20553 1903 20587
rect 1903 20553 1912 20587
rect 1860 20544 1912 20553
rect 2044 20544 2096 20596
rect 5080 20587 5132 20596
rect 1676 20476 1728 20528
rect 2044 20451 2096 20460
rect 2044 20417 2053 20451
rect 2053 20417 2087 20451
rect 2087 20417 2096 20451
rect 2044 20408 2096 20417
rect 2228 20408 2280 20460
rect 2688 20408 2740 20460
rect 2596 20340 2648 20392
rect 3056 20383 3108 20392
rect 3056 20349 3065 20383
rect 3065 20349 3099 20383
rect 3099 20349 3108 20383
rect 3056 20340 3108 20349
rect 2228 20247 2280 20256
rect 2228 20213 2237 20247
rect 2237 20213 2271 20247
rect 2271 20213 2280 20247
rect 2228 20204 2280 20213
rect 5080 20553 5089 20587
rect 5089 20553 5123 20587
rect 5123 20553 5132 20587
rect 5080 20544 5132 20553
rect 6184 20544 6236 20596
rect 6828 20544 6880 20596
rect 4988 20476 5040 20528
rect 6644 20476 6696 20528
rect 4712 20408 4764 20460
rect 5356 20408 5408 20460
rect 6920 20451 6972 20460
rect 4252 20340 4304 20392
rect 6920 20417 6929 20451
rect 6929 20417 6963 20451
rect 6963 20417 6972 20451
rect 6920 20408 6972 20417
rect 7380 20476 7432 20528
rect 8116 20476 8168 20528
rect 8484 20544 8536 20596
rect 9772 20544 9824 20596
rect 10508 20544 10560 20596
rect 10692 20544 10744 20596
rect 5172 20272 5224 20324
rect 8024 20451 8076 20460
rect 8024 20417 8033 20451
rect 8033 20417 8067 20451
rect 8067 20417 8076 20451
rect 8208 20451 8260 20460
rect 8024 20408 8076 20417
rect 8208 20417 8217 20451
rect 8217 20417 8251 20451
rect 8251 20417 8260 20451
rect 8208 20408 8260 20417
rect 9036 20408 9088 20460
rect 9128 20408 9180 20460
rect 11244 20544 11296 20596
rect 11336 20544 11388 20596
rect 17224 20544 17276 20596
rect 11060 20476 11112 20528
rect 9956 20408 10008 20460
rect 7656 20272 7708 20324
rect 10784 20451 10836 20460
rect 10784 20417 10793 20451
rect 10793 20417 10827 20451
rect 10827 20417 10836 20451
rect 10784 20408 10836 20417
rect 11244 20340 11296 20392
rect 11888 20476 11940 20528
rect 14188 20476 14240 20528
rect 14556 20476 14608 20528
rect 15108 20476 15160 20528
rect 15476 20476 15528 20528
rect 16120 20476 16172 20528
rect 16672 20476 16724 20528
rect 16764 20476 16816 20528
rect 11612 20451 11664 20460
rect 11612 20417 11621 20451
rect 11621 20417 11655 20451
rect 11655 20417 11664 20451
rect 11612 20408 11664 20417
rect 11796 20451 11848 20460
rect 11796 20417 11804 20451
rect 11804 20417 11838 20451
rect 11838 20417 11848 20451
rect 11796 20408 11848 20417
rect 12164 20451 12216 20460
rect 12164 20417 12173 20451
rect 12173 20417 12207 20451
rect 12207 20417 12216 20451
rect 12164 20408 12216 20417
rect 12532 20408 12584 20460
rect 14924 20408 14976 20460
rect 15384 20451 15436 20460
rect 15384 20417 15393 20451
rect 15393 20417 15427 20451
rect 15427 20417 15436 20451
rect 15384 20408 15436 20417
rect 15660 20408 15712 20460
rect 16028 20408 16080 20460
rect 8116 20272 8168 20324
rect 5356 20204 5408 20256
rect 6920 20204 6972 20256
rect 7380 20204 7432 20256
rect 8484 20204 8536 20256
rect 9404 20204 9456 20256
rect 11060 20204 11112 20256
rect 11704 20272 11756 20324
rect 12348 20340 12400 20392
rect 12808 20340 12860 20392
rect 14648 20340 14700 20392
rect 16948 20451 17000 20460
rect 16948 20417 16957 20451
rect 16957 20417 16991 20451
rect 16991 20417 17000 20451
rect 18604 20544 18656 20596
rect 18880 20544 18932 20596
rect 23480 20587 23532 20596
rect 18236 20519 18288 20528
rect 18236 20485 18259 20519
rect 18259 20485 18288 20519
rect 18236 20476 18288 20485
rect 19616 20476 19668 20528
rect 20076 20476 20128 20528
rect 16948 20408 17000 20417
rect 16672 20340 16724 20392
rect 18696 20408 18748 20460
rect 18972 20408 19024 20460
rect 19984 20340 20036 20392
rect 20720 20408 20772 20460
rect 21456 20476 21508 20528
rect 23480 20553 23489 20587
rect 23489 20553 23523 20587
rect 23523 20553 23532 20587
rect 23480 20544 23532 20553
rect 24584 20544 24636 20596
rect 27252 20587 27304 20596
rect 27252 20553 27261 20587
rect 27261 20553 27295 20587
rect 27295 20553 27304 20587
rect 27252 20544 27304 20553
rect 27620 20587 27672 20596
rect 27620 20553 27629 20587
rect 27629 20553 27663 20587
rect 27663 20553 27672 20587
rect 27620 20544 27672 20553
rect 27804 20544 27856 20596
rect 29092 20544 29144 20596
rect 29184 20544 29236 20596
rect 29644 20544 29696 20596
rect 31116 20544 31168 20596
rect 21824 20408 21876 20460
rect 22928 20408 22980 20460
rect 12164 20272 12216 20324
rect 15568 20272 15620 20324
rect 16028 20272 16080 20324
rect 16304 20272 16356 20324
rect 20996 20340 21048 20392
rect 21732 20340 21784 20392
rect 23756 20408 23808 20460
rect 24768 20408 24820 20460
rect 24860 20408 24912 20460
rect 26976 20408 27028 20460
rect 24216 20340 24268 20392
rect 25412 20340 25464 20392
rect 25596 20340 25648 20392
rect 27712 20340 27764 20392
rect 29736 20408 29788 20460
rect 30564 20476 30616 20528
rect 12348 20204 12400 20256
rect 14740 20204 14792 20256
rect 15476 20204 15528 20256
rect 16856 20204 16908 20256
rect 20260 20272 20312 20324
rect 21916 20272 21968 20324
rect 22560 20272 22612 20324
rect 23020 20272 23072 20324
rect 24860 20272 24912 20324
rect 27620 20272 27672 20324
rect 28448 20272 28500 20324
rect 29092 20272 29144 20324
rect 29368 20340 29420 20392
rect 30840 20340 30892 20392
rect 30196 20272 30248 20324
rect 20076 20204 20128 20256
rect 20628 20204 20680 20256
rect 22008 20204 22060 20256
rect 22284 20204 22336 20256
rect 22468 20204 22520 20256
rect 23388 20204 23440 20256
rect 24308 20204 24360 20256
rect 24676 20204 24728 20256
rect 25136 20204 25188 20256
rect 26056 20204 26108 20256
rect 26332 20247 26384 20256
rect 26332 20213 26341 20247
rect 26341 20213 26375 20247
rect 26375 20213 26384 20247
rect 26332 20204 26384 20213
rect 28816 20247 28868 20256
rect 28816 20213 28825 20247
rect 28825 20213 28859 20247
rect 28859 20213 28868 20247
rect 28816 20204 28868 20213
rect 29460 20204 29512 20256
rect 30288 20204 30340 20256
rect 30748 20247 30800 20256
rect 30748 20213 30757 20247
rect 30757 20213 30791 20247
rect 30791 20213 30800 20247
rect 30748 20204 30800 20213
rect 30840 20204 30892 20256
rect 31208 20204 31260 20256
rect 2136 20102 2188 20154
rect 12440 20102 12492 20154
rect 22744 20102 22796 20154
rect 2044 20000 2096 20052
rect 5172 20043 5224 20052
rect 5172 20009 5181 20043
rect 5181 20009 5215 20043
rect 5215 20009 5224 20043
rect 5172 20000 5224 20009
rect 6000 20000 6052 20052
rect 6368 20000 6420 20052
rect 7012 20043 7064 20052
rect 7012 20009 7021 20043
rect 7021 20009 7055 20043
rect 7055 20009 7064 20043
rect 7012 20000 7064 20009
rect 8760 20000 8812 20052
rect 8852 20000 8904 20052
rect 8668 19932 8720 19984
rect 9312 19932 9364 19984
rect 1308 19796 1360 19848
rect 3516 19864 3568 19916
rect 5632 19907 5684 19916
rect 5632 19873 5641 19907
rect 5641 19873 5675 19907
rect 5675 19873 5684 19907
rect 5632 19864 5684 19873
rect 8392 19864 8444 19916
rect 10692 19932 10744 19984
rect 11980 19932 12032 19984
rect 15660 20000 15712 20052
rect 1124 19728 1176 19780
rect 1676 19728 1728 19780
rect 1584 19660 1636 19712
rect 2872 19796 2924 19848
rect 3884 19796 3936 19848
rect 3056 19728 3108 19780
rect 6368 19728 6420 19780
rect 10416 19864 10468 19916
rect 9128 19796 9180 19848
rect 9956 19839 10008 19848
rect 9956 19805 9965 19839
rect 9965 19805 9999 19839
rect 9999 19805 10008 19839
rect 9956 19796 10008 19805
rect 10508 19839 10560 19848
rect 3608 19660 3660 19712
rect 4344 19660 4396 19712
rect 9772 19728 9824 19780
rect 10508 19805 10517 19839
rect 10517 19805 10551 19839
rect 10551 19805 10560 19839
rect 10508 19796 10560 19805
rect 10140 19728 10192 19780
rect 14280 19932 14332 19984
rect 18052 20000 18104 20052
rect 18236 20000 18288 20052
rect 19984 20000 20036 20052
rect 21272 20000 21324 20052
rect 21640 20000 21692 20052
rect 22284 20000 22336 20052
rect 18328 19932 18380 19984
rect 18604 19932 18656 19984
rect 19248 19932 19300 19984
rect 21916 19932 21968 19984
rect 23480 20000 23532 20052
rect 24768 20043 24820 20052
rect 24768 20009 24777 20043
rect 24777 20009 24811 20043
rect 24811 20009 24820 20043
rect 24768 20000 24820 20009
rect 26240 20000 26292 20052
rect 11244 19839 11296 19848
rect 11244 19805 11253 19839
rect 11253 19805 11287 19839
rect 11287 19805 11296 19839
rect 11244 19796 11296 19805
rect 11520 19796 11572 19848
rect 11060 19728 11112 19780
rect 12348 19796 12400 19848
rect 14188 19864 14240 19916
rect 13084 19839 13136 19848
rect 13084 19805 13093 19839
rect 13093 19805 13127 19839
rect 13127 19805 13136 19839
rect 13084 19796 13136 19805
rect 11980 19728 12032 19780
rect 7656 19660 7708 19712
rect 8116 19703 8168 19712
rect 8116 19669 8125 19703
rect 8125 19669 8159 19703
rect 8159 19669 8168 19703
rect 8116 19660 8168 19669
rect 8576 19660 8628 19712
rect 12072 19660 12124 19712
rect 12992 19728 13044 19780
rect 14004 19796 14056 19848
rect 14372 19796 14424 19848
rect 14464 19796 14516 19848
rect 14924 19796 14976 19848
rect 15292 19796 15344 19848
rect 15476 19839 15528 19848
rect 15476 19805 15485 19839
rect 15485 19805 15519 19839
rect 15519 19805 15528 19839
rect 15476 19796 15528 19805
rect 16028 19864 16080 19916
rect 16856 19907 16908 19916
rect 16856 19873 16865 19907
rect 16865 19873 16899 19907
rect 16899 19873 16908 19907
rect 16856 19864 16908 19873
rect 17224 19907 17276 19916
rect 17224 19873 17233 19907
rect 17233 19873 17267 19907
rect 17267 19873 17276 19907
rect 17224 19864 17276 19873
rect 17500 19864 17552 19916
rect 18052 19864 18104 19916
rect 18880 19864 18932 19916
rect 18972 19864 19024 19916
rect 19156 19864 19208 19916
rect 17776 19796 17828 19848
rect 17868 19796 17920 19848
rect 14096 19728 14148 19780
rect 14188 19660 14240 19712
rect 15108 19728 15160 19780
rect 19984 19796 20036 19848
rect 20352 19796 20404 19848
rect 14740 19660 14792 19712
rect 15568 19703 15620 19712
rect 15568 19669 15577 19703
rect 15577 19669 15611 19703
rect 15611 19669 15620 19703
rect 15568 19660 15620 19669
rect 20076 19728 20128 19780
rect 20628 19728 20680 19780
rect 22008 19796 22060 19848
rect 25228 19932 25280 19984
rect 27804 20000 27856 20052
rect 28264 20000 28316 20052
rect 27436 19932 27488 19984
rect 27528 19932 27580 19984
rect 24860 19864 24912 19916
rect 27620 19864 27672 19916
rect 29460 20000 29512 20052
rect 29552 20000 29604 20052
rect 30564 20000 30616 20052
rect 25780 19796 25832 19848
rect 26148 19839 26200 19848
rect 26148 19805 26182 19839
rect 26182 19805 26200 19839
rect 26148 19796 26200 19805
rect 22100 19728 22152 19780
rect 18604 19660 18656 19712
rect 24676 19728 24728 19780
rect 25136 19728 25188 19780
rect 28724 19796 28776 19848
rect 28908 19932 28960 19984
rect 29920 19907 29972 19916
rect 29920 19873 29929 19907
rect 29929 19873 29963 19907
rect 29963 19873 29972 19907
rect 29920 19864 29972 19873
rect 28908 19839 28960 19848
rect 28908 19805 28917 19839
rect 28917 19805 28951 19839
rect 28951 19805 28960 19839
rect 28908 19796 28960 19805
rect 30748 19796 30800 19848
rect 27804 19728 27856 19780
rect 28356 19728 28408 19780
rect 30380 19728 30432 19780
rect 31208 19728 31260 19780
rect 23480 19660 23532 19712
rect 28172 19660 28224 19712
rect 29368 19660 29420 19712
rect 29828 19660 29880 19712
rect 30564 19660 30616 19712
rect 31116 19660 31168 19712
rect 7288 19558 7340 19610
rect 17592 19558 17644 19610
rect 27896 19558 27948 19610
rect 2780 19456 2832 19508
rect 3884 19456 3936 19508
rect 4344 19499 4396 19508
rect 4344 19465 4353 19499
rect 4353 19465 4387 19499
rect 4387 19465 4396 19499
rect 4344 19456 4396 19465
rect 6092 19456 6144 19508
rect 6828 19456 6880 19508
rect 7012 19499 7064 19508
rect 7012 19465 7021 19499
rect 7021 19465 7055 19499
rect 7055 19465 7064 19499
rect 7012 19456 7064 19465
rect 8208 19456 8260 19508
rect 8760 19456 8812 19508
rect 1584 19388 1636 19440
rect 1860 19388 1912 19440
rect 1676 19363 1728 19372
rect 1676 19329 1710 19363
rect 1710 19329 1728 19363
rect 1676 19320 1728 19329
rect 1952 19320 2004 19372
rect 2688 19320 2740 19372
rect 3516 19320 3568 19372
rect 3792 19320 3844 19372
rect 7564 19388 7616 19440
rect 5172 19320 5224 19372
rect 3976 19252 4028 19304
rect 4436 19252 4488 19304
rect 5632 19320 5684 19372
rect 8944 19388 8996 19440
rect 6644 19295 6696 19304
rect 6644 19261 6653 19295
rect 6653 19261 6687 19295
rect 6687 19261 6696 19295
rect 6644 19252 6696 19261
rect 8760 19320 8812 19372
rect 9956 19320 10008 19372
rect 10784 19388 10836 19440
rect 11980 19456 12032 19508
rect 12900 19499 12952 19508
rect 12900 19465 12909 19499
rect 12909 19465 12943 19499
rect 12943 19465 12952 19499
rect 12900 19456 12952 19465
rect 13084 19456 13136 19508
rect 14832 19456 14884 19508
rect 15568 19456 15620 19508
rect 15752 19499 15804 19508
rect 15752 19465 15761 19499
rect 15761 19465 15795 19499
rect 15795 19465 15804 19499
rect 15752 19456 15804 19465
rect 16488 19499 16540 19508
rect 16488 19465 16497 19499
rect 16497 19465 16531 19499
rect 16531 19465 16540 19499
rect 16488 19456 16540 19465
rect 16948 19456 17000 19508
rect 18328 19456 18380 19508
rect 19616 19456 19668 19508
rect 21824 19499 21876 19508
rect 21824 19465 21833 19499
rect 21833 19465 21867 19499
rect 21867 19465 21876 19499
rect 21824 19456 21876 19465
rect 11612 19388 11664 19440
rect 12072 19388 12124 19440
rect 6460 19184 6512 19236
rect 11336 19320 11388 19372
rect 11520 19363 11572 19372
rect 11520 19329 11529 19363
rect 11529 19329 11563 19363
rect 11563 19329 11572 19363
rect 11520 19320 11572 19329
rect 12624 19320 12676 19372
rect 13084 19320 13136 19372
rect 13728 19363 13780 19372
rect 13728 19329 13737 19363
rect 13737 19329 13771 19363
rect 13771 19329 13780 19363
rect 13728 19320 13780 19329
rect 14464 19363 14516 19372
rect 14464 19329 14473 19363
rect 14473 19329 14507 19363
rect 14507 19329 14516 19363
rect 14464 19320 14516 19329
rect 1308 19116 1360 19168
rect 2596 19116 2648 19168
rect 2964 19116 3016 19168
rect 4620 19116 4672 19168
rect 10600 19184 10652 19236
rect 11244 19184 11296 19236
rect 13360 19252 13412 19304
rect 14648 19252 14700 19304
rect 15384 19320 15436 19372
rect 16488 19320 16540 19372
rect 16672 19363 16724 19372
rect 16672 19329 16681 19363
rect 16681 19329 16715 19363
rect 16715 19329 16724 19363
rect 16672 19320 16724 19329
rect 15292 19252 15344 19304
rect 17132 19320 17184 19372
rect 18144 19388 18196 19440
rect 18512 19388 18564 19440
rect 23296 19456 23348 19508
rect 18420 19320 18472 19372
rect 23388 19388 23440 19440
rect 9036 19159 9088 19168
rect 9036 19125 9045 19159
rect 9045 19125 9079 19159
rect 9079 19125 9088 19159
rect 9036 19116 9088 19125
rect 9220 19116 9272 19168
rect 11060 19116 11112 19168
rect 11704 19116 11756 19168
rect 15016 19184 15068 19236
rect 13636 19116 13688 19168
rect 18420 19227 18472 19236
rect 18420 19193 18429 19227
rect 18429 19193 18463 19227
rect 18463 19193 18472 19227
rect 18420 19184 18472 19193
rect 18512 19184 18564 19236
rect 19156 19363 19208 19372
rect 19156 19329 19165 19363
rect 19165 19329 19199 19363
rect 19199 19329 19208 19363
rect 19156 19320 19208 19329
rect 19432 19320 19484 19372
rect 20352 19320 20404 19372
rect 19524 19295 19576 19304
rect 19524 19261 19533 19295
rect 19533 19261 19567 19295
rect 19567 19261 19576 19295
rect 19524 19252 19576 19261
rect 20168 19252 20220 19304
rect 21180 19363 21232 19372
rect 21180 19329 21189 19363
rect 21189 19329 21223 19363
rect 21223 19329 21232 19363
rect 21180 19320 21232 19329
rect 22100 19320 22152 19372
rect 21548 19252 21600 19304
rect 22560 19252 22612 19304
rect 23388 19295 23440 19304
rect 23388 19261 23397 19295
rect 23397 19261 23431 19295
rect 23431 19261 23440 19295
rect 23388 19252 23440 19261
rect 25044 19456 25096 19508
rect 25596 19499 25648 19508
rect 25596 19465 25605 19499
rect 25605 19465 25639 19499
rect 25639 19465 25648 19499
rect 25596 19456 25648 19465
rect 25688 19456 25740 19508
rect 25780 19388 25832 19440
rect 24308 19320 24360 19372
rect 24952 19320 25004 19372
rect 28356 19456 28408 19508
rect 28540 19499 28592 19508
rect 28540 19465 28549 19499
rect 28549 19465 28583 19499
rect 28583 19465 28592 19499
rect 28540 19456 28592 19465
rect 29552 19456 29604 19508
rect 29184 19388 29236 19440
rect 28448 19320 28500 19372
rect 18880 19184 18932 19236
rect 23848 19252 23900 19304
rect 25872 19252 25924 19304
rect 27344 19252 27396 19304
rect 28632 19252 28684 19304
rect 29368 19320 29420 19372
rect 30472 19388 30524 19440
rect 29828 19329 29833 19346
rect 29833 19329 29867 19346
rect 29867 19329 29880 19346
rect 29828 19294 29880 19329
rect 30104 19320 30156 19372
rect 30288 19320 30340 19372
rect 31024 19363 31076 19372
rect 15568 19116 15620 19168
rect 17040 19159 17092 19168
rect 17040 19125 17049 19159
rect 17049 19125 17083 19159
rect 17083 19125 17092 19159
rect 17040 19116 17092 19125
rect 17224 19116 17276 19168
rect 17960 19116 18012 19168
rect 21824 19116 21876 19168
rect 22008 19116 22060 19168
rect 28908 19184 28960 19236
rect 31024 19329 31033 19363
rect 31033 19329 31067 19363
rect 31067 19329 31076 19363
rect 31024 19320 31076 19329
rect 31300 19184 31352 19236
rect 26148 19159 26200 19168
rect 26148 19125 26157 19159
rect 26157 19125 26191 19159
rect 26191 19125 26200 19159
rect 26148 19116 26200 19125
rect 27252 19159 27304 19168
rect 27252 19125 27261 19159
rect 27261 19125 27295 19159
rect 27295 19125 27304 19159
rect 27252 19116 27304 19125
rect 28080 19116 28132 19168
rect 2136 19014 2188 19066
rect 12440 19014 12492 19066
rect 22744 19014 22796 19066
rect 5448 18912 5500 18964
rect 6644 18955 6696 18964
rect 6644 18921 6653 18955
rect 6653 18921 6687 18955
rect 6687 18921 6696 18955
rect 6644 18912 6696 18921
rect 10508 18912 10560 18964
rect 10600 18912 10652 18964
rect 13912 18912 13964 18964
rect 21180 18955 21232 18964
rect 1952 18776 2004 18828
rect 3976 18776 4028 18828
rect 1952 18572 2004 18624
rect 2596 18640 2648 18692
rect 4712 18708 4764 18760
rect 4896 18708 4948 18760
rect 2872 18640 2924 18692
rect 5172 18640 5224 18692
rect 7196 18844 7248 18896
rect 8576 18844 8628 18896
rect 7012 18776 7064 18828
rect 8668 18776 8720 18828
rect 8024 18708 8076 18760
rect 8760 18708 8812 18760
rect 7564 18640 7616 18692
rect 9036 18640 9088 18692
rect 9956 18844 10008 18896
rect 9404 18776 9456 18828
rect 9312 18708 9364 18760
rect 9680 18708 9732 18760
rect 10600 18776 10652 18828
rect 11060 18708 11112 18760
rect 11428 18776 11480 18828
rect 11704 18776 11756 18828
rect 11336 18708 11388 18760
rect 12256 18844 12308 18896
rect 12624 18844 12676 18896
rect 12808 18844 12860 18896
rect 16672 18776 16724 18828
rect 18972 18844 19024 18896
rect 21180 18921 21189 18955
rect 21189 18921 21223 18955
rect 21223 18921 21232 18955
rect 21180 18912 21232 18921
rect 22192 18912 22244 18964
rect 23020 18912 23072 18964
rect 23848 18955 23900 18964
rect 23848 18921 23857 18955
rect 23857 18921 23891 18955
rect 23891 18921 23900 18955
rect 23848 18912 23900 18921
rect 24492 18912 24544 18964
rect 25688 18912 25740 18964
rect 27344 18844 27396 18896
rect 28908 18887 28960 18896
rect 18236 18819 18288 18828
rect 18236 18785 18245 18819
rect 18245 18785 18279 18819
rect 18279 18785 18288 18819
rect 18236 18776 18288 18785
rect 18512 18776 18564 18828
rect 13176 18751 13228 18760
rect 13176 18717 13185 18751
rect 13185 18717 13219 18751
rect 13219 18717 13228 18751
rect 13176 18708 13228 18717
rect 13452 18708 13504 18760
rect 14188 18708 14240 18760
rect 15108 18708 15160 18760
rect 15384 18708 15436 18760
rect 16764 18708 16816 18760
rect 17224 18708 17276 18760
rect 10140 18683 10192 18692
rect 10140 18649 10149 18683
rect 10149 18649 10183 18683
rect 10183 18649 10192 18683
rect 10140 18640 10192 18649
rect 5448 18572 5500 18624
rect 6000 18572 6052 18624
rect 6460 18572 6512 18624
rect 6736 18572 6788 18624
rect 7748 18572 7800 18624
rect 10784 18572 10836 18624
rect 10968 18572 11020 18624
rect 12164 18572 12216 18624
rect 12900 18640 12952 18692
rect 15936 18640 15988 18692
rect 17040 18640 17092 18692
rect 18328 18708 18380 18760
rect 18788 18776 18840 18828
rect 19248 18776 19300 18828
rect 20996 18776 21048 18828
rect 23756 18776 23808 18828
rect 28908 18853 28917 18887
rect 28917 18853 28951 18887
rect 28951 18853 28960 18887
rect 28908 18844 28960 18853
rect 30196 18887 30248 18896
rect 30196 18853 30205 18887
rect 30205 18853 30239 18887
rect 30239 18853 30248 18887
rect 30196 18844 30248 18853
rect 17684 18640 17736 18692
rect 20904 18708 20956 18760
rect 21732 18708 21784 18760
rect 23296 18708 23348 18760
rect 24032 18708 24084 18760
rect 24584 18708 24636 18760
rect 25780 18751 25832 18760
rect 25780 18717 25789 18751
rect 25789 18717 25823 18751
rect 25823 18717 25832 18751
rect 25780 18708 25832 18717
rect 26056 18751 26108 18760
rect 26056 18717 26090 18751
rect 26090 18717 26108 18751
rect 26056 18708 26108 18717
rect 28080 18751 28132 18760
rect 28080 18717 28089 18751
rect 28089 18717 28123 18751
rect 28123 18717 28132 18751
rect 28080 18708 28132 18717
rect 28540 18708 28592 18760
rect 13360 18615 13412 18624
rect 13360 18581 13369 18615
rect 13369 18581 13403 18615
rect 13403 18581 13412 18615
rect 13360 18572 13412 18581
rect 13820 18572 13872 18624
rect 17224 18572 17276 18624
rect 19524 18640 19576 18692
rect 21640 18640 21692 18692
rect 24676 18640 24728 18692
rect 27988 18683 28040 18692
rect 27988 18649 27997 18683
rect 27997 18649 28031 18683
rect 28031 18649 28040 18683
rect 27988 18640 28040 18649
rect 28632 18640 28684 18692
rect 30196 18640 30248 18692
rect 30472 18708 30524 18760
rect 30656 18751 30708 18760
rect 30656 18717 30665 18751
rect 30665 18717 30699 18751
rect 30699 18717 30708 18751
rect 30656 18708 30708 18717
rect 31116 18708 31168 18760
rect 30748 18640 30800 18692
rect 17960 18572 18012 18624
rect 19340 18572 19392 18624
rect 20720 18572 20772 18624
rect 22376 18572 22428 18624
rect 23020 18572 23072 18624
rect 23848 18572 23900 18624
rect 24124 18572 24176 18624
rect 24492 18572 24544 18624
rect 27068 18572 27120 18624
rect 27528 18572 27580 18624
rect 28816 18572 28868 18624
rect 29000 18572 29052 18624
rect 30840 18572 30892 18624
rect 7288 18470 7340 18522
rect 17592 18470 17644 18522
rect 27896 18470 27948 18522
rect 1676 18368 1728 18420
rect 6092 18368 6144 18420
rect 6368 18411 6420 18420
rect 6368 18377 6377 18411
rect 6377 18377 6411 18411
rect 6411 18377 6420 18411
rect 6368 18368 6420 18377
rect 7196 18368 7248 18420
rect 7472 18411 7524 18420
rect 7472 18377 7481 18411
rect 7481 18377 7515 18411
rect 7515 18377 7524 18411
rect 7472 18368 7524 18377
rect 7564 18368 7616 18420
rect 14464 18368 14516 18420
rect 15016 18368 15068 18420
rect 1952 18275 2004 18284
rect 1952 18241 1961 18275
rect 1961 18241 1995 18275
rect 1995 18241 2004 18275
rect 1952 18232 2004 18241
rect 2228 18300 2280 18352
rect 2688 18164 2740 18216
rect 3792 18300 3844 18352
rect 4160 18343 4212 18352
rect 4160 18309 4194 18343
rect 4194 18309 4212 18343
rect 4160 18300 4212 18309
rect 5448 18300 5500 18352
rect 2964 18275 3016 18284
rect 2964 18241 2973 18275
rect 2973 18241 3007 18275
rect 3007 18241 3016 18275
rect 2964 18232 3016 18241
rect 3148 18275 3200 18284
rect 3148 18241 3157 18275
rect 3157 18241 3191 18275
rect 3191 18241 3200 18275
rect 3148 18232 3200 18241
rect 3884 18207 3936 18216
rect 3884 18173 3893 18207
rect 3893 18173 3927 18207
rect 3927 18173 3936 18207
rect 3884 18164 3936 18173
rect 4896 18164 4948 18216
rect 7104 18300 7156 18352
rect 8760 18300 8812 18352
rect 7656 18275 7708 18284
rect 7656 18241 7665 18275
rect 7665 18241 7699 18275
rect 7699 18241 7708 18275
rect 7656 18232 7708 18241
rect 7748 18275 7800 18284
rect 7748 18241 7757 18275
rect 7757 18241 7791 18275
rect 7791 18241 7800 18275
rect 7932 18275 7984 18284
rect 7748 18232 7800 18241
rect 7932 18241 7941 18275
rect 7941 18241 7975 18275
rect 7975 18241 7984 18275
rect 7932 18232 7984 18241
rect 8024 18275 8076 18284
rect 8024 18241 8033 18275
rect 8033 18241 8067 18275
rect 8067 18241 8076 18275
rect 9036 18300 9088 18352
rect 13636 18300 13688 18352
rect 8024 18232 8076 18241
rect 9312 18232 9364 18284
rect 10416 18275 10468 18284
rect 10416 18241 10425 18275
rect 10425 18241 10459 18275
rect 10459 18241 10468 18275
rect 10416 18232 10468 18241
rect 10876 18275 10928 18284
rect 3148 18096 3200 18148
rect 6644 18096 6696 18148
rect 9220 18164 9272 18216
rect 9588 18164 9640 18216
rect 10048 18164 10100 18216
rect 10600 18164 10652 18216
rect 10876 18241 10885 18275
rect 10885 18241 10919 18275
rect 10919 18241 10928 18275
rect 10876 18232 10928 18241
rect 11704 18232 11756 18284
rect 11888 18232 11940 18284
rect 12256 18232 12308 18284
rect 12532 18232 12584 18284
rect 13176 18232 13228 18284
rect 13820 18300 13872 18352
rect 17408 18368 17460 18420
rect 17776 18368 17828 18420
rect 17960 18368 18012 18420
rect 18236 18368 18288 18420
rect 18328 18368 18380 18420
rect 19248 18368 19300 18420
rect 19524 18411 19576 18420
rect 19524 18377 19533 18411
rect 19533 18377 19567 18411
rect 19567 18377 19576 18411
rect 19524 18368 19576 18377
rect 22008 18411 22060 18420
rect 22008 18377 22017 18411
rect 22017 18377 22051 18411
rect 22051 18377 22060 18411
rect 22008 18368 22060 18377
rect 22100 18368 22152 18420
rect 22376 18368 22428 18420
rect 23388 18368 23440 18420
rect 24216 18368 24268 18420
rect 26148 18368 26200 18420
rect 26976 18411 27028 18420
rect 26976 18377 26985 18411
rect 26985 18377 27019 18411
rect 27019 18377 27028 18411
rect 26976 18368 27028 18377
rect 27712 18368 27764 18420
rect 28448 18368 28500 18420
rect 16028 18275 16080 18284
rect 2228 18028 2280 18080
rect 5080 18028 5132 18080
rect 5908 18028 5960 18080
rect 9220 18028 9272 18080
rect 10048 18028 10100 18080
rect 10324 18096 10376 18148
rect 10968 18096 11020 18148
rect 11060 18096 11112 18148
rect 12164 18164 12216 18216
rect 12808 18096 12860 18148
rect 14832 18164 14884 18216
rect 16028 18241 16037 18275
rect 16037 18241 16071 18275
rect 16071 18241 16080 18275
rect 16028 18232 16080 18241
rect 18604 18300 18656 18352
rect 16764 18232 16816 18284
rect 17408 18232 17460 18284
rect 15936 18207 15988 18216
rect 15936 18173 15945 18207
rect 15945 18173 15979 18207
rect 15979 18173 15988 18207
rect 15936 18164 15988 18173
rect 17960 18232 18012 18284
rect 18144 18232 18196 18284
rect 18420 18232 18472 18284
rect 20260 18300 20312 18352
rect 21824 18343 21876 18352
rect 21824 18309 21833 18343
rect 21833 18309 21867 18343
rect 21867 18309 21876 18343
rect 21824 18300 21876 18309
rect 19340 18232 19392 18284
rect 12164 18028 12216 18080
rect 12348 18028 12400 18080
rect 12900 18028 12952 18080
rect 15476 18028 15528 18080
rect 15844 18028 15896 18080
rect 16028 18028 16080 18080
rect 17868 18096 17920 18148
rect 18328 18096 18380 18148
rect 20260 18164 20312 18216
rect 20352 18164 20404 18216
rect 20996 18232 21048 18284
rect 21180 18232 21232 18284
rect 21364 18232 21416 18284
rect 24124 18300 24176 18352
rect 24492 18300 24544 18352
rect 25136 18300 25188 18352
rect 27068 18300 27120 18352
rect 22100 18275 22152 18284
rect 22100 18241 22109 18275
rect 22109 18241 22143 18275
rect 22143 18241 22152 18275
rect 22100 18232 22152 18241
rect 23112 18232 23164 18284
rect 23756 18232 23808 18284
rect 25872 18232 25924 18284
rect 27344 18232 27396 18284
rect 27528 18232 27580 18284
rect 29184 18368 29236 18420
rect 29000 18232 29052 18284
rect 29092 18275 29144 18284
rect 29092 18241 29101 18275
rect 29101 18241 29135 18275
rect 29135 18241 29144 18275
rect 30012 18411 30064 18420
rect 30012 18377 30021 18411
rect 30021 18377 30055 18411
rect 30055 18377 30064 18411
rect 30012 18368 30064 18377
rect 29092 18232 29144 18241
rect 21916 18164 21968 18216
rect 18880 18028 18932 18080
rect 19248 18028 19300 18080
rect 19340 18028 19392 18080
rect 19800 18028 19852 18080
rect 20168 18028 20220 18080
rect 21640 18028 21692 18080
rect 21824 18071 21876 18080
rect 21824 18037 21833 18071
rect 21833 18037 21867 18071
rect 21867 18037 21876 18071
rect 21824 18028 21876 18037
rect 24032 18096 24084 18148
rect 24492 18096 24544 18148
rect 22560 18028 22612 18080
rect 23204 18028 23256 18080
rect 28172 18164 28224 18216
rect 28540 18164 28592 18216
rect 29184 18164 29236 18216
rect 30187 18275 30239 18284
rect 30187 18241 30205 18275
rect 30205 18241 30239 18275
rect 30840 18275 30892 18284
rect 30187 18232 30239 18241
rect 30840 18241 30849 18275
rect 30849 18241 30883 18275
rect 30883 18241 30892 18275
rect 30840 18232 30892 18241
rect 31300 18275 31352 18284
rect 30472 18164 30524 18216
rect 31300 18241 31309 18275
rect 31309 18241 31343 18275
rect 31343 18241 31352 18275
rect 31300 18232 31352 18241
rect 31024 18096 31076 18148
rect 25504 18028 25556 18080
rect 26148 18028 26200 18080
rect 27804 18028 27856 18080
rect 30748 18028 30800 18080
rect 2136 17926 2188 17978
rect 12440 17926 12492 17978
rect 22744 17926 22796 17978
rect 3056 17824 3108 17876
rect 3148 17867 3200 17876
rect 3148 17833 3157 17867
rect 3157 17833 3191 17867
rect 3191 17833 3200 17867
rect 3148 17824 3200 17833
rect 4068 17824 4120 17876
rect 4988 17824 5040 17876
rect 5540 17824 5592 17876
rect 6828 17824 6880 17876
rect 7380 17824 7432 17876
rect 7656 17824 7708 17876
rect 10140 17824 10192 17876
rect 14188 17824 14240 17876
rect 940 17756 992 17808
rect 4620 17756 4672 17808
rect 8208 17756 8260 17808
rect 2688 17688 2740 17740
rect 3056 17688 3108 17740
rect 5632 17688 5684 17740
rect 8392 17688 8444 17740
rect 10048 17756 10100 17808
rect 10784 17756 10836 17808
rect 11520 17756 11572 17808
rect 11244 17688 11296 17740
rect 12624 17756 12676 17808
rect 12992 17756 13044 17808
rect 17224 17756 17276 17808
rect 17500 17756 17552 17808
rect 17960 17756 18012 17808
rect 2872 17620 2924 17672
rect 1492 17552 1544 17604
rect 3608 17620 3660 17672
rect 4068 17620 4120 17672
rect 4436 17663 4488 17672
rect 4436 17629 4445 17663
rect 4445 17629 4479 17663
rect 4479 17629 4488 17663
rect 4436 17620 4488 17629
rect 6552 17620 6604 17672
rect 8208 17620 8260 17672
rect 10416 17620 10468 17672
rect 11520 17620 11572 17672
rect 11980 17663 12032 17672
rect 2044 17484 2096 17536
rect 5080 17595 5132 17604
rect 5080 17561 5089 17595
rect 5089 17561 5123 17595
rect 5123 17561 5132 17595
rect 5080 17552 5132 17561
rect 6920 17552 6972 17604
rect 2872 17484 2924 17536
rect 3516 17484 3568 17536
rect 11980 17629 11989 17663
rect 11989 17629 12023 17663
rect 12023 17629 12032 17663
rect 11980 17620 12032 17629
rect 13360 17688 13412 17740
rect 17868 17688 17920 17740
rect 18972 17824 19024 17876
rect 19800 17756 19852 17808
rect 20996 17824 21048 17876
rect 21732 17824 21784 17876
rect 23756 17867 23808 17876
rect 23756 17833 23765 17867
rect 23765 17833 23799 17867
rect 23799 17833 23808 17867
rect 23756 17824 23808 17833
rect 24124 17824 24176 17876
rect 25596 17824 25648 17876
rect 25964 17824 26016 17876
rect 26148 17824 26200 17876
rect 27344 17824 27396 17876
rect 27436 17824 27488 17876
rect 30564 17824 30616 17876
rect 23480 17756 23532 17808
rect 23020 17731 23072 17740
rect 23020 17697 23029 17731
rect 23029 17697 23063 17731
rect 23063 17697 23072 17731
rect 23020 17688 23072 17697
rect 13912 17620 13964 17672
rect 14464 17620 14516 17672
rect 15016 17663 15068 17672
rect 15016 17629 15025 17663
rect 15025 17629 15059 17663
rect 15059 17629 15068 17663
rect 15016 17620 15068 17629
rect 15476 17663 15528 17672
rect 7196 17484 7248 17536
rect 8668 17484 8720 17536
rect 8944 17484 8996 17536
rect 11704 17484 11756 17536
rect 14096 17552 14148 17604
rect 14832 17595 14884 17604
rect 14004 17484 14056 17536
rect 14832 17561 14841 17595
rect 14841 17561 14875 17595
rect 14875 17561 14884 17595
rect 14832 17552 14884 17561
rect 15476 17629 15485 17663
rect 15485 17629 15519 17663
rect 15519 17629 15528 17663
rect 15476 17620 15528 17629
rect 16672 17620 16724 17672
rect 15384 17552 15436 17604
rect 15844 17552 15896 17604
rect 15936 17552 15988 17604
rect 16948 17552 17000 17604
rect 18052 17620 18104 17672
rect 18236 17663 18288 17672
rect 18236 17629 18245 17663
rect 18245 17629 18279 17663
rect 18279 17629 18288 17663
rect 18236 17620 18288 17629
rect 19984 17663 20036 17672
rect 19984 17629 19993 17663
rect 19993 17629 20027 17663
rect 20027 17629 20036 17663
rect 19984 17620 20036 17629
rect 20168 17663 20220 17672
rect 20168 17629 20177 17663
rect 20177 17629 20211 17663
rect 20211 17629 20220 17663
rect 20168 17620 20220 17629
rect 21916 17620 21968 17672
rect 22560 17620 22612 17672
rect 24032 17756 24084 17808
rect 26608 17756 26660 17808
rect 28632 17756 28684 17808
rect 24584 17663 24636 17672
rect 24584 17629 24593 17663
rect 24593 17629 24627 17663
rect 24627 17629 24636 17663
rect 24584 17620 24636 17629
rect 25504 17688 25556 17740
rect 26700 17688 26752 17740
rect 29920 17731 29972 17740
rect 29920 17697 29929 17731
rect 29929 17697 29963 17731
rect 29963 17697 29972 17731
rect 29920 17688 29972 17697
rect 25044 17663 25096 17672
rect 25044 17629 25053 17663
rect 25053 17629 25087 17663
rect 25087 17629 25096 17663
rect 25044 17620 25096 17629
rect 26056 17620 26108 17672
rect 15108 17484 15160 17536
rect 17132 17484 17184 17536
rect 17684 17527 17736 17536
rect 17684 17493 17693 17527
rect 17693 17493 17727 17527
rect 17727 17493 17736 17527
rect 17684 17484 17736 17493
rect 18972 17484 19024 17536
rect 19340 17484 19392 17536
rect 20352 17484 20404 17536
rect 20628 17484 20680 17536
rect 26148 17552 26200 17604
rect 27804 17552 27856 17604
rect 29276 17552 29328 17604
rect 30564 17552 30616 17604
rect 23020 17484 23072 17536
rect 24216 17484 24268 17536
rect 24952 17484 25004 17536
rect 25780 17484 25832 17536
rect 27620 17484 27672 17536
rect 28264 17527 28316 17536
rect 28264 17493 28273 17527
rect 28273 17493 28307 17527
rect 28307 17493 28316 17527
rect 28264 17484 28316 17493
rect 7288 17382 7340 17434
rect 17592 17382 17644 17434
rect 27896 17382 27948 17434
rect 3516 17212 3568 17264
rect 2688 17144 2740 17196
rect 3884 17280 3936 17332
rect 5448 17323 5500 17332
rect 5448 17289 5457 17323
rect 5457 17289 5491 17323
rect 5491 17289 5500 17323
rect 5448 17280 5500 17289
rect 7196 17280 7248 17332
rect 7932 17280 7984 17332
rect 8024 17280 8076 17332
rect 11612 17280 11664 17332
rect 4988 17255 5040 17264
rect 4988 17221 4997 17255
rect 4997 17221 5031 17255
rect 5031 17221 5040 17255
rect 4988 17212 5040 17221
rect 17684 17280 17736 17332
rect 18052 17280 18104 17332
rect 18144 17280 18196 17332
rect 18696 17280 18748 17332
rect 19156 17280 19208 17332
rect 19984 17280 20036 17332
rect 22560 17280 22612 17332
rect 23112 17323 23164 17332
rect 23112 17289 23121 17323
rect 23121 17289 23155 17323
rect 23155 17289 23164 17323
rect 23112 17280 23164 17289
rect 23204 17280 23256 17332
rect 7748 17144 7800 17196
rect 8944 17187 8996 17196
rect 8944 17153 8953 17187
rect 8953 17153 8987 17187
rect 8987 17153 8996 17187
rect 8944 17144 8996 17153
rect 9220 17187 9272 17196
rect 9220 17153 9254 17187
rect 9254 17153 9272 17187
rect 9220 17144 9272 17153
rect 9496 17144 9548 17196
rect 11704 17187 11756 17196
rect 11704 17153 11713 17187
rect 11713 17153 11747 17187
rect 11747 17153 11756 17187
rect 11704 17144 11756 17153
rect 13820 17212 13872 17264
rect 14004 17212 14056 17264
rect 15384 17212 15436 17264
rect 14740 17144 14792 17196
rect 15016 17144 15068 17196
rect 15844 17144 15896 17196
rect 1860 17008 1912 17060
rect 3884 17008 3936 17060
rect 5172 17008 5224 17060
rect 1768 16940 1820 16992
rect 7472 17008 7524 17060
rect 8484 17076 8536 17128
rect 10600 17076 10652 17128
rect 13544 17076 13596 17128
rect 8024 17008 8076 17060
rect 8208 17008 8260 17060
rect 10232 17008 10284 17060
rect 12256 17008 12308 17060
rect 7012 16940 7064 16992
rect 7380 16940 7432 16992
rect 8392 16940 8444 16992
rect 9680 16940 9732 16992
rect 10876 16940 10928 16992
rect 11888 16983 11940 16992
rect 11888 16949 11897 16983
rect 11897 16949 11931 16983
rect 11931 16949 11940 16983
rect 11888 16940 11940 16949
rect 12164 16940 12216 16992
rect 16672 17144 16724 17196
rect 17132 17212 17184 17264
rect 17408 17212 17460 17264
rect 17868 17255 17920 17264
rect 17040 17187 17092 17196
rect 17040 17153 17049 17187
rect 17049 17153 17083 17187
rect 17083 17153 17092 17187
rect 17040 17144 17092 17153
rect 17868 17221 17902 17255
rect 17902 17221 17920 17255
rect 17868 17212 17920 17221
rect 17960 17212 18012 17264
rect 18880 17144 18932 17196
rect 19800 17212 19852 17264
rect 19984 17144 20036 17196
rect 20352 17187 20404 17196
rect 20352 17153 20361 17187
rect 20361 17153 20395 17187
rect 20395 17153 20404 17187
rect 20352 17144 20404 17153
rect 21824 17212 21876 17264
rect 24308 17280 24360 17332
rect 27160 17280 27212 17332
rect 29092 17280 29144 17332
rect 21732 17144 21784 17196
rect 22192 17187 22244 17196
rect 15752 17008 15804 17060
rect 13912 16983 13964 16992
rect 13912 16949 13921 16983
rect 13921 16949 13955 16983
rect 13955 16949 13964 16983
rect 13912 16940 13964 16949
rect 15476 16940 15528 16992
rect 16948 17008 17000 17060
rect 17408 17008 17460 17060
rect 16212 16940 16264 16992
rect 18880 16940 18932 16992
rect 20720 17076 20772 17128
rect 20904 17076 20956 17128
rect 22192 17153 22201 17187
rect 22201 17153 22235 17187
rect 22235 17153 22244 17187
rect 22192 17144 22244 17153
rect 24676 17212 24728 17264
rect 27252 17212 27304 17264
rect 24216 17187 24268 17196
rect 24216 17153 24225 17187
rect 24225 17153 24259 17187
rect 24259 17153 24268 17187
rect 24216 17144 24268 17153
rect 24492 17187 24544 17196
rect 24492 17153 24501 17187
rect 24501 17153 24535 17187
rect 24535 17153 24544 17187
rect 24492 17144 24544 17153
rect 24860 17144 24912 17196
rect 26608 17144 26660 17196
rect 27620 17187 27672 17196
rect 27620 17153 27629 17187
rect 27629 17153 27663 17187
rect 27663 17153 27672 17187
rect 27620 17144 27672 17153
rect 29092 17144 29144 17196
rect 29828 17144 29880 17196
rect 30840 17212 30892 17264
rect 24952 17119 25004 17128
rect 20168 17008 20220 17060
rect 22928 17008 22980 17060
rect 23204 17008 23256 17060
rect 24952 17085 24961 17119
rect 24961 17085 24995 17119
rect 24995 17085 25004 17119
rect 24952 17076 25004 17085
rect 30012 17076 30064 17128
rect 30472 17076 30524 17128
rect 30656 17144 30708 17196
rect 31024 17144 31076 17196
rect 22100 16940 22152 16992
rect 23388 16940 23440 16992
rect 23756 16940 23808 16992
rect 24492 16940 24544 16992
rect 24768 16940 24820 16992
rect 25228 16940 25280 16992
rect 26056 16940 26108 16992
rect 29184 16940 29236 16992
rect 29460 16983 29512 16992
rect 29460 16949 29469 16983
rect 29469 16949 29503 16983
rect 29503 16949 29512 16983
rect 29460 16940 29512 16949
rect 30840 16940 30892 16992
rect 2136 16838 2188 16890
rect 12440 16838 12492 16890
rect 22744 16838 22796 16890
rect 6920 16736 6972 16788
rect 8852 16736 8904 16788
rect 2596 16600 2648 16652
rect 3792 16643 3844 16652
rect 3792 16609 3801 16643
rect 3801 16609 3835 16643
rect 3835 16609 3844 16643
rect 3792 16600 3844 16609
rect 5264 16600 5316 16652
rect 7840 16600 7892 16652
rect 8392 16643 8444 16652
rect 8392 16609 8401 16643
rect 8401 16609 8435 16643
rect 8435 16609 8444 16643
rect 8392 16600 8444 16609
rect 2044 16532 2096 16584
rect 2780 16532 2832 16584
rect 4252 16532 4304 16584
rect 5448 16532 5500 16584
rect 6552 16532 6604 16584
rect 7196 16575 7248 16584
rect 7196 16541 7205 16575
rect 7205 16541 7239 16575
rect 7239 16541 7248 16575
rect 7380 16575 7432 16584
rect 7196 16532 7248 16541
rect 7380 16541 7389 16575
rect 7389 16541 7423 16575
rect 7423 16541 7432 16575
rect 7380 16532 7432 16541
rect 7564 16532 7616 16584
rect 8576 16532 8628 16584
rect 8944 16600 8996 16652
rect 11428 16736 11480 16788
rect 11980 16736 12032 16788
rect 12164 16736 12216 16788
rect 12624 16779 12676 16788
rect 12624 16745 12633 16779
rect 12633 16745 12667 16779
rect 12667 16745 12676 16779
rect 12624 16736 12676 16745
rect 12256 16668 12308 16720
rect 17316 16668 17368 16720
rect 13820 16600 13872 16652
rect 15108 16600 15160 16652
rect 15292 16600 15344 16652
rect 15384 16600 15436 16652
rect 16764 16643 16816 16652
rect 10508 16532 10560 16584
rect 11060 16532 11112 16584
rect 11980 16532 12032 16584
rect 2596 16507 2648 16516
rect 2596 16473 2605 16507
rect 2605 16473 2639 16507
rect 2639 16473 2648 16507
rect 2596 16464 2648 16473
rect 5540 16507 5592 16516
rect 1492 16396 1544 16448
rect 2044 16396 2096 16448
rect 2412 16396 2464 16448
rect 3148 16439 3200 16448
rect 3148 16405 3157 16439
rect 3157 16405 3191 16439
rect 3191 16405 3200 16439
rect 3148 16396 3200 16405
rect 4804 16439 4856 16448
rect 4804 16405 4813 16439
rect 4813 16405 4847 16439
rect 4847 16405 4856 16439
rect 4804 16396 4856 16405
rect 5540 16473 5549 16507
rect 5549 16473 5583 16507
rect 5583 16473 5592 16507
rect 5540 16464 5592 16473
rect 8208 16464 8260 16516
rect 9220 16464 9272 16516
rect 10968 16464 11020 16516
rect 12808 16464 12860 16516
rect 13176 16464 13228 16516
rect 15476 16532 15528 16584
rect 15108 16464 15160 16516
rect 16764 16609 16773 16643
rect 16773 16609 16807 16643
rect 16807 16609 16816 16643
rect 16764 16600 16816 16609
rect 17408 16600 17460 16652
rect 18880 16600 18932 16652
rect 19156 16600 19208 16652
rect 20996 16668 21048 16720
rect 22376 16736 22428 16788
rect 22928 16736 22980 16788
rect 23388 16736 23440 16788
rect 24032 16736 24084 16788
rect 24216 16736 24268 16788
rect 24400 16779 24452 16788
rect 24400 16745 24409 16779
rect 24409 16745 24443 16779
rect 24443 16745 24452 16779
rect 24400 16736 24452 16745
rect 24676 16736 24728 16788
rect 26056 16736 26108 16788
rect 29920 16668 29972 16720
rect 20904 16600 20956 16652
rect 16304 16532 16356 16584
rect 17040 16532 17092 16584
rect 17776 16575 17828 16584
rect 17776 16541 17785 16575
rect 17785 16541 17819 16575
rect 17819 16541 17828 16575
rect 17776 16532 17828 16541
rect 18236 16532 18288 16584
rect 19524 16575 19576 16584
rect 19524 16541 19533 16575
rect 19533 16541 19567 16575
rect 19567 16541 19576 16575
rect 19524 16532 19576 16541
rect 5724 16396 5776 16448
rect 6736 16396 6788 16448
rect 9496 16396 9548 16448
rect 9772 16396 9824 16448
rect 10600 16396 10652 16448
rect 10784 16439 10836 16448
rect 10784 16405 10793 16439
rect 10793 16405 10827 16439
rect 10827 16405 10836 16439
rect 10784 16396 10836 16405
rect 11428 16396 11480 16448
rect 12164 16396 12216 16448
rect 12256 16396 12308 16448
rect 14832 16396 14884 16448
rect 15384 16396 15436 16448
rect 15568 16396 15620 16448
rect 15844 16396 15896 16448
rect 19800 16464 19852 16516
rect 18604 16396 18656 16448
rect 22284 16532 22336 16584
rect 22376 16532 22428 16584
rect 25044 16600 25096 16652
rect 23112 16532 23164 16584
rect 24308 16532 24360 16584
rect 24492 16532 24544 16584
rect 24584 16532 24636 16584
rect 26148 16600 26200 16652
rect 25228 16532 25280 16584
rect 25780 16532 25832 16584
rect 26700 16532 26752 16584
rect 26792 16532 26844 16584
rect 27252 16532 27304 16584
rect 28356 16532 28408 16584
rect 20076 16396 20128 16448
rect 23480 16464 23532 16516
rect 28540 16464 28592 16516
rect 31392 16464 31444 16516
rect 22284 16396 22336 16448
rect 22560 16396 22612 16448
rect 24032 16396 24084 16448
rect 26056 16396 26108 16448
rect 7288 16294 7340 16346
rect 17592 16294 17644 16346
rect 27896 16294 27948 16346
rect 5540 16192 5592 16244
rect 6368 16192 6420 16244
rect 7380 16192 7432 16244
rect 8208 16192 8260 16244
rect 9220 16235 9272 16244
rect 9220 16201 9229 16235
rect 9229 16201 9263 16235
rect 9263 16201 9272 16235
rect 9220 16192 9272 16201
rect 11796 16235 11848 16244
rect 11796 16201 11805 16235
rect 11805 16201 11839 16235
rect 11839 16201 11848 16235
rect 11796 16192 11848 16201
rect 12348 16192 12400 16244
rect 14372 16192 14424 16244
rect 18052 16192 18104 16244
rect 2228 16124 2280 16176
rect 3148 16124 3200 16176
rect 14832 16124 14884 16176
rect 15292 16124 15344 16176
rect 15844 16124 15896 16176
rect 3884 16056 3936 16108
rect 4436 16056 4488 16108
rect 6000 16056 6052 16108
rect 7564 16056 7616 16108
rect 7840 16056 7892 16108
rect 10324 16099 10376 16108
rect 10324 16065 10333 16099
rect 10333 16065 10367 16099
rect 10367 16065 10376 16099
rect 10324 16056 10376 16065
rect 10784 16099 10836 16108
rect 1400 15988 1452 16040
rect 1860 16031 1912 16040
rect 1860 15997 1869 16031
rect 1869 15997 1903 16031
rect 1903 15997 1912 16031
rect 1860 15988 1912 15997
rect 4344 15920 4396 15972
rect 5080 15920 5132 15972
rect 7472 15988 7524 16040
rect 9680 16031 9732 16040
rect 9680 15997 9689 16031
rect 9689 15997 9723 16031
rect 9723 15997 9732 16031
rect 9680 15988 9732 15997
rect 10784 16065 10793 16099
rect 10793 16065 10827 16099
rect 10827 16065 10836 16099
rect 10784 16056 10836 16065
rect 11520 16056 11572 16108
rect 12072 15988 12124 16040
rect 12624 16056 12676 16108
rect 13636 16056 13688 16108
rect 14372 15988 14424 16040
rect 15016 16056 15068 16108
rect 15476 16056 15528 16108
rect 15660 16056 15712 16108
rect 20260 16235 20312 16244
rect 20260 16201 20269 16235
rect 20269 16201 20303 16235
rect 20303 16201 20312 16235
rect 20260 16192 20312 16201
rect 21272 16192 21324 16244
rect 23480 16192 23532 16244
rect 23664 16235 23716 16244
rect 23664 16201 23673 16235
rect 23673 16201 23707 16235
rect 23707 16201 23716 16235
rect 23664 16192 23716 16201
rect 24400 16192 24452 16244
rect 28264 16192 28316 16244
rect 19156 16167 19208 16176
rect 19156 16133 19190 16167
rect 19190 16133 19208 16167
rect 19156 16124 19208 16133
rect 18880 16099 18932 16108
rect 18880 16065 18889 16099
rect 18889 16065 18923 16099
rect 18923 16065 18932 16099
rect 18880 16056 18932 16065
rect 21456 16124 21508 16176
rect 17040 16031 17092 16040
rect 7196 15920 7248 15972
rect 10048 15920 10100 15972
rect 12164 15920 12216 15972
rect 1860 15852 1912 15904
rect 6644 15852 6696 15904
rect 7380 15852 7432 15904
rect 9496 15852 9548 15904
rect 17040 15997 17049 16031
rect 17049 15997 17083 16031
rect 17083 15997 17092 16031
rect 17040 15988 17092 15997
rect 18052 15988 18104 16040
rect 20260 16056 20312 16108
rect 21916 16056 21968 16108
rect 22100 16099 22152 16108
rect 22100 16065 22134 16099
rect 22134 16065 22152 16099
rect 23204 16124 23256 16176
rect 25228 16124 25280 16176
rect 30380 16124 30432 16176
rect 31300 16192 31352 16244
rect 31484 16124 31536 16176
rect 22100 16056 22152 16065
rect 23572 16056 23624 16108
rect 23940 16056 23992 16108
rect 23388 15988 23440 16040
rect 24400 16056 24452 16108
rect 25964 16056 26016 16108
rect 26056 16099 26108 16108
rect 26056 16065 26065 16099
rect 26065 16065 26099 16099
rect 26099 16065 26108 16099
rect 26056 16056 26108 16065
rect 26976 16056 27028 16108
rect 24676 15988 24728 16040
rect 16948 15920 17000 15972
rect 14832 15852 14884 15904
rect 16304 15852 16356 15904
rect 18512 15852 18564 15904
rect 20996 15852 21048 15904
rect 21272 15895 21324 15904
rect 21272 15861 21281 15895
rect 21281 15861 21315 15895
rect 21315 15861 21324 15895
rect 21272 15852 21324 15861
rect 23112 15852 23164 15904
rect 24400 15920 24452 15972
rect 24584 15920 24636 15972
rect 27252 15988 27304 16040
rect 27528 15988 27580 16040
rect 23664 15852 23716 15904
rect 26240 15852 26292 15904
rect 27436 15895 27488 15904
rect 27436 15861 27445 15895
rect 27445 15861 27479 15895
rect 27479 15861 27488 15895
rect 27436 15852 27488 15861
rect 29000 16056 29052 16108
rect 29276 16056 29328 16108
rect 29920 16056 29972 16108
rect 30656 16056 30708 16108
rect 28448 15920 28500 15972
rect 28908 15852 28960 15904
rect 2136 15750 2188 15802
rect 12440 15750 12492 15802
rect 22744 15750 22796 15802
rect 1492 15648 1544 15700
rect 2596 15648 2648 15700
rect 4804 15648 4856 15700
rect 2872 15623 2924 15632
rect 2872 15589 2881 15623
rect 2881 15589 2915 15623
rect 2915 15589 2924 15623
rect 2872 15580 2924 15589
rect 5080 15580 5132 15632
rect 7472 15648 7524 15700
rect 3792 15512 3844 15564
rect 4344 15555 4396 15564
rect 4344 15521 4353 15555
rect 4353 15521 4387 15555
rect 4387 15521 4396 15555
rect 4344 15512 4396 15521
rect 5448 15555 5500 15564
rect 5448 15521 5457 15555
rect 5457 15521 5491 15555
rect 5491 15521 5500 15555
rect 5448 15512 5500 15521
rect 6644 15580 6696 15632
rect 6552 15512 6604 15564
rect 6828 15555 6880 15564
rect 6828 15521 6837 15555
rect 6837 15521 6871 15555
rect 6871 15521 6880 15555
rect 6828 15512 6880 15521
rect 1860 15444 1912 15496
rect 2412 15444 2464 15496
rect 1492 15376 1544 15428
rect 2320 15376 2372 15428
rect 2412 15308 2464 15360
rect 2504 15308 2556 15360
rect 3056 15351 3108 15360
rect 3056 15317 3065 15351
rect 3065 15317 3099 15351
rect 3099 15317 3108 15351
rect 3056 15308 3108 15317
rect 5540 15376 5592 15428
rect 6276 15308 6328 15360
rect 6736 15351 6788 15360
rect 6736 15317 6745 15351
rect 6745 15317 6779 15351
rect 6779 15317 6788 15351
rect 6736 15308 6788 15317
rect 7748 15580 7800 15632
rect 10508 15580 10560 15632
rect 13820 15648 13872 15700
rect 16488 15648 16540 15700
rect 17960 15648 18012 15700
rect 18328 15648 18380 15700
rect 19524 15691 19576 15700
rect 19524 15657 19533 15691
rect 19533 15657 19567 15691
rect 19567 15657 19576 15691
rect 19524 15648 19576 15657
rect 19892 15648 19944 15700
rect 23664 15648 23716 15700
rect 23940 15648 23992 15700
rect 8576 15512 8628 15564
rect 8944 15555 8996 15564
rect 8944 15521 8953 15555
rect 8953 15521 8987 15555
rect 8987 15521 8996 15555
rect 8944 15512 8996 15521
rect 7196 15444 7248 15496
rect 14004 15512 14056 15564
rect 8484 15376 8536 15428
rect 9312 15376 9364 15428
rect 11428 15487 11480 15496
rect 11428 15453 11437 15487
rect 11437 15453 11471 15487
rect 11471 15453 11480 15487
rect 11428 15444 11480 15453
rect 11796 15376 11848 15428
rect 11980 15444 12032 15496
rect 12348 15444 12400 15496
rect 14188 15444 14240 15496
rect 14464 15487 14516 15496
rect 14464 15453 14473 15487
rect 14473 15453 14507 15487
rect 14507 15453 14516 15487
rect 14464 15444 14516 15453
rect 15936 15444 15988 15496
rect 16488 15444 16540 15496
rect 13176 15376 13228 15428
rect 17040 15512 17092 15564
rect 17868 15555 17920 15564
rect 17868 15521 17877 15555
rect 17877 15521 17911 15555
rect 17911 15521 17920 15555
rect 17868 15512 17920 15521
rect 17960 15512 18012 15564
rect 18696 15512 18748 15564
rect 20352 15512 20404 15564
rect 22928 15512 22980 15564
rect 23112 15512 23164 15564
rect 24768 15580 24820 15632
rect 25596 15648 25648 15700
rect 29000 15691 29052 15700
rect 29000 15657 29009 15691
rect 29009 15657 29043 15691
rect 29043 15657 29052 15691
rect 29000 15648 29052 15657
rect 30564 15648 30616 15700
rect 17684 15444 17736 15496
rect 18788 15444 18840 15496
rect 19708 15487 19760 15496
rect 19708 15453 19717 15487
rect 19717 15453 19751 15487
rect 19751 15453 19760 15487
rect 19708 15444 19760 15453
rect 19984 15487 20036 15496
rect 19984 15453 19993 15487
rect 19993 15453 20027 15487
rect 20027 15453 20036 15487
rect 19984 15444 20036 15453
rect 20260 15444 20312 15496
rect 20812 15487 20864 15496
rect 20812 15453 20821 15487
rect 20821 15453 20855 15487
rect 20855 15453 20864 15487
rect 20812 15444 20864 15453
rect 23756 15487 23808 15496
rect 19248 15376 19300 15428
rect 7656 15351 7708 15360
rect 7656 15317 7665 15351
rect 7665 15317 7699 15351
rect 7699 15317 7708 15351
rect 7656 15308 7708 15317
rect 10508 15308 10560 15360
rect 12164 15308 12216 15360
rect 14188 15308 14240 15360
rect 16212 15308 16264 15360
rect 16856 15308 16908 15360
rect 19524 15308 19576 15360
rect 23388 15376 23440 15428
rect 23756 15453 23765 15487
rect 23765 15453 23799 15487
rect 23799 15453 23808 15487
rect 23756 15444 23808 15453
rect 23664 15376 23716 15428
rect 24308 15444 24360 15496
rect 24768 15487 24820 15496
rect 24768 15453 24777 15487
rect 24777 15453 24811 15487
rect 24811 15453 24820 15487
rect 24768 15444 24820 15453
rect 25596 15487 25648 15496
rect 25596 15453 25605 15487
rect 25605 15453 25639 15487
rect 25639 15453 25648 15487
rect 25596 15444 25648 15453
rect 27620 15512 27672 15564
rect 30380 15580 30432 15632
rect 27712 15487 27764 15496
rect 27712 15453 27721 15487
rect 27721 15453 27755 15487
rect 27755 15453 27764 15487
rect 27712 15444 27764 15453
rect 24860 15376 24912 15428
rect 26884 15376 26936 15428
rect 27252 15376 27304 15428
rect 22008 15308 22060 15360
rect 22836 15308 22888 15360
rect 25780 15308 25832 15360
rect 26976 15351 27028 15360
rect 26976 15317 26985 15351
rect 26985 15317 27019 15351
rect 27019 15317 27028 15351
rect 28264 15376 28316 15428
rect 28908 15444 28960 15496
rect 29828 15444 29880 15496
rect 30012 15487 30064 15496
rect 30012 15453 30021 15487
rect 30021 15453 30055 15487
rect 30055 15453 30064 15487
rect 30012 15444 30064 15453
rect 30196 15487 30248 15496
rect 30196 15453 30205 15487
rect 30205 15453 30239 15487
rect 30239 15453 30248 15487
rect 30196 15444 30248 15453
rect 30840 15487 30892 15496
rect 30840 15453 30849 15487
rect 30849 15453 30883 15487
rect 30883 15453 30892 15487
rect 30840 15444 30892 15453
rect 31116 15487 31168 15496
rect 31116 15453 31125 15487
rect 31125 15453 31159 15487
rect 31159 15453 31168 15487
rect 31116 15444 31168 15453
rect 26976 15308 27028 15317
rect 28724 15308 28776 15360
rect 7288 15206 7340 15258
rect 17592 15206 17644 15258
rect 27896 15206 27948 15258
rect 1676 15104 1728 15156
rect 2228 15104 2280 15156
rect 2872 15104 2924 15156
rect 3884 15104 3936 15156
rect 3976 15104 4028 15156
rect 4896 15104 4948 15156
rect 5448 15104 5500 15156
rect 1492 15079 1544 15088
rect 1492 15045 1501 15079
rect 1501 15045 1535 15079
rect 1535 15045 1544 15079
rect 1492 15036 1544 15045
rect 2320 15036 2372 15088
rect 6092 15104 6144 15156
rect 14096 15104 14148 15156
rect 14924 15104 14976 15156
rect 6828 15079 6880 15088
rect 1032 14968 1084 15020
rect 1676 14968 1728 15020
rect 2504 15011 2556 15020
rect 2504 14977 2513 15011
rect 2513 14977 2547 15011
rect 2547 14977 2556 15011
rect 2504 14968 2556 14977
rect 1952 14900 2004 14952
rect 3608 14968 3660 15020
rect 3976 15011 4028 15020
rect 3976 14977 3985 15011
rect 3985 14977 4019 15011
rect 4019 14977 4028 15011
rect 3976 14968 4028 14977
rect 5080 14968 5132 15020
rect 6828 15045 6837 15079
rect 6837 15045 6871 15079
rect 6871 15045 6880 15079
rect 6828 15036 6880 15045
rect 7656 14968 7708 15020
rect 8944 15036 8996 15088
rect 4436 14943 4488 14952
rect 4436 14909 4445 14943
rect 4445 14909 4479 14943
rect 4479 14909 4488 14943
rect 4436 14900 4488 14909
rect 7012 14900 7064 14952
rect 8392 14968 8444 15020
rect 10048 15011 10100 15020
rect 1860 14764 1912 14816
rect 3516 14764 3568 14816
rect 7748 14832 7800 14884
rect 10048 14977 10057 15011
rect 10057 14977 10091 15011
rect 10091 14977 10100 15011
rect 10048 14968 10100 14977
rect 9220 14900 9272 14952
rect 11336 15036 11388 15088
rect 12164 15079 12216 15088
rect 12164 15045 12198 15079
rect 12198 15045 12216 15079
rect 12164 15036 12216 15045
rect 15660 15104 15712 15156
rect 16212 15104 16264 15156
rect 16948 15104 17000 15156
rect 17776 15104 17828 15156
rect 18144 15104 18196 15156
rect 10508 15011 10560 15020
rect 10508 14977 10517 15011
rect 10517 14977 10551 15011
rect 10551 14977 10560 15011
rect 10508 14968 10560 14977
rect 11244 14968 11296 15020
rect 13820 14968 13872 15020
rect 14648 14968 14700 15020
rect 11060 14900 11112 14952
rect 11888 14943 11940 14952
rect 11888 14909 11897 14943
rect 11897 14909 11931 14943
rect 11931 14909 11940 14943
rect 11888 14900 11940 14909
rect 15844 15036 15896 15088
rect 20996 15104 21048 15156
rect 22100 15147 22152 15156
rect 22100 15113 22109 15147
rect 22109 15113 22143 15147
rect 22143 15113 22152 15147
rect 22100 15104 22152 15113
rect 23664 15104 23716 15156
rect 24032 15104 24084 15156
rect 20260 15036 20312 15088
rect 15108 14968 15160 15020
rect 16120 14968 16172 15020
rect 16764 15011 16816 15020
rect 16764 14977 16773 15011
rect 16773 14977 16807 15011
rect 16807 14977 16816 15011
rect 16764 14968 16816 14977
rect 16948 14968 17000 15020
rect 18512 14968 18564 15020
rect 18880 15011 18932 15020
rect 18880 14977 18889 15011
rect 18889 14977 18923 15011
rect 18923 14977 18932 15011
rect 18880 14968 18932 14977
rect 20904 15011 20956 15020
rect 20904 14977 20913 15011
rect 20913 14977 20947 15011
rect 20947 14977 20956 15011
rect 20904 14968 20956 14977
rect 22192 15036 22244 15088
rect 21272 14968 21324 15020
rect 22284 15011 22336 15020
rect 22284 14977 22293 15011
rect 22293 14977 22327 15011
rect 22327 14977 22336 15011
rect 22284 14968 22336 14977
rect 23388 15011 23440 15020
rect 23388 14977 23422 15011
rect 23422 14977 23440 15011
rect 23940 15036 23992 15088
rect 27436 15104 27488 15156
rect 27712 15104 27764 15156
rect 29368 15104 29420 15156
rect 30196 15104 30248 15156
rect 30656 15147 30708 15156
rect 30656 15113 30665 15147
rect 30665 15113 30699 15147
rect 30699 15113 30708 15147
rect 30656 15104 30708 15113
rect 24952 15036 25004 15088
rect 25596 15036 25648 15088
rect 26332 15036 26384 15088
rect 28264 15036 28316 15088
rect 23388 14968 23440 14977
rect 24768 14968 24820 15020
rect 25228 15011 25280 15020
rect 25228 14977 25237 15011
rect 25237 14977 25271 15011
rect 25271 14977 25280 15011
rect 25228 14968 25280 14977
rect 18144 14900 18196 14952
rect 7196 14764 7248 14816
rect 7380 14764 7432 14816
rect 7472 14764 7524 14816
rect 9404 14764 9456 14816
rect 9496 14764 9548 14816
rect 13544 14832 13596 14884
rect 17868 14832 17920 14884
rect 18328 14875 18380 14884
rect 18328 14841 18337 14875
rect 18337 14841 18371 14875
rect 18371 14841 18380 14875
rect 18328 14832 18380 14841
rect 22192 14900 22244 14952
rect 22928 14900 22980 14952
rect 24492 14900 24544 14952
rect 26148 14968 26200 15020
rect 26976 14968 27028 15020
rect 27252 14968 27304 15020
rect 29000 15036 29052 15088
rect 29920 15036 29972 15088
rect 28632 15011 28684 15020
rect 28632 14977 28666 15011
rect 28666 14977 28684 15011
rect 28632 14968 28684 14977
rect 30748 14968 30800 15020
rect 31024 14968 31076 15020
rect 26792 14900 26844 14952
rect 27344 14943 27396 14952
rect 27344 14909 27353 14943
rect 27353 14909 27387 14943
rect 27387 14909 27396 14943
rect 27344 14900 27396 14909
rect 14740 14764 14792 14816
rect 14924 14764 14976 14816
rect 15660 14764 15712 14816
rect 15752 14764 15804 14816
rect 16028 14764 16080 14816
rect 16212 14764 16264 14816
rect 17408 14764 17460 14816
rect 17684 14764 17736 14816
rect 19892 14764 19944 14816
rect 20720 14764 20772 14816
rect 25228 14832 25280 14884
rect 30380 14832 30432 14884
rect 25044 14764 25096 14816
rect 27068 14764 27120 14816
rect 27160 14807 27212 14816
rect 27160 14773 27169 14807
rect 27169 14773 27203 14807
rect 27203 14773 27212 14807
rect 27160 14764 27212 14773
rect 2136 14662 2188 14714
rect 12440 14662 12492 14714
rect 22744 14662 22796 14714
rect 2688 14560 2740 14612
rect 3516 14560 3568 14612
rect 5448 14560 5500 14612
rect 6828 14560 6880 14612
rect 8208 14560 8260 14612
rect 2412 14492 2464 14544
rect 4068 14492 4120 14544
rect 4620 14424 4672 14476
rect 1400 14399 1452 14408
rect 1400 14365 1409 14399
rect 1409 14365 1443 14399
rect 1443 14365 1452 14399
rect 1400 14356 1452 14365
rect 4160 14356 4212 14408
rect 6092 14424 6144 14476
rect 6276 14467 6328 14476
rect 6276 14433 6285 14467
rect 6285 14433 6319 14467
rect 6319 14433 6328 14467
rect 6276 14424 6328 14433
rect 8760 14424 8812 14476
rect 5172 14399 5224 14408
rect 5172 14365 5181 14399
rect 5181 14365 5215 14399
rect 5215 14365 5224 14399
rect 5172 14356 5224 14365
rect 5356 14356 5408 14408
rect 9772 14560 9824 14612
rect 10508 14560 10560 14612
rect 14004 14560 14056 14612
rect 14188 14560 14240 14612
rect 15200 14560 15252 14612
rect 23388 14603 23440 14612
rect 9956 14492 10008 14544
rect 13544 14535 13596 14544
rect 13544 14501 13553 14535
rect 13553 14501 13587 14535
rect 13587 14501 13596 14535
rect 13544 14492 13596 14501
rect 8944 14424 8996 14476
rect 13176 14424 13228 14476
rect 9588 14356 9640 14408
rect 11704 14356 11756 14408
rect 11888 14356 11940 14408
rect 12164 14399 12216 14408
rect 12164 14365 12173 14399
rect 12173 14365 12207 14399
rect 12207 14365 12216 14399
rect 12164 14356 12216 14365
rect 13820 14356 13872 14408
rect 15476 14424 15528 14476
rect 14740 14399 14792 14408
rect 2688 14288 2740 14340
rect 6920 14288 6972 14340
rect 7748 14331 7800 14340
rect 2780 14263 2832 14272
rect 2780 14229 2789 14263
rect 2789 14229 2823 14263
rect 2823 14229 2832 14263
rect 2780 14220 2832 14229
rect 3516 14220 3568 14272
rect 4344 14220 4396 14272
rect 5448 14220 5500 14272
rect 5724 14220 5776 14272
rect 6184 14220 6236 14272
rect 6552 14220 6604 14272
rect 7748 14297 7757 14331
rect 7757 14297 7791 14331
rect 7791 14297 7800 14331
rect 7748 14288 7800 14297
rect 11980 14288 12032 14340
rect 13452 14288 13504 14340
rect 14740 14365 14749 14399
rect 14749 14365 14783 14399
rect 14783 14365 14792 14399
rect 14740 14356 14792 14365
rect 15016 14356 15068 14408
rect 15936 14424 15988 14476
rect 17316 14424 17368 14476
rect 23388 14569 23397 14603
rect 23397 14569 23431 14603
rect 23431 14569 23440 14603
rect 23388 14560 23440 14569
rect 25964 14603 26016 14612
rect 25964 14569 25973 14603
rect 25973 14569 26007 14603
rect 26007 14569 26016 14603
rect 25964 14560 26016 14569
rect 27436 14603 27488 14612
rect 27436 14569 27445 14603
rect 27445 14569 27479 14603
rect 27479 14569 27488 14603
rect 27436 14560 27488 14569
rect 27620 14560 27672 14612
rect 28632 14560 28684 14612
rect 18696 14492 18748 14544
rect 23296 14492 23348 14544
rect 16120 14356 16172 14408
rect 15108 14288 15160 14340
rect 17040 14356 17092 14408
rect 7932 14220 7984 14272
rect 8208 14220 8260 14272
rect 8300 14220 8352 14272
rect 9404 14220 9456 14272
rect 11612 14263 11664 14272
rect 11612 14229 11621 14263
rect 11621 14229 11655 14263
rect 11655 14229 11664 14263
rect 11612 14220 11664 14229
rect 12992 14220 13044 14272
rect 13728 14220 13780 14272
rect 15752 14220 15804 14272
rect 18236 14220 18288 14272
rect 18696 14288 18748 14340
rect 22836 14424 22888 14476
rect 19432 14356 19484 14408
rect 20628 14356 20680 14408
rect 22376 14356 22428 14408
rect 22560 14356 22612 14408
rect 22928 14399 22980 14408
rect 22928 14365 22937 14399
rect 22937 14365 22971 14399
rect 22971 14365 22980 14399
rect 22928 14356 22980 14365
rect 23664 14356 23716 14408
rect 24308 14356 24360 14408
rect 24952 14492 25004 14544
rect 25044 14492 25096 14544
rect 26240 14492 26292 14544
rect 26332 14492 26384 14544
rect 29736 14492 29788 14544
rect 25964 14424 26016 14476
rect 23388 14288 23440 14340
rect 21180 14220 21232 14272
rect 21364 14263 21416 14272
rect 21364 14229 21373 14263
rect 21373 14229 21407 14263
rect 21407 14229 21416 14263
rect 21364 14220 21416 14229
rect 21824 14220 21876 14272
rect 23296 14220 23348 14272
rect 24032 14220 24084 14272
rect 24492 14288 24544 14340
rect 24860 14220 24912 14272
rect 26240 14356 26292 14408
rect 27160 14399 27212 14408
rect 27160 14365 27169 14399
rect 27169 14365 27203 14399
rect 27203 14365 27212 14399
rect 27160 14356 27212 14365
rect 27252 14356 27304 14408
rect 28724 14399 28776 14408
rect 28724 14365 28733 14399
rect 28733 14365 28767 14399
rect 28767 14365 28776 14399
rect 28724 14356 28776 14365
rect 29184 14356 29236 14408
rect 29460 14356 29512 14408
rect 29920 14288 29972 14340
rect 29276 14220 29328 14272
rect 29644 14220 29696 14272
rect 7288 14118 7340 14170
rect 17592 14118 17644 14170
rect 27896 14118 27948 14170
rect 1860 14016 1912 14068
rect 3056 13991 3108 14000
rect 3056 13957 3065 13991
rect 3065 13957 3099 13991
rect 3099 13957 3108 13991
rect 3056 13948 3108 13957
rect 3148 13991 3200 14000
rect 3148 13957 3157 13991
rect 3157 13957 3191 13991
rect 3191 13957 3200 13991
rect 3516 13991 3568 14000
rect 3148 13948 3200 13957
rect 3516 13957 3525 13991
rect 3525 13957 3559 13991
rect 3559 13957 3568 13991
rect 3516 13948 3568 13957
rect 4252 13948 4304 14000
rect 5540 13948 5592 14000
rect 6184 13948 6236 14000
rect 1308 13880 1360 13932
rect 3976 13880 4028 13932
rect 5264 13880 5316 13932
rect 7932 14016 7984 14068
rect 7656 13948 7708 14000
rect 9588 14016 9640 14068
rect 10508 14016 10560 14068
rect 12624 14016 12676 14068
rect 14648 14059 14700 14068
rect 8392 13880 8444 13932
rect 12992 13948 13044 14000
rect 9128 13880 9180 13932
rect 9496 13923 9548 13932
rect 9496 13889 9505 13923
rect 9505 13889 9539 13923
rect 9539 13889 9548 13923
rect 9496 13880 9548 13889
rect 9956 13880 10008 13932
rect 10048 13880 10100 13932
rect 10232 13880 10284 13932
rect 10508 13923 10560 13932
rect 10508 13889 10517 13923
rect 10517 13889 10551 13923
rect 10551 13889 10560 13923
rect 10508 13880 10560 13889
rect 10876 13880 10928 13932
rect 2320 13812 2372 13864
rect 2780 13812 2832 13864
rect 4620 13855 4672 13864
rect 4620 13821 4629 13855
rect 4629 13821 4663 13855
rect 4663 13821 4672 13855
rect 4620 13812 4672 13821
rect 5448 13812 5500 13864
rect 6552 13787 6604 13796
rect 6552 13753 6561 13787
rect 6561 13753 6595 13787
rect 6595 13753 6604 13787
rect 6552 13744 6604 13753
rect 8300 13812 8352 13864
rect 8760 13812 8812 13864
rect 11612 13880 11664 13932
rect 11980 13923 12032 13932
rect 11980 13889 11989 13923
rect 11989 13889 12023 13923
rect 12023 13889 12032 13923
rect 11980 13880 12032 13889
rect 14648 14025 14657 14059
rect 14657 14025 14691 14059
rect 14691 14025 14700 14059
rect 14648 14016 14700 14025
rect 14740 14016 14792 14068
rect 16212 14016 16264 14068
rect 16672 14059 16724 14068
rect 16672 14025 16681 14059
rect 16681 14025 16715 14059
rect 16715 14025 16724 14059
rect 16672 14016 16724 14025
rect 13176 13880 13228 13932
rect 13452 13880 13504 13932
rect 13544 13923 13596 13932
rect 13544 13889 13553 13923
rect 13553 13889 13587 13923
rect 13587 13889 13596 13923
rect 13544 13880 13596 13889
rect 12348 13855 12400 13864
rect 12348 13821 12357 13855
rect 12357 13821 12391 13855
rect 12391 13821 12400 13855
rect 12348 13812 12400 13821
rect 13912 13812 13964 13864
rect 14648 13880 14700 13932
rect 14832 13923 14884 13932
rect 14832 13889 14841 13923
rect 14841 13889 14875 13923
rect 14875 13889 14884 13923
rect 14832 13880 14884 13889
rect 15384 13880 15436 13932
rect 15844 13880 15896 13932
rect 15936 13923 15988 13932
rect 15936 13889 15945 13923
rect 15945 13889 15979 13923
rect 15979 13889 15988 13923
rect 15936 13880 15988 13889
rect 16488 13880 16540 13932
rect 19248 14016 19300 14068
rect 19984 14016 20036 14068
rect 20996 14016 21048 14068
rect 21732 14016 21784 14068
rect 16948 13880 17000 13932
rect 18144 13948 18196 14000
rect 21364 13948 21416 14000
rect 22928 14016 22980 14068
rect 24676 14016 24728 14068
rect 24860 14016 24912 14068
rect 25136 14016 25188 14068
rect 25964 14016 26016 14068
rect 15568 13812 15620 13864
rect 16212 13812 16264 13864
rect 16764 13812 16816 13864
rect 16856 13812 16908 13864
rect 19892 13880 19944 13932
rect 21180 13880 21232 13932
rect 22928 13880 22980 13932
rect 25228 13880 25280 13932
rect 25504 13880 25556 13932
rect 26148 13948 26200 14000
rect 29092 14016 29144 14068
rect 30932 14016 30984 14068
rect 25780 13923 25832 13932
rect 25780 13889 25789 13923
rect 25789 13889 25823 13923
rect 25823 13889 25832 13923
rect 25780 13880 25832 13889
rect 27068 13880 27120 13932
rect 27528 13880 27580 13932
rect 7656 13744 7708 13796
rect 8024 13787 8076 13796
rect 8024 13753 8033 13787
rect 8033 13753 8067 13787
rect 8067 13753 8076 13787
rect 8024 13744 8076 13753
rect 9312 13787 9364 13796
rect 4344 13676 4396 13728
rect 8668 13719 8720 13728
rect 8668 13685 8677 13719
rect 8677 13685 8711 13719
rect 8711 13685 8720 13719
rect 8668 13676 8720 13685
rect 9312 13753 9321 13787
rect 9321 13753 9355 13787
rect 9355 13753 9364 13787
rect 9312 13744 9364 13753
rect 11060 13676 11112 13728
rect 11520 13676 11572 13728
rect 11704 13676 11756 13728
rect 12992 13676 13044 13728
rect 13544 13676 13596 13728
rect 15016 13719 15068 13728
rect 15016 13685 15025 13719
rect 15025 13685 15059 13719
rect 15059 13685 15068 13719
rect 15016 13676 15068 13685
rect 15384 13676 15436 13728
rect 15568 13719 15620 13728
rect 15568 13685 15577 13719
rect 15577 13685 15611 13719
rect 15611 13685 15620 13719
rect 15568 13676 15620 13685
rect 16120 13744 16172 13796
rect 21364 13812 21416 13864
rect 23756 13812 23808 13864
rect 24676 13855 24728 13864
rect 24676 13821 24685 13855
rect 24685 13821 24719 13855
rect 24719 13821 24728 13855
rect 24676 13812 24728 13821
rect 17408 13744 17460 13796
rect 17684 13676 17736 13728
rect 22836 13744 22888 13796
rect 18328 13676 18380 13728
rect 18696 13676 18748 13728
rect 20996 13676 21048 13728
rect 22008 13676 22060 13728
rect 24216 13719 24268 13728
rect 24216 13685 24225 13719
rect 24225 13685 24259 13719
rect 24259 13685 24268 13719
rect 24216 13676 24268 13685
rect 26884 13744 26936 13796
rect 27160 13744 27212 13796
rect 27804 13812 27856 13864
rect 28724 13948 28776 14000
rect 29184 13880 29236 13932
rect 30932 13880 30984 13932
rect 31116 13923 31168 13932
rect 31116 13889 31125 13923
rect 31125 13889 31159 13923
rect 31159 13889 31168 13923
rect 31116 13880 31168 13889
rect 29092 13812 29144 13864
rect 29736 13812 29788 13864
rect 30840 13855 30892 13864
rect 30840 13821 30849 13855
rect 30849 13821 30883 13855
rect 30883 13821 30892 13855
rect 30840 13812 30892 13821
rect 28632 13719 28684 13728
rect 28632 13685 28641 13719
rect 28641 13685 28675 13719
rect 28675 13685 28684 13719
rect 28632 13676 28684 13685
rect 29644 13719 29696 13728
rect 29644 13685 29653 13719
rect 29653 13685 29687 13719
rect 29687 13685 29696 13719
rect 29644 13676 29696 13685
rect 2136 13574 2188 13626
rect 12440 13574 12492 13626
rect 22744 13574 22796 13626
rect 2688 13515 2740 13524
rect 2688 13481 2697 13515
rect 2697 13481 2731 13515
rect 2731 13481 2740 13515
rect 2688 13472 2740 13481
rect 3056 13515 3108 13524
rect 3056 13481 3065 13515
rect 3065 13481 3099 13515
rect 3099 13481 3108 13515
rect 3056 13472 3108 13481
rect 3148 13472 3200 13524
rect 7104 13515 7156 13524
rect 7104 13481 7113 13515
rect 7113 13481 7147 13515
rect 7147 13481 7156 13515
rect 7104 13472 7156 13481
rect 7472 13472 7524 13524
rect 7748 13472 7800 13524
rect 8668 13472 8720 13524
rect 2320 13404 2372 13456
rect 3608 13404 3660 13456
rect 4712 13404 4764 13456
rect 7564 13404 7616 13456
rect 8024 13404 8076 13456
rect 1492 13336 1544 13388
rect 2504 13268 2556 13320
rect 3976 13336 4028 13388
rect 5448 13336 5500 13388
rect 6828 13336 6880 13388
rect 3792 13268 3844 13320
rect 4988 13268 5040 13320
rect 3976 13243 4028 13252
rect 3976 13209 3985 13243
rect 3985 13209 4019 13243
rect 4019 13209 4028 13243
rect 3976 13200 4028 13209
rect 3516 13132 3568 13184
rect 5540 13200 5592 13252
rect 5724 13268 5776 13320
rect 6920 13268 6972 13320
rect 8392 13404 8444 13456
rect 8484 13404 8536 13456
rect 10416 13404 10468 13456
rect 11520 13404 11572 13456
rect 9404 13379 9456 13388
rect 9404 13345 9413 13379
rect 9413 13345 9447 13379
rect 9447 13345 9456 13379
rect 9404 13336 9456 13345
rect 8760 13200 8812 13252
rect 4804 13132 4856 13184
rect 6184 13175 6236 13184
rect 6184 13141 6193 13175
rect 6193 13141 6227 13175
rect 6227 13141 6236 13175
rect 6184 13132 6236 13141
rect 7104 13132 7156 13184
rect 7656 13132 7708 13184
rect 12164 13268 12216 13320
rect 12624 13268 12676 13320
rect 15108 13404 15160 13456
rect 15936 13404 15988 13456
rect 16764 13472 16816 13524
rect 16856 13472 16908 13524
rect 17132 13472 17184 13524
rect 17776 13472 17828 13524
rect 18144 13404 18196 13456
rect 18328 13472 18380 13524
rect 19340 13472 19392 13524
rect 19800 13404 19852 13456
rect 21732 13472 21784 13524
rect 22100 13472 22152 13524
rect 23572 13472 23624 13524
rect 24308 13472 24360 13524
rect 25504 13472 25556 13524
rect 25780 13472 25832 13524
rect 26516 13472 26568 13524
rect 27160 13472 27212 13524
rect 27344 13472 27396 13524
rect 28632 13472 28684 13524
rect 29092 13472 29144 13524
rect 29920 13515 29972 13524
rect 29920 13481 29929 13515
rect 29929 13481 29963 13515
rect 29963 13481 29972 13515
rect 29920 13472 29972 13481
rect 30932 13515 30984 13524
rect 30932 13481 30941 13515
rect 30941 13481 30975 13515
rect 30975 13481 30984 13515
rect 30932 13472 30984 13481
rect 31116 13515 31168 13524
rect 31116 13481 31125 13515
rect 31125 13481 31159 13515
rect 31159 13481 31168 13515
rect 31116 13472 31168 13481
rect 25964 13404 26016 13456
rect 12992 13311 13044 13320
rect 12992 13277 13001 13311
rect 13001 13277 13035 13311
rect 13035 13277 13044 13311
rect 12992 13268 13044 13277
rect 14188 13268 14240 13320
rect 14648 13268 14700 13320
rect 11336 13200 11388 13252
rect 13912 13200 13964 13252
rect 14924 13200 14976 13252
rect 15108 13268 15160 13320
rect 12348 13175 12400 13184
rect 12348 13141 12357 13175
rect 12357 13141 12391 13175
rect 12391 13141 12400 13175
rect 12348 13132 12400 13141
rect 12808 13132 12860 13184
rect 15108 13132 15160 13184
rect 15752 13336 15804 13388
rect 16212 13379 16264 13388
rect 16212 13345 16221 13379
rect 16221 13345 16255 13379
rect 16255 13345 16264 13379
rect 16212 13336 16264 13345
rect 16304 13268 16356 13320
rect 16488 13268 16540 13320
rect 19432 13336 19484 13388
rect 19984 13379 20036 13388
rect 19984 13345 19993 13379
rect 19993 13345 20027 13379
rect 20027 13345 20036 13379
rect 19984 13336 20036 13345
rect 20996 13336 21048 13388
rect 22376 13336 22428 13388
rect 22560 13336 22612 13388
rect 24768 13379 24820 13388
rect 15844 13200 15896 13252
rect 17500 13200 17552 13252
rect 18788 13268 18840 13320
rect 19156 13268 19208 13320
rect 17960 13243 18012 13252
rect 17960 13209 17969 13243
rect 17969 13209 18003 13243
rect 18003 13209 18012 13243
rect 17960 13200 18012 13209
rect 18144 13200 18196 13252
rect 21824 13268 21876 13320
rect 23388 13311 23440 13320
rect 23388 13277 23397 13311
rect 23397 13277 23431 13311
rect 23431 13277 23440 13311
rect 23388 13268 23440 13277
rect 24768 13345 24777 13379
rect 24777 13345 24811 13379
rect 24811 13345 24820 13379
rect 24768 13336 24820 13345
rect 27068 13379 27120 13388
rect 27068 13345 27077 13379
rect 27077 13345 27111 13379
rect 27111 13345 27120 13379
rect 27068 13336 27120 13345
rect 23940 13268 23992 13320
rect 24216 13268 24268 13320
rect 26792 13311 26844 13320
rect 26792 13277 26801 13311
rect 26801 13277 26835 13311
rect 26835 13277 26844 13311
rect 26792 13268 26844 13277
rect 22560 13200 22612 13252
rect 22928 13200 22980 13252
rect 19248 13132 19300 13184
rect 21916 13132 21968 13184
rect 23572 13132 23624 13184
rect 24676 13200 24728 13252
rect 25688 13200 25740 13252
rect 27712 13336 27764 13388
rect 28724 13336 28776 13388
rect 26332 13132 26384 13184
rect 26976 13132 27028 13184
rect 28908 13268 28960 13320
rect 30196 13268 30248 13320
rect 29644 13200 29696 13252
rect 27620 13132 27672 13184
rect 28724 13132 28776 13184
rect 28816 13175 28868 13184
rect 28816 13141 28841 13175
rect 28841 13141 28868 13175
rect 29552 13175 29604 13184
rect 28816 13132 28868 13141
rect 29552 13141 29561 13175
rect 29561 13141 29595 13175
rect 29595 13141 29604 13175
rect 29552 13132 29604 13141
rect 31024 13132 31076 13184
rect 7288 13030 7340 13082
rect 17592 13030 17644 13082
rect 27896 13030 27948 13082
rect 3516 12928 3568 12980
rect 1492 12903 1544 12912
rect 1492 12869 1501 12903
rect 1501 12869 1535 12903
rect 1535 12869 1544 12903
rect 1492 12860 1544 12869
rect 2320 12835 2372 12844
rect 2320 12801 2329 12835
rect 2329 12801 2363 12835
rect 2363 12801 2372 12835
rect 2320 12792 2372 12801
rect 2872 12860 2924 12912
rect 2780 12835 2832 12844
rect 2780 12801 2789 12835
rect 2789 12801 2823 12835
rect 2823 12801 2832 12835
rect 2780 12792 2832 12801
rect 1308 12724 1360 12776
rect 1860 12656 1912 12708
rect 2412 12724 2464 12776
rect 4804 12971 4856 12980
rect 4804 12937 4813 12971
rect 4813 12937 4847 12971
rect 4847 12937 4856 12971
rect 4804 12928 4856 12937
rect 7564 12928 7616 12980
rect 4068 12860 4120 12912
rect 5356 12860 5408 12912
rect 4344 12835 4396 12844
rect 4344 12801 4353 12835
rect 4353 12801 4387 12835
rect 4387 12801 4396 12835
rect 4344 12792 4396 12801
rect 5908 12792 5960 12844
rect 6276 12792 6328 12844
rect 7104 12860 7156 12912
rect 8208 12928 8260 12980
rect 8668 12928 8720 12980
rect 14188 12928 14240 12980
rect 14924 12928 14976 12980
rect 20168 12928 20220 12980
rect 20720 12928 20772 12980
rect 25964 12928 26016 12980
rect 26792 12928 26844 12980
rect 29644 12971 29696 12980
rect 29644 12937 29653 12971
rect 29653 12937 29687 12971
rect 29687 12937 29696 12971
rect 29644 12928 29696 12937
rect 11520 12860 11572 12912
rect 7840 12835 7892 12844
rect 7840 12801 7869 12835
rect 7869 12801 7892 12835
rect 7840 12792 7892 12801
rect 8208 12792 8260 12844
rect 8392 12792 8444 12844
rect 8760 12835 8812 12844
rect 8760 12801 8769 12835
rect 8769 12801 8803 12835
rect 8803 12801 8812 12835
rect 8760 12792 8812 12801
rect 9680 12792 9732 12844
rect 9772 12835 9824 12844
rect 9772 12801 9781 12835
rect 9781 12801 9815 12835
rect 9815 12801 9824 12835
rect 9772 12792 9824 12801
rect 10784 12792 10836 12844
rect 15568 12860 15620 12912
rect 16580 12860 16632 12912
rect 12348 12792 12400 12844
rect 12532 12835 12584 12844
rect 12532 12801 12541 12835
rect 12541 12801 12575 12835
rect 12575 12801 12584 12835
rect 12532 12792 12584 12801
rect 12624 12792 12676 12844
rect 13268 12835 13320 12844
rect 13268 12801 13277 12835
rect 13277 12801 13311 12835
rect 13311 12801 13320 12835
rect 13268 12792 13320 12801
rect 13912 12835 13964 12844
rect 13912 12801 13921 12835
rect 13921 12801 13955 12835
rect 13955 12801 13964 12835
rect 13912 12792 13964 12801
rect 14096 12835 14148 12844
rect 14096 12801 14105 12835
rect 14105 12801 14139 12835
rect 14139 12801 14148 12835
rect 14096 12792 14148 12801
rect 14556 12792 14608 12844
rect 14740 12835 14792 12844
rect 14740 12801 14749 12835
rect 14749 12801 14783 12835
rect 14783 12801 14792 12835
rect 14740 12792 14792 12801
rect 16764 12835 16816 12844
rect 16764 12801 16773 12835
rect 16773 12801 16807 12835
rect 16807 12801 16816 12835
rect 16764 12792 16816 12801
rect 3976 12724 4028 12776
rect 5632 12724 5684 12776
rect 6552 12724 6604 12776
rect 8300 12724 8352 12776
rect 11888 12767 11940 12776
rect 11888 12733 11897 12767
rect 11897 12733 11931 12767
rect 11931 12733 11940 12767
rect 11888 12724 11940 12733
rect 13176 12724 13228 12776
rect 16028 12724 16080 12776
rect 16488 12724 16540 12776
rect 18604 12860 18656 12912
rect 19156 12860 19208 12912
rect 19892 12860 19944 12912
rect 17868 12792 17920 12844
rect 18144 12835 18196 12844
rect 17500 12724 17552 12776
rect 18144 12801 18153 12835
rect 18153 12801 18187 12835
rect 18187 12801 18196 12835
rect 18144 12792 18196 12801
rect 22376 12860 22428 12912
rect 24492 12860 24544 12912
rect 20536 12835 20588 12844
rect 16120 12699 16172 12708
rect 2228 12588 2280 12640
rect 3608 12631 3660 12640
rect 3608 12597 3617 12631
rect 3617 12597 3651 12631
rect 3651 12597 3660 12631
rect 3608 12588 3660 12597
rect 5172 12588 5224 12640
rect 7656 12588 7708 12640
rect 9220 12588 9272 12640
rect 10416 12631 10468 12640
rect 10416 12597 10425 12631
rect 10425 12597 10459 12631
rect 10459 12597 10468 12631
rect 10416 12588 10468 12597
rect 11336 12588 11388 12640
rect 13360 12631 13412 12640
rect 13360 12597 13369 12631
rect 13369 12597 13403 12631
rect 13403 12597 13412 12631
rect 13360 12588 13412 12597
rect 16120 12665 16129 12699
rect 16129 12665 16163 12699
rect 16163 12665 16172 12699
rect 16120 12656 16172 12665
rect 16948 12588 17000 12640
rect 17040 12588 17092 12640
rect 20536 12801 20545 12835
rect 20545 12801 20579 12835
rect 20579 12801 20588 12835
rect 20536 12792 20588 12801
rect 21916 12792 21968 12844
rect 23296 12792 23348 12844
rect 25044 12835 25096 12844
rect 25044 12801 25053 12835
rect 25053 12801 25087 12835
rect 25087 12801 25096 12835
rect 25044 12792 25096 12801
rect 25504 12860 25556 12912
rect 25688 12792 25740 12844
rect 25872 12792 25924 12844
rect 27712 12860 27764 12912
rect 27436 12835 27488 12844
rect 20260 12724 20312 12776
rect 20444 12724 20496 12776
rect 21548 12724 21600 12776
rect 21364 12656 21416 12708
rect 19800 12631 19852 12640
rect 19800 12597 19809 12631
rect 19809 12597 19843 12631
rect 19843 12597 19852 12631
rect 20352 12631 20404 12640
rect 19800 12588 19852 12597
rect 20352 12597 20361 12631
rect 20361 12597 20395 12631
rect 20395 12597 20404 12631
rect 20352 12588 20404 12597
rect 20812 12588 20864 12640
rect 22560 12588 22612 12640
rect 23940 12588 23992 12640
rect 24952 12724 25004 12776
rect 26148 12724 26200 12776
rect 27436 12801 27445 12835
rect 27445 12801 27479 12835
rect 27479 12801 27488 12835
rect 27436 12792 27488 12801
rect 27620 12835 27672 12844
rect 27620 12801 27629 12835
rect 27629 12801 27663 12835
rect 27663 12801 27672 12835
rect 27620 12792 27672 12801
rect 29000 12860 29052 12912
rect 29552 12792 29604 12844
rect 30288 12792 30340 12844
rect 30932 12792 30984 12844
rect 31208 12792 31260 12844
rect 29920 12724 29972 12776
rect 27344 12656 27396 12708
rect 25228 12631 25280 12640
rect 25228 12597 25237 12631
rect 25237 12597 25271 12631
rect 25271 12597 25280 12631
rect 25228 12588 25280 12597
rect 25964 12588 26016 12640
rect 30196 12588 30248 12640
rect 2136 12486 2188 12538
rect 12440 12486 12492 12538
rect 22744 12486 22796 12538
rect 2964 12384 3016 12436
rect 3884 12384 3936 12436
rect 5908 12427 5960 12436
rect 3056 12248 3108 12300
rect 3608 12248 3660 12300
rect 5908 12393 5917 12427
rect 5917 12393 5951 12427
rect 5951 12393 5960 12427
rect 5908 12384 5960 12393
rect 6184 12384 6236 12436
rect 7656 12384 7708 12436
rect 8668 12384 8720 12436
rect 9128 12384 9180 12436
rect 13268 12384 13320 12436
rect 13728 12384 13780 12436
rect 6460 12316 6512 12368
rect 6644 12316 6696 12368
rect 7380 12316 7432 12368
rect 11520 12316 11572 12368
rect 15384 12384 15436 12436
rect 16304 12316 16356 12368
rect 6276 12248 6328 12300
rect 1400 12223 1452 12232
rect 1400 12189 1409 12223
rect 1409 12189 1443 12223
rect 1443 12189 1452 12223
rect 1400 12180 1452 12189
rect 4436 12180 4488 12232
rect 6460 12223 6512 12232
rect 6460 12189 6469 12223
rect 6469 12189 6503 12223
rect 6503 12189 6512 12223
rect 6460 12180 6512 12189
rect 6644 12180 6696 12232
rect 7472 12180 7524 12232
rect 7840 12180 7892 12232
rect 2228 12112 2280 12164
rect 2320 12112 2372 12164
rect 3792 12112 3844 12164
rect 4896 12112 4948 12164
rect 5356 12112 5408 12164
rect 8576 12248 8628 12300
rect 8944 12291 8996 12300
rect 8944 12257 8953 12291
rect 8953 12257 8987 12291
rect 8987 12257 8996 12291
rect 8944 12248 8996 12257
rect 9220 12223 9272 12232
rect 9220 12189 9254 12223
rect 9254 12189 9272 12223
rect 10784 12223 10836 12232
rect 9220 12180 9272 12189
rect 10784 12189 10793 12223
rect 10793 12189 10827 12223
rect 10827 12189 10836 12223
rect 10784 12180 10836 12189
rect 11060 12223 11112 12232
rect 11060 12189 11069 12223
rect 11069 12189 11103 12223
rect 11103 12189 11112 12223
rect 11060 12180 11112 12189
rect 12624 12180 12676 12232
rect 13636 12248 13688 12300
rect 15108 12248 15160 12300
rect 16028 12248 16080 12300
rect 13544 12223 13596 12232
rect 13544 12189 13553 12223
rect 13553 12189 13587 12223
rect 13587 12189 13596 12223
rect 13544 12180 13596 12189
rect 13820 12180 13872 12232
rect 14740 12180 14792 12232
rect 17960 12384 18012 12436
rect 18144 12384 18196 12436
rect 19340 12384 19392 12436
rect 17776 12316 17828 12368
rect 18972 12316 19024 12368
rect 20536 12384 20588 12436
rect 20904 12384 20956 12436
rect 21640 12427 21692 12436
rect 21640 12393 21649 12427
rect 21649 12393 21683 12427
rect 21683 12393 21692 12427
rect 21640 12384 21692 12393
rect 23296 12384 23348 12436
rect 23480 12384 23532 12436
rect 26516 12384 26568 12436
rect 20720 12316 20772 12368
rect 24124 12316 24176 12368
rect 27712 12384 27764 12436
rect 28080 12384 28132 12436
rect 28724 12427 28776 12436
rect 28724 12393 28733 12427
rect 28733 12393 28767 12427
rect 28767 12393 28776 12427
rect 28724 12384 28776 12393
rect 31024 12384 31076 12436
rect 11244 12112 11296 12164
rect 16856 12112 16908 12164
rect 16948 12112 17000 12164
rect 18328 12112 18380 12164
rect 3700 12044 3752 12096
rect 4712 12044 4764 12096
rect 5724 12044 5776 12096
rect 7012 12044 7064 12096
rect 7472 12044 7524 12096
rect 7656 12087 7708 12096
rect 7656 12053 7665 12087
rect 7665 12053 7699 12087
rect 7699 12053 7708 12087
rect 7656 12044 7708 12053
rect 7840 12044 7892 12096
rect 8760 12044 8812 12096
rect 9404 12044 9456 12096
rect 12808 12087 12860 12096
rect 12808 12053 12817 12087
rect 12817 12053 12851 12087
rect 12851 12053 12860 12087
rect 12808 12044 12860 12053
rect 14556 12044 14608 12096
rect 15936 12044 15988 12096
rect 16764 12044 16816 12096
rect 18420 12044 18472 12096
rect 19156 12180 19208 12232
rect 19708 12180 19760 12232
rect 20076 12223 20128 12232
rect 20076 12189 20085 12223
rect 20085 12189 20119 12223
rect 20119 12189 20128 12223
rect 20076 12180 20128 12189
rect 20260 12223 20312 12232
rect 20260 12189 20269 12223
rect 20269 12189 20303 12223
rect 20303 12189 20312 12223
rect 20260 12180 20312 12189
rect 20536 12180 20588 12232
rect 21456 12223 21508 12232
rect 21456 12189 21465 12223
rect 21465 12189 21499 12223
rect 21499 12189 21508 12223
rect 21456 12180 21508 12189
rect 18972 12112 19024 12164
rect 21364 12112 21416 12164
rect 23112 12248 23164 12300
rect 23480 12248 23532 12300
rect 23664 12248 23716 12300
rect 22560 12223 22612 12232
rect 22560 12189 22569 12223
rect 22569 12189 22603 12223
rect 22603 12189 22612 12223
rect 22560 12180 22612 12189
rect 23572 12223 23624 12232
rect 23572 12189 23581 12223
rect 23581 12189 23615 12223
rect 23615 12189 23624 12223
rect 23572 12180 23624 12189
rect 24952 12223 25004 12232
rect 24952 12189 24961 12223
rect 24961 12189 24995 12223
rect 24995 12189 25004 12223
rect 24952 12180 25004 12189
rect 25044 12180 25096 12232
rect 25964 12223 26016 12232
rect 23664 12112 23716 12164
rect 24032 12112 24084 12164
rect 25964 12189 25973 12223
rect 25973 12189 26007 12223
rect 26007 12189 26016 12223
rect 25964 12180 26016 12189
rect 26700 12223 26752 12232
rect 25412 12112 25464 12164
rect 26700 12189 26709 12223
rect 26709 12189 26743 12223
rect 26743 12189 26752 12223
rect 26700 12180 26752 12189
rect 26976 12223 27028 12232
rect 26976 12189 27010 12223
rect 27010 12189 27028 12223
rect 26976 12180 27028 12189
rect 27620 12112 27672 12164
rect 27988 12112 28040 12164
rect 29000 12248 29052 12300
rect 30196 12223 30248 12232
rect 30196 12189 30230 12223
rect 30230 12189 30248 12223
rect 30196 12180 30248 12189
rect 23388 12044 23440 12096
rect 23572 12044 23624 12096
rect 24308 12044 24360 12096
rect 24768 12087 24820 12096
rect 24768 12053 24777 12087
rect 24777 12053 24811 12087
rect 24811 12053 24820 12087
rect 24768 12044 24820 12053
rect 26792 12044 26844 12096
rect 30840 12112 30892 12164
rect 28172 12044 28224 12096
rect 30012 12044 30064 12096
rect 7288 11942 7340 11994
rect 17592 11942 17644 11994
rect 27896 11942 27948 11994
rect 2504 11840 2556 11892
rect 9956 11840 10008 11892
rect 11152 11840 11204 11892
rect 13176 11883 13228 11892
rect 13176 11849 13185 11883
rect 13185 11849 13219 11883
rect 13219 11849 13228 11883
rect 13176 11840 13228 11849
rect 3700 11772 3752 11824
rect 1952 11747 2004 11756
rect 1952 11713 1961 11747
rect 1961 11713 1995 11747
rect 1995 11713 2004 11747
rect 1952 11704 2004 11713
rect 1584 11636 1636 11688
rect 1768 11568 1820 11620
rect 4528 11704 4580 11756
rect 4988 11704 5040 11756
rect 7196 11704 7248 11756
rect 7564 11704 7616 11756
rect 7932 11704 7984 11756
rect 8668 11704 8720 11756
rect 9404 11747 9456 11756
rect 9404 11713 9413 11747
rect 9413 11713 9447 11747
rect 9447 11713 9456 11747
rect 9404 11704 9456 11713
rect 9772 11704 9824 11756
rect 10140 11704 10192 11756
rect 12072 11747 12124 11756
rect 12072 11713 12106 11747
rect 12106 11713 12124 11747
rect 12072 11704 12124 11713
rect 13268 11772 13320 11824
rect 15844 11840 15896 11892
rect 23664 11883 23716 11892
rect 16856 11815 16908 11824
rect 16856 11781 16865 11815
rect 16865 11781 16899 11815
rect 16899 11781 16908 11815
rect 16856 11772 16908 11781
rect 17500 11772 17552 11824
rect 12624 11704 12676 11756
rect 12808 11704 12860 11756
rect 17040 11747 17092 11756
rect 17040 11713 17049 11747
rect 17049 11713 17083 11747
rect 17083 11713 17092 11747
rect 17040 11704 17092 11713
rect 17684 11704 17736 11756
rect 17868 11704 17920 11756
rect 18972 11772 19024 11824
rect 20168 11772 20220 11824
rect 21364 11772 21416 11824
rect 23664 11849 23673 11883
rect 23673 11849 23707 11883
rect 23707 11849 23716 11883
rect 23664 11840 23716 11849
rect 24768 11840 24820 11892
rect 28172 11840 28224 11892
rect 28908 11883 28960 11892
rect 28908 11849 28917 11883
rect 28917 11849 28951 11883
rect 28951 11849 28960 11883
rect 28908 11840 28960 11849
rect 29552 11840 29604 11892
rect 30288 11883 30340 11892
rect 30288 11849 30297 11883
rect 30297 11849 30331 11883
rect 30331 11849 30340 11883
rect 30288 11840 30340 11849
rect 2688 11679 2740 11688
rect 2688 11645 2697 11679
rect 2697 11645 2731 11679
rect 2731 11645 2740 11679
rect 2688 11636 2740 11645
rect 4620 11636 4672 11688
rect 6092 11636 6144 11688
rect 6644 11636 6696 11688
rect 7104 11636 7156 11688
rect 7840 11636 7892 11688
rect 10324 11636 10376 11688
rect 11796 11679 11848 11688
rect 11796 11645 11805 11679
rect 11805 11645 11839 11679
rect 11839 11645 11848 11679
rect 11796 11636 11848 11645
rect 14280 11679 14332 11688
rect 3056 11500 3108 11552
rect 5264 11500 5316 11552
rect 6184 11500 6236 11552
rect 8300 11500 8352 11552
rect 9128 11500 9180 11552
rect 12900 11568 12952 11620
rect 14280 11645 14289 11679
rect 14289 11645 14323 11679
rect 14323 11645 14332 11679
rect 14280 11636 14332 11645
rect 16120 11636 16172 11688
rect 19156 11636 19208 11688
rect 12992 11500 13044 11552
rect 13636 11543 13688 11552
rect 13636 11509 13645 11543
rect 13645 11509 13679 11543
rect 13679 11509 13688 11543
rect 13636 11500 13688 11509
rect 18512 11568 18564 11620
rect 17316 11500 17368 11552
rect 17500 11500 17552 11552
rect 20352 11704 20404 11756
rect 23572 11747 23624 11756
rect 23572 11713 23581 11747
rect 23581 11713 23615 11747
rect 23615 11713 23624 11747
rect 23572 11704 23624 11713
rect 23940 11747 23992 11756
rect 20628 11636 20680 11688
rect 21640 11568 21692 11620
rect 22100 11611 22152 11620
rect 22100 11577 22109 11611
rect 22109 11577 22143 11611
rect 22143 11577 22152 11611
rect 22100 11568 22152 11577
rect 23020 11568 23072 11620
rect 23204 11568 23256 11620
rect 23940 11713 23949 11747
rect 23949 11713 23983 11747
rect 23983 11713 23992 11747
rect 23940 11704 23992 11713
rect 20444 11500 20496 11552
rect 20628 11500 20680 11552
rect 23296 11500 23348 11552
rect 24584 11772 24636 11824
rect 25412 11772 25464 11824
rect 27988 11772 28040 11824
rect 29092 11747 29144 11756
rect 29092 11713 29101 11747
rect 29101 11713 29135 11747
rect 29135 11713 29144 11747
rect 29092 11704 29144 11713
rect 29368 11747 29420 11756
rect 29368 11713 29377 11747
rect 29377 11713 29411 11747
rect 29411 11713 29420 11747
rect 29368 11704 29420 11713
rect 29644 11704 29696 11756
rect 29736 11704 29788 11756
rect 28080 11636 28132 11688
rect 31024 11704 31076 11756
rect 31300 11568 31352 11620
rect 25228 11543 25280 11552
rect 25228 11509 25237 11543
rect 25237 11509 25271 11543
rect 25271 11509 25280 11543
rect 25228 11500 25280 11509
rect 26056 11543 26108 11552
rect 26056 11509 26065 11543
rect 26065 11509 26099 11543
rect 26099 11509 26108 11543
rect 26056 11500 26108 11509
rect 29092 11500 29144 11552
rect 29736 11500 29788 11552
rect 2136 11398 2188 11450
rect 12440 11398 12492 11450
rect 22744 11398 22796 11450
rect 2412 11296 2464 11348
rect 3608 11296 3660 11348
rect 4160 11296 4212 11348
rect 5080 11339 5132 11348
rect 5080 11305 5089 11339
rect 5089 11305 5123 11339
rect 5123 11305 5132 11339
rect 5080 11296 5132 11305
rect 12348 11296 12400 11348
rect 13728 11296 13780 11348
rect 15200 11296 15252 11348
rect 15384 11296 15436 11348
rect 1860 11092 1912 11144
rect 3148 11160 3200 11212
rect 5540 11203 5592 11212
rect 5540 11169 5549 11203
rect 5549 11169 5583 11203
rect 5583 11169 5592 11203
rect 5540 11160 5592 11169
rect 6368 11160 6420 11212
rect 2780 11135 2832 11144
rect 2780 11101 2789 11135
rect 2789 11101 2823 11135
rect 2823 11101 2832 11135
rect 2964 11135 3016 11144
rect 2780 11092 2832 11101
rect 2964 11101 2973 11135
rect 2973 11101 3007 11135
rect 3007 11101 3016 11135
rect 2964 11092 3016 11101
rect 2872 11024 2924 11076
rect 4252 11092 4304 11144
rect 4436 11092 4488 11144
rect 5264 11135 5316 11144
rect 5264 11101 5273 11135
rect 5273 11101 5307 11135
rect 5307 11101 5316 11135
rect 5264 11092 5316 11101
rect 9496 11228 9548 11280
rect 13636 11228 13688 11280
rect 17316 11296 17368 11348
rect 17684 11228 17736 11280
rect 7656 11160 7708 11212
rect 9680 11203 9732 11212
rect 7932 11092 7984 11144
rect 8208 11135 8260 11144
rect 8208 11101 8217 11135
rect 8217 11101 8251 11135
rect 8251 11101 8260 11135
rect 8208 11092 8260 11101
rect 6184 11067 6236 11076
rect 6184 11033 6193 11067
rect 6193 11033 6227 11067
rect 6227 11033 6236 11067
rect 6184 11024 6236 11033
rect 6460 11067 6512 11076
rect 6460 11033 6469 11067
rect 6469 11033 6503 11067
rect 6503 11033 6512 11067
rect 6460 11024 6512 11033
rect 6552 11067 6604 11076
rect 6552 11033 6561 11067
rect 6561 11033 6595 11067
rect 6595 11033 6604 11067
rect 6552 11024 6604 11033
rect 6736 11024 6788 11076
rect 2228 10956 2280 11008
rect 6000 10956 6052 11008
rect 7104 10956 7156 11008
rect 7932 10956 7984 11008
rect 8024 10956 8076 11008
rect 9036 11092 9088 11144
rect 9680 11169 9689 11203
rect 9689 11169 9723 11203
rect 9723 11169 9732 11203
rect 9680 11160 9732 11169
rect 9864 11135 9916 11144
rect 9864 11101 9873 11135
rect 9873 11101 9907 11135
rect 9907 11101 9916 11135
rect 9864 11092 9916 11101
rect 10416 11160 10468 11212
rect 10324 11135 10376 11144
rect 10324 11101 10333 11135
rect 10333 11101 10367 11135
rect 10367 11101 10376 11135
rect 10324 11092 10376 11101
rect 12624 11160 12676 11212
rect 11796 11092 11848 11144
rect 12992 11160 13044 11212
rect 14096 11092 14148 11144
rect 17500 11160 17552 11212
rect 18328 11160 18380 11212
rect 8944 11067 8996 11076
rect 8944 11033 8953 11067
rect 8953 11033 8987 11067
rect 8987 11033 8996 11067
rect 8944 11024 8996 11033
rect 9128 11067 9180 11076
rect 9128 11033 9137 11067
rect 9137 11033 9171 11067
rect 9171 11033 9180 11067
rect 9128 11024 9180 11033
rect 12716 11024 12768 11076
rect 18236 11135 18288 11144
rect 18236 11101 18245 11135
rect 18245 11101 18279 11135
rect 18279 11101 18288 11135
rect 18236 11092 18288 11101
rect 21180 11296 21232 11348
rect 22192 11228 22244 11280
rect 23480 11228 23532 11280
rect 28080 11271 28132 11280
rect 28080 11237 28089 11271
rect 28089 11237 28123 11271
rect 28123 11237 28132 11271
rect 28080 11228 28132 11237
rect 29920 11296 29972 11348
rect 29184 11228 29236 11280
rect 20444 11160 20496 11212
rect 20812 11203 20864 11212
rect 20812 11169 20821 11203
rect 20821 11169 20855 11203
rect 20855 11169 20864 11203
rect 20812 11160 20864 11169
rect 21916 11160 21968 11212
rect 20904 11092 20956 11144
rect 22560 11092 22612 11144
rect 18512 11024 18564 11076
rect 15200 10956 15252 11008
rect 17500 10956 17552 11008
rect 17868 10956 17920 11008
rect 17960 10956 18012 11008
rect 18052 10956 18104 11008
rect 19616 10956 19668 11008
rect 21732 11024 21784 11076
rect 22284 11024 22336 11076
rect 22468 10956 22520 11008
rect 22928 11024 22980 11076
rect 23204 11092 23256 11144
rect 25688 11135 25740 11144
rect 25688 11101 25697 11135
rect 25697 11101 25731 11135
rect 25731 11101 25740 11135
rect 25688 11092 25740 11101
rect 25872 11135 25924 11144
rect 25872 11101 25881 11135
rect 25881 11101 25915 11135
rect 25915 11101 25924 11135
rect 25872 11092 25924 11101
rect 26700 11135 26752 11144
rect 23388 11024 23440 11076
rect 25504 11067 25556 11076
rect 23204 10956 23256 11008
rect 24400 10956 24452 11008
rect 25504 11033 25513 11067
rect 25513 11033 25547 11067
rect 25547 11033 25556 11067
rect 25504 11024 25556 11033
rect 26700 11101 26709 11135
rect 26709 11101 26743 11135
rect 26743 11101 26752 11135
rect 26700 11092 26752 11101
rect 26792 11092 26844 11144
rect 29644 11092 29696 11144
rect 29736 11135 29788 11144
rect 29736 11101 29745 11135
rect 29745 11101 29779 11135
rect 29779 11101 29788 11135
rect 29736 11092 29788 11101
rect 30196 11135 30248 11144
rect 27252 11024 27304 11076
rect 29276 11024 29328 11076
rect 29368 11024 29420 11076
rect 30196 11101 30205 11135
rect 30205 11101 30239 11135
rect 30239 11101 30248 11135
rect 30840 11135 30892 11144
rect 30196 11092 30248 11101
rect 30840 11101 30849 11135
rect 30849 11101 30883 11135
rect 30883 11101 30892 11135
rect 30840 11092 30892 11101
rect 30104 11024 30156 11076
rect 25964 10956 26016 11008
rect 29000 10956 29052 11008
rect 29644 10956 29696 11008
rect 7288 10854 7340 10906
rect 17592 10854 17644 10906
rect 27896 10854 27948 10906
rect 2872 10752 2924 10804
rect 6736 10795 6788 10804
rect 1860 10684 1912 10736
rect 4528 10684 4580 10736
rect 6736 10761 6745 10795
rect 6745 10761 6779 10795
rect 6779 10761 6788 10795
rect 6736 10752 6788 10761
rect 2044 10616 2096 10668
rect 2228 10659 2280 10668
rect 2228 10625 2237 10659
rect 2237 10625 2271 10659
rect 2271 10625 2280 10659
rect 2228 10616 2280 10625
rect 2320 10616 2372 10668
rect 7923 10727 7975 10736
rect 7923 10693 7931 10727
rect 7931 10693 7965 10727
rect 7965 10693 7975 10727
rect 7923 10684 7975 10693
rect 8576 10752 8628 10804
rect 15016 10752 15068 10804
rect 4988 10659 5040 10668
rect 1492 10548 1544 10600
rect 1768 10548 1820 10600
rect 3056 10548 3108 10600
rect 2780 10480 2832 10532
rect 4528 10548 4580 10600
rect 4988 10625 4997 10659
rect 4997 10625 5031 10659
rect 5031 10625 5040 10659
rect 4988 10616 5040 10625
rect 5632 10616 5684 10668
rect 6000 10616 6052 10668
rect 7012 10616 7064 10668
rect 7656 10616 7708 10668
rect 8116 10616 8168 10668
rect 10140 10684 10192 10736
rect 8576 10616 8628 10668
rect 9496 10659 9548 10668
rect 4804 10548 4856 10600
rect 7196 10591 7248 10600
rect 3608 10480 3660 10532
rect 7196 10557 7205 10591
rect 7205 10557 7239 10591
rect 7239 10557 7248 10591
rect 7196 10548 7248 10557
rect 6920 10480 6972 10532
rect 9496 10625 9505 10659
rect 9505 10625 9539 10659
rect 9539 10625 9548 10659
rect 9496 10616 9548 10625
rect 9864 10616 9916 10668
rect 12624 10684 12676 10736
rect 13360 10684 13412 10736
rect 15936 10684 15988 10736
rect 9680 10548 9732 10600
rect 10232 10548 10284 10600
rect 12992 10616 13044 10668
rect 14648 10616 14700 10668
rect 15200 10659 15252 10668
rect 11060 10548 11112 10600
rect 11888 10548 11940 10600
rect 15200 10625 15209 10659
rect 15209 10625 15243 10659
rect 15243 10625 15252 10659
rect 15200 10616 15252 10625
rect 16028 10659 16080 10668
rect 16028 10625 16037 10659
rect 16037 10625 16071 10659
rect 16071 10625 16080 10659
rect 16028 10616 16080 10625
rect 16120 10659 16172 10668
rect 16120 10625 16129 10659
rect 16129 10625 16163 10659
rect 16163 10625 16172 10659
rect 16120 10616 16172 10625
rect 17868 10752 17920 10804
rect 18420 10752 18472 10804
rect 20904 10752 20956 10804
rect 17960 10684 18012 10736
rect 19064 10684 19116 10736
rect 19432 10684 19484 10736
rect 16672 10591 16724 10600
rect 1768 10455 1820 10464
rect 1768 10421 1777 10455
rect 1777 10421 1811 10455
rect 1811 10421 1820 10455
rect 1768 10412 1820 10421
rect 4436 10412 4488 10464
rect 5080 10412 5132 10464
rect 5724 10412 5776 10464
rect 7748 10412 7800 10464
rect 9588 10480 9640 10532
rect 10324 10480 10376 10532
rect 14280 10480 14332 10532
rect 8668 10412 8720 10464
rect 11152 10412 11204 10464
rect 11520 10455 11572 10464
rect 11520 10421 11529 10455
rect 11529 10421 11563 10455
rect 11563 10421 11572 10455
rect 11520 10412 11572 10421
rect 11980 10412 12032 10464
rect 16672 10557 16681 10591
rect 16681 10557 16715 10591
rect 16715 10557 16724 10591
rect 16672 10548 16724 10557
rect 17500 10616 17552 10668
rect 20628 10684 20680 10736
rect 22100 10752 22152 10804
rect 22560 10752 22612 10804
rect 21180 10659 21232 10668
rect 21180 10625 21189 10659
rect 21189 10625 21223 10659
rect 21223 10625 21232 10659
rect 21180 10616 21232 10625
rect 22100 10616 22152 10668
rect 22284 10659 22336 10668
rect 22284 10625 22293 10659
rect 22293 10625 22327 10659
rect 22327 10625 22336 10659
rect 22468 10659 22520 10668
rect 22284 10616 22336 10625
rect 22468 10625 22477 10659
rect 22477 10625 22511 10659
rect 22511 10625 22520 10659
rect 22468 10616 22520 10625
rect 17684 10548 17736 10600
rect 19340 10548 19392 10600
rect 23204 10616 23256 10668
rect 23940 10752 23992 10804
rect 25688 10752 25740 10804
rect 26148 10752 26200 10804
rect 29828 10752 29880 10804
rect 30196 10752 30248 10804
rect 30840 10752 30892 10804
rect 24032 10684 24084 10736
rect 23112 10591 23164 10600
rect 23112 10557 23121 10591
rect 23121 10557 23155 10591
rect 23155 10557 23164 10591
rect 23112 10548 23164 10557
rect 23296 10548 23348 10600
rect 23756 10616 23808 10668
rect 23848 10616 23900 10668
rect 25964 10659 26016 10668
rect 25964 10625 25973 10659
rect 25973 10625 26007 10659
rect 26007 10625 26016 10659
rect 25964 10616 26016 10625
rect 26240 10616 26292 10668
rect 27252 10684 27304 10736
rect 29000 10727 29052 10736
rect 27436 10659 27488 10668
rect 27436 10625 27445 10659
rect 27445 10625 27479 10659
rect 27479 10625 27488 10659
rect 27436 10616 27488 10625
rect 29000 10693 29034 10727
rect 29034 10693 29052 10727
rect 29000 10684 29052 10693
rect 29184 10684 29236 10736
rect 29644 10684 29696 10736
rect 20444 10412 20496 10464
rect 24952 10480 25004 10532
rect 27528 10548 27580 10600
rect 29736 10616 29788 10668
rect 31208 10659 31260 10668
rect 31208 10625 31217 10659
rect 31217 10625 31251 10659
rect 31251 10625 31260 10659
rect 31208 10616 31260 10625
rect 26240 10480 26292 10532
rect 21548 10412 21600 10464
rect 21824 10455 21876 10464
rect 21824 10421 21833 10455
rect 21833 10421 21867 10455
rect 21867 10421 21876 10455
rect 21824 10412 21876 10421
rect 24216 10455 24268 10464
rect 24216 10421 24225 10455
rect 24225 10421 24259 10455
rect 24259 10421 24268 10455
rect 24216 10412 24268 10421
rect 25872 10412 25924 10464
rect 26332 10412 26384 10464
rect 2136 10310 2188 10362
rect 12440 10310 12492 10362
rect 22744 10310 22796 10362
rect 1124 10208 1176 10260
rect 3056 10208 3108 10260
rect 3884 10208 3936 10260
rect 5448 10208 5500 10260
rect 6460 10208 6512 10260
rect 6276 10140 6328 10192
rect 7656 10140 7708 10192
rect 8208 10251 8260 10260
rect 8208 10217 8217 10251
rect 8217 10217 8251 10251
rect 8251 10217 8260 10251
rect 8208 10208 8260 10217
rect 8944 10208 8996 10260
rect 11152 10251 11204 10260
rect 11152 10217 11161 10251
rect 11161 10217 11195 10251
rect 11195 10217 11204 10251
rect 11152 10208 11204 10217
rect 13084 10208 13136 10260
rect 16028 10208 16080 10260
rect 11244 10140 11296 10192
rect 16672 10140 16724 10192
rect 18328 10208 18380 10260
rect 23848 10208 23900 10260
rect 24032 10208 24084 10260
rect 25964 10208 26016 10260
rect 27252 10208 27304 10260
rect 31208 10251 31260 10260
rect 31208 10217 31217 10251
rect 31217 10217 31251 10251
rect 31251 10217 31260 10251
rect 31208 10208 31260 10217
rect 18512 10140 18564 10192
rect 9220 10072 9272 10124
rect 14280 10072 14332 10124
rect 2688 10004 2740 10056
rect 4160 10047 4212 10056
rect 4160 10013 4169 10047
rect 4169 10013 4203 10047
rect 4203 10013 4212 10047
rect 4160 10004 4212 10013
rect 6000 10004 6052 10056
rect 6736 10004 6788 10056
rect 7380 10047 7432 10056
rect 1768 9936 1820 9988
rect 7104 9936 7156 9988
rect 7380 10013 7389 10047
rect 7389 10013 7423 10047
rect 7423 10013 7432 10047
rect 7380 10004 7432 10013
rect 8392 9936 8444 9988
rect 8760 9936 8812 9988
rect 8944 9936 8996 9988
rect 11796 10047 11848 10056
rect 11796 10013 11805 10047
rect 11805 10013 11839 10047
rect 11839 10013 11848 10047
rect 11796 10004 11848 10013
rect 9864 9936 9916 9988
rect 11520 9936 11572 9988
rect 12072 9979 12124 9988
rect 12072 9945 12106 9979
rect 12106 9945 12124 9979
rect 14464 9979 14516 9988
rect 12072 9936 12124 9945
rect 14464 9945 14473 9979
rect 14473 9945 14507 9979
rect 14507 9945 14516 9979
rect 14464 9936 14516 9945
rect 2228 9868 2280 9920
rect 3424 9868 3476 9920
rect 3792 9868 3844 9920
rect 6000 9868 6052 9920
rect 7196 9868 7248 9920
rect 8300 9868 8352 9920
rect 8852 9868 8904 9920
rect 14096 9868 14148 9920
rect 18328 10004 18380 10056
rect 18604 10004 18656 10056
rect 21916 10140 21968 10192
rect 20812 10072 20864 10124
rect 21088 10004 21140 10056
rect 21640 10004 21692 10056
rect 19340 9979 19392 9988
rect 19340 9945 19349 9979
rect 19349 9945 19383 9979
rect 19383 9945 19392 9979
rect 19340 9936 19392 9945
rect 23664 10004 23716 10056
rect 26792 10004 26844 10056
rect 27528 10004 27580 10056
rect 29184 10004 29236 10056
rect 30104 10047 30156 10056
rect 30104 10013 30138 10047
rect 30138 10013 30156 10047
rect 30104 10004 30156 10013
rect 22652 9936 22704 9988
rect 23296 9936 23348 9988
rect 16120 9868 16172 9920
rect 19524 9868 19576 9920
rect 22468 9868 22520 9920
rect 23112 9868 23164 9920
rect 24216 9936 24268 9988
rect 26148 9936 26200 9988
rect 26240 9868 26292 9920
rect 28540 9868 28592 9920
rect 29092 9868 29144 9920
rect 7288 9766 7340 9818
rect 17592 9766 17644 9818
rect 27896 9766 27948 9818
rect 3700 9664 3752 9716
rect 3884 9664 3936 9716
rect 6644 9664 6696 9716
rect 7656 9664 7708 9716
rect 1768 9596 1820 9648
rect 2320 9596 2372 9648
rect 1400 9571 1452 9580
rect 1400 9537 1409 9571
rect 1409 9537 1443 9571
rect 1443 9537 1452 9571
rect 1400 9528 1452 9537
rect 2228 9528 2280 9580
rect 2688 9528 2740 9580
rect 4712 9596 4764 9648
rect 4896 9639 4948 9648
rect 4896 9605 4905 9639
rect 4905 9605 4939 9639
rect 4939 9605 4948 9639
rect 4896 9596 4948 9605
rect 4528 9528 4580 9580
rect 5080 9571 5132 9580
rect 5080 9537 5089 9571
rect 5089 9537 5123 9571
rect 5123 9537 5132 9571
rect 5080 9528 5132 9537
rect 2320 9503 2372 9512
rect 2320 9469 2329 9503
rect 2329 9469 2363 9503
rect 2363 9469 2372 9503
rect 2320 9460 2372 9469
rect 2412 9460 2464 9512
rect 5724 9528 5776 9580
rect 6552 9528 6604 9580
rect 6828 9596 6880 9648
rect 8024 9596 8076 9648
rect 8392 9596 8444 9648
rect 9036 9664 9088 9716
rect 9220 9664 9272 9716
rect 8668 9528 8720 9580
rect 7380 9503 7432 9512
rect 3608 9435 3660 9444
rect 3608 9401 3617 9435
rect 3617 9401 3651 9435
rect 3651 9401 3660 9435
rect 3608 9392 3660 9401
rect 3976 9392 4028 9444
rect 7380 9469 7389 9503
rect 7389 9469 7423 9503
rect 7423 9469 7432 9503
rect 7380 9460 7432 9469
rect 7564 9460 7616 9512
rect 8760 9460 8812 9512
rect 9588 9596 9640 9648
rect 13912 9596 13964 9648
rect 14372 9639 14424 9648
rect 14372 9605 14406 9639
rect 14406 9605 14424 9639
rect 14372 9596 14424 9605
rect 9680 9528 9732 9580
rect 10968 9537 10973 9564
rect 10973 9537 11007 9564
rect 11007 9537 11020 9564
rect 10968 9512 11020 9537
rect 11152 9528 11204 9580
rect 11612 9528 11664 9580
rect 11888 9528 11940 9580
rect 12164 9571 12216 9580
rect 12164 9537 12173 9571
rect 12173 9537 12207 9571
rect 12207 9537 12216 9571
rect 12164 9528 12216 9537
rect 12992 9528 13044 9580
rect 14096 9571 14148 9580
rect 14096 9537 14105 9571
rect 14105 9537 14139 9571
rect 14139 9537 14148 9571
rect 14096 9528 14148 9537
rect 21916 9596 21968 9648
rect 22652 9664 22704 9716
rect 26240 9664 26292 9716
rect 26424 9664 26476 9716
rect 26700 9664 26752 9716
rect 23020 9596 23072 9648
rect 24124 9596 24176 9648
rect 24860 9596 24912 9648
rect 25504 9596 25556 9648
rect 1952 9324 2004 9376
rect 6276 9324 6328 9376
rect 9036 9392 9088 9444
rect 7656 9324 7708 9376
rect 8576 9324 8628 9376
rect 10324 9460 10376 9512
rect 10876 9460 10928 9512
rect 14648 9528 14700 9580
rect 16120 9571 16172 9580
rect 16120 9537 16129 9571
rect 16129 9537 16163 9571
rect 16163 9537 16172 9571
rect 16120 9528 16172 9537
rect 16212 9528 16264 9580
rect 17500 9528 17552 9580
rect 17776 9528 17828 9580
rect 17868 9528 17920 9580
rect 18420 9571 18472 9580
rect 18420 9537 18429 9571
rect 18429 9537 18463 9571
rect 18463 9537 18472 9571
rect 18420 9528 18472 9537
rect 9680 9392 9732 9444
rect 18144 9503 18196 9512
rect 14004 9392 14056 9444
rect 15108 9392 15160 9444
rect 18144 9469 18153 9503
rect 18153 9469 18187 9503
rect 18187 9469 18196 9503
rect 18144 9460 18196 9469
rect 18512 9460 18564 9512
rect 9496 9324 9548 9376
rect 10600 9324 10652 9376
rect 11244 9324 11296 9376
rect 11980 9324 12032 9376
rect 13084 9324 13136 9376
rect 15752 9324 15804 9376
rect 17776 9392 17828 9444
rect 19340 9528 19392 9580
rect 18696 9460 18748 9512
rect 19156 9460 19208 9512
rect 20260 9460 20312 9512
rect 20536 9528 20588 9580
rect 21272 9528 21324 9580
rect 21824 9528 21876 9580
rect 22468 9528 22520 9580
rect 22100 9460 22152 9512
rect 23296 9528 23348 9580
rect 25044 9528 25096 9580
rect 25596 9528 25648 9580
rect 25780 9528 25832 9580
rect 29092 9596 29144 9648
rect 27712 9528 27764 9580
rect 29276 9528 29328 9580
rect 30012 9528 30064 9580
rect 29644 9460 29696 9512
rect 19064 9392 19116 9444
rect 19524 9392 19576 9444
rect 20628 9392 20680 9444
rect 21732 9392 21784 9444
rect 22928 9392 22980 9444
rect 23572 9392 23624 9444
rect 16304 9324 16356 9376
rect 17040 9367 17092 9376
rect 17040 9333 17049 9367
rect 17049 9333 17083 9367
rect 17083 9333 17092 9367
rect 17040 9324 17092 9333
rect 17960 9367 18012 9376
rect 17960 9333 17969 9367
rect 17969 9333 18003 9367
rect 18003 9333 18012 9367
rect 17960 9324 18012 9333
rect 18144 9324 18196 9376
rect 19616 9324 19668 9376
rect 23204 9324 23256 9376
rect 23296 9324 23348 9376
rect 23756 9324 23808 9376
rect 24124 9324 24176 9376
rect 25964 9324 26016 9376
rect 28632 9392 28684 9444
rect 30932 9392 30984 9444
rect 28356 9324 28408 9376
rect 29000 9367 29052 9376
rect 29000 9333 29009 9367
rect 29009 9333 29043 9367
rect 29043 9333 29052 9367
rect 29000 9324 29052 9333
rect 31116 9367 31168 9376
rect 31116 9333 31125 9367
rect 31125 9333 31159 9367
rect 31159 9333 31168 9367
rect 31116 9324 31168 9333
rect 2136 9222 2188 9274
rect 12440 9222 12492 9274
rect 22744 9222 22796 9274
rect 3332 9120 3384 9172
rect 3884 9120 3936 9172
rect 7564 9120 7616 9172
rect 2596 9052 2648 9104
rect 9680 9052 9732 9104
rect 11520 9052 11572 9104
rect 12164 9052 12216 9104
rect 13084 9052 13136 9104
rect 14004 9120 14056 9172
rect 17776 9120 17828 9172
rect 17960 9120 18012 9172
rect 24952 9120 25004 9172
rect 26148 9163 26200 9172
rect 26148 9129 26157 9163
rect 26157 9129 26191 9163
rect 26191 9129 26200 9163
rect 26148 9120 26200 9129
rect 27712 9120 27764 9172
rect 28264 9120 28316 9172
rect 28356 9120 28408 9172
rect 14372 9052 14424 9104
rect 18236 9052 18288 9104
rect 2228 8984 2280 9036
rect 5632 8984 5684 9036
rect 8116 8984 8168 9036
rect 12716 8984 12768 9036
rect 13544 8984 13596 9036
rect 14096 8984 14148 9036
rect 15936 8984 15988 9036
rect 19708 9052 19760 9104
rect 21272 9052 21324 9104
rect 1676 8916 1728 8968
rect 3240 8916 3292 8968
rect 4896 8916 4948 8968
rect 5264 8959 5316 8968
rect 5264 8925 5273 8959
rect 5273 8925 5307 8959
rect 5307 8925 5316 8959
rect 5264 8916 5316 8925
rect 5448 8959 5500 8968
rect 5448 8925 5457 8959
rect 5457 8925 5491 8959
rect 5491 8925 5500 8959
rect 5448 8916 5500 8925
rect 4068 8848 4120 8900
rect 6276 8959 6328 8968
rect 6276 8925 6285 8959
rect 6285 8925 6319 8959
rect 6319 8925 6328 8959
rect 6920 8959 6972 8968
rect 6276 8916 6328 8925
rect 6920 8925 6929 8959
rect 6929 8925 6963 8959
rect 6963 8925 6972 8959
rect 6920 8916 6972 8925
rect 7104 8916 7156 8968
rect 9220 8959 9272 8968
rect 9220 8925 9229 8959
rect 9229 8925 9263 8959
rect 9263 8925 9272 8959
rect 9220 8916 9272 8925
rect 6000 8848 6052 8900
rect 6644 8848 6696 8900
rect 1952 8823 2004 8832
rect 1952 8789 1961 8823
rect 1961 8789 1995 8823
rect 1995 8789 2004 8823
rect 1952 8780 2004 8789
rect 3056 8780 3108 8832
rect 4344 8823 4396 8832
rect 4344 8789 4353 8823
rect 4353 8789 4387 8823
rect 4387 8789 4396 8823
rect 4344 8780 4396 8789
rect 7472 8780 7524 8832
rect 8024 8780 8076 8832
rect 8300 8848 8352 8900
rect 9588 8916 9640 8968
rect 10600 8916 10652 8968
rect 16304 8916 16356 8968
rect 16580 8916 16632 8968
rect 17040 8916 17092 8968
rect 17500 8916 17552 8968
rect 17868 8916 17920 8968
rect 18236 8959 18288 8968
rect 18236 8925 18245 8959
rect 18245 8925 18279 8959
rect 18279 8925 18288 8959
rect 18236 8916 18288 8925
rect 18512 8959 18564 8968
rect 18512 8925 18521 8959
rect 18521 8925 18555 8959
rect 18555 8925 18564 8959
rect 19616 8984 19668 9036
rect 21548 8984 21600 9036
rect 21824 8984 21876 9036
rect 22468 9052 22520 9104
rect 23204 9052 23256 9104
rect 25872 9052 25924 9104
rect 28080 9052 28132 9104
rect 29276 9052 29328 9104
rect 18512 8916 18564 8925
rect 19708 8959 19760 8968
rect 19708 8925 19717 8959
rect 19717 8925 19751 8959
rect 19751 8925 19760 8959
rect 19708 8916 19760 8925
rect 20168 8916 20220 8968
rect 21088 8916 21140 8968
rect 23204 8916 23256 8968
rect 11704 8848 11756 8900
rect 8484 8780 8536 8832
rect 18144 8848 18196 8900
rect 22284 8891 22336 8900
rect 22284 8857 22293 8891
rect 22293 8857 22327 8891
rect 22327 8857 22336 8891
rect 22284 8848 22336 8857
rect 22652 8891 22704 8900
rect 22652 8857 22661 8891
rect 22661 8857 22695 8891
rect 22695 8857 22704 8891
rect 22652 8848 22704 8857
rect 24860 8848 24912 8900
rect 26332 8959 26384 8968
rect 26332 8925 26341 8959
rect 26341 8925 26375 8959
rect 26375 8925 26384 8959
rect 26332 8916 26384 8925
rect 28540 8959 28592 8968
rect 28540 8925 28549 8959
rect 28549 8925 28583 8959
rect 28583 8925 28592 8959
rect 28540 8916 28592 8925
rect 29644 8984 29696 9036
rect 29000 8959 29052 8968
rect 29000 8925 29009 8959
rect 29009 8925 29043 8959
rect 29043 8925 29052 8959
rect 29000 8916 29052 8925
rect 13636 8780 13688 8832
rect 13912 8780 13964 8832
rect 15752 8780 15804 8832
rect 15936 8780 15988 8832
rect 16488 8823 16540 8832
rect 16488 8789 16497 8823
rect 16497 8789 16531 8823
rect 16531 8789 16540 8823
rect 16488 8780 16540 8789
rect 18328 8780 18380 8832
rect 19432 8780 19484 8832
rect 19984 8780 20036 8832
rect 20720 8780 20772 8832
rect 23020 8823 23072 8832
rect 23020 8789 23029 8823
rect 23029 8789 23063 8823
rect 23063 8789 23072 8823
rect 23020 8780 23072 8789
rect 23756 8780 23808 8832
rect 25044 8780 25096 8832
rect 25964 8780 26016 8832
rect 27344 8780 27396 8832
rect 30380 8848 30432 8900
rect 30932 8916 30984 8968
rect 31300 8959 31352 8968
rect 31300 8925 31309 8959
rect 31309 8925 31343 8959
rect 31343 8925 31352 8959
rect 31300 8916 31352 8925
rect 31392 8848 31444 8900
rect 29828 8780 29880 8832
rect 30656 8780 30708 8832
rect 7288 8678 7340 8730
rect 17592 8678 17644 8730
rect 27896 8678 27948 8730
rect 4344 8576 4396 8628
rect 5540 8619 5592 8628
rect 5540 8585 5549 8619
rect 5549 8585 5583 8619
rect 5583 8585 5592 8619
rect 5540 8576 5592 8585
rect 1952 8508 2004 8560
rect 1768 8440 1820 8492
rect 3608 8508 3660 8560
rect 6920 8576 6972 8628
rect 8300 8576 8352 8628
rect 8576 8619 8628 8628
rect 8576 8585 8585 8619
rect 8585 8585 8619 8619
rect 8619 8585 8628 8619
rect 8576 8576 8628 8585
rect 8668 8576 8720 8628
rect 19294 8576 19346 8628
rect 19984 8576 20036 8628
rect 31116 8576 31168 8628
rect 3332 8440 3384 8492
rect 3976 8440 4028 8492
rect 4160 8483 4212 8492
rect 4160 8449 4169 8483
rect 4169 8449 4203 8483
rect 4203 8449 4212 8483
rect 4160 8440 4212 8449
rect 6276 8440 6328 8492
rect 6460 8440 6512 8492
rect 9680 8508 9732 8560
rect 9864 8508 9916 8560
rect 8944 8440 8996 8492
rect 10600 8483 10652 8492
rect 10600 8449 10609 8483
rect 10609 8449 10643 8483
rect 10643 8449 10652 8483
rect 10600 8440 10652 8449
rect 10784 8508 10836 8560
rect 14096 8508 14148 8560
rect 16488 8508 16540 8560
rect 17040 8508 17092 8560
rect 17500 8508 17552 8560
rect 18696 8508 18748 8560
rect 18880 8508 18932 8560
rect 22560 8508 22612 8560
rect 15660 8440 15712 8492
rect 2320 8372 2372 8424
rect 3240 8415 3292 8424
rect 2412 8304 2464 8356
rect 3240 8381 3249 8415
rect 3249 8381 3283 8415
rect 3283 8381 3292 8415
rect 3240 8372 3292 8381
rect 6000 8372 6052 8424
rect 8208 8372 8260 8424
rect 10968 8372 11020 8424
rect 3976 8304 4028 8356
rect 7656 8304 7708 8356
rect 9312 8304 9364 8356
rect 2596 8279 2648 8288
rect 2596 8245 2605 8279
rect 2605 8245 2639 8279
rect 2639 8245 2648 8279
rect 2596 8236 2648 8245
rect 2688 8236 2740 8288
rect 4896 8236 4948 8288
rect 5080 8236 5132 8288
rect 6644 8236 6696 8288
rect 9128 8236 9180 8288
rect 10508 8304 10560 8356
rect 11244 8372 11296 8424
rect 9772 8279 9824 8288
rect 9772 8245 9781 8279
rect 9781 8245 9815 8279
rect 9815 8245 9824 8279
rect 9772 8236 9824 8245
rect 10140 8236 10192 8288
rect 14372 8347 14424 8356
rect 13360 8236 13412 8288
rect 14372 8313 14381 8347
rect 14381 8313 14415 8347
rect 14415 8313 14424 8347
rect 14372 8304 14424 8313
rect 14648 8304 14700 8356
rect 15384 8372 15436 8424
rect 18236 8440 18288 8492
rect 19156 8483 19208 8492
rect 19156 8449 19165 8483
rect 19165 8449 19199 8483
rect 19199 8449 19208 8483
rect 19156 8440 19208 8449
rect 16672 8415 16724 8424
rect 16672 8381 16681 8415
rect 16681 8381 16715 8415
rect 16715 8381 16724 8415
rect 16672 8372 16724 8381
rect 19800 8440 19852 8492
rect 20260 8483 20312 8492
rect 20260 8449 20269 8483
rect 20269 8449 20303 8483
rect 20303 8449 20312 8483
rect 20260 8440 20312 8449
rect 20536 8483 20588 8492
rect 20536 8449 20545 8483
rect 20545 8449 20579 8483
rect 20579 8449 20588 8483
rect 20536 8440 20588 8449
rect 20720 8483 20772 8492
rect 20720 8449 20729 8483
rect 20729 8449 20763 8483
rect 20763 8449 20772 8483
rect 20720 8440 20772 8449
rect 21732 8440 21784 8492
rect 23020 8508 23072 8560
rect 25044 8508 25096 8560
rect 25136 8508 25188 8560
rect 23112 8440 23164 8492
rect 23204 8440 23256 8492
rect 24400 8440 24452 8492
rect 25228 8483 25280 8492
rect 25228 8449 25237 8483
rect 25237 8449 25271 8483
rect 25271 8449 25280 8483
rect 25228 8440 25280 8449
rect 26056 8508 26108 8560
rect 27804 8508 27856 8560
rect 27620 8440 27672 8492
rect 29736 8440 29788 8492
rect 31024 8483 31076 8492
rect 31024 8449 31033 8483
rect 31033 8449 31067 8483
rect 31067 8449 31076 8483
rect 31024 8440 31076 8449
rect 17960 8304 18012 8356
rect 18512 8304 18564 8356
rect 19616 8304 19668 8356
rect 22560 8372 22612 8424
rect 22836 8415 22888 8424
rect 22836 8381 22845 8415
rect 22845 8381 22879 8415
rect 22879 8381 22888 8415
rect 22836 8372 22888 8381
rect 20628 8304 20680 8356
rect 25780 8372 25832 8424
rect 27344 8372 27396 8424
rect 31300 8415 31352 8424
rect 23756 8304 23808 8356
rect 24584 8304 24636 8356
rect 26608 8304 26660 8356
rect 27528 8304 27580 8356
rect 28264 8304 28316 8356
rect 30196 8304 30248 8356
rect 31300 8381 31309 8415
rect 31309 8381 31343 8415
rect 31343 8381 31352 8415
rect 31300 8372 31352 8381
rect 31392 8304 31444 8356
rect 22284 8236 22336 8288
rect 23296 8236 23348 8288
rect 24492 8236 24544 8288
rect 25596 8279 25648 8288
rect 25596 8245 25605 8279
rect 25605 8245 25639 8279
rect 25639 8245 25648 8279
rect 25596 8236 25648 8245
rect 27252 8236 27304 8288
rect 27988 8236 28040 8288
rect 29092 8236 29144 8288
rect 29644 8236 29696 8288
rect 2136 8134 2188 8186
rect 12440 8134 12492 8186
rect 22744 8134 22796 8186
rect 2688 8032 2740 8084
rect 6460 8032 6512 8084
rect 8208 8075 8260 8084
rect 8208 8041 8217 8075
rect 8217 8041 8251 8075
rect 8251 8041 8260 8075
rect 8208 8032 8260 8041
rect 9220 8032 9272 8084
rect 10600 8032 10652 8084
rect 13452 8075 13504 8084
rect 13452 8041 13461 8075
rect 13461 8041 13495 8075
rect 13495 8041 13504 8075
rect 13452 8032 13504 8041
rect 16212 8032 16264 8084
rect 16856 8032 16908 8084
rect 17224 8032 17276 8084
rect 18788 8032 18840 8084
rect 20720 8075 20772 8084
rect 20720 8041 20729 8075
rect 20729 8041 20763 8075
rect 20763 8041 20772 8075
rect 21640 8075 21692 8084
rect 20720 8032 20772 8041
rect 21640 8041 21649 8075
rect 21649 8041 21683 8075
rect 21683 8041 21692 8075
rect 21640 8032 21692 8041
rect 21732 8032 21784 8084
rect 22376 8032 22428 8084
rect 1400 7896 1452 7948
rect 2412 7896 2464 7948
rect 1768 7828 1820 7880
rect 2228 7871 2280 7880
rect 2228 7837 2237 7871
rect 2237 7837 2271 7871
rect 2271 7837 2280 7871
rect 2228 7828 2280 7837
rect 2504 7871 2556 7880
rect 2504 7837 2513 7871
rect 2513 7837 2547 7871
rect 2547 7837 2556 7871
rect 2504 7828 2556 7837
rect 3056 7896 3108 7948
rect 6184 7964 6236 8016
rect 8024 8007 8076 8016
rect 8024 7973 8033 8007
rect 8033 7973 8067 8007
rect 8067 7973 8076 8007
rect 8024 7964 8076 7973
rect 10232 7964 10284 8016
rect 11612 7964 11664 8016
rect 12624 7964 12676 8016
rect 16028 7964 16080 8016
rect 5080 7896 5132 7948
rect 3608 7760 3660 7812
rect 4804 7828 4856 7880
rect 5264 7896 5316 7948
rect 5448 7896 5500 7948
rect 5540 7828 5592 7880
rect 6736 7896 6788 7948
rect 7104 7828 7156 7880
rect 7380 7896 7432 7948
rect 9772 7896 9824 7948
rect 9128 7871 9180 7880
rect 9128 7837 9137 7871
rect 9137 7837 9171 7871
rect 9171 7837 9180 7871
rect 9128 7828 9180 7837
rect 6920 7760 6972 7812
rect 9036 7760 9088 7812
rect 9680 7828 9732 7880
rect 10416 7828 10468 7880
rect 10968 7828 11020 7880
rect 11704 7828 11756 7880
rect 10784 7760 10836 7812
rect 16304 7896 16356 7948
rect 21916 7896 21968 7948
rect 29276 8032 29328 8084
rect 12532 7871 12584 7880
rect 12532 7837 12541 7871
rect 12541 7837 12575 7871
rect 12575 7837 12584 7871
rect 12532 7828 12584 7837
rect 12808 7871 12860 7880
rect 12808 7837 12817 7871
rect 12817 7837 12851 7871
rect 12851 7837 12860 7871
rect 12808 7828 12860 7837
rect 14096 7871 14148 7880
rect 14096 7837 14105 7871
rect 14105 7837 14139 7871
rect 14139 7837 14148 7871
rect 14096 7828 14148 7837
rect 14280 7828 14332 7880
rect 14740 7828 14792 7880
rect 15108 7828 15160 7880
rect 15016 7760 15068 7812
rect 15936 7828 15988 7880
rect 16672 7828 16724 7880
rect 17684 7828 17736 7880
rect 20168 7828 20220 7880
rect 21272 7871 21324 7880
rect 21272 7837 21281 7871
rect 21281 7837 21315 7871
rect 21315 7837 21324 7871
rect 21272 7828 21324 7837
rect 22008 7828 22060 7880
rect 22100 7828 22152 7880
rect 24124 7828 24176 7880
rect 24952 7871 25004 7880
rect 24952 7837 24961 7871
rect 24961 7837 24995 7871
rect 24995 7837 25004 7871
rect 24952 7828 25004 7837
rect 25596 7871 25648 7880
rect 25596 7837 25605 7871
rect 25605 7837 25639 7871
rect 25639 7837 25648 7871
rect 25596 7828 25648 7837
rect 26976 7896 27028 7948
rect 31300 8032 31352 8084
rect 27344 7871 27396 7880
rect 27344 7837 27353 7871
rect 27353 7837 27387 7871
rect 27387 7837 27396 7871
rect 27344 7828 27396 7837
rect 28080 7871 28132 7880
rect 28080 7837 28089 7871
rect 28089 7837 28123 7871
rect 28123 7837 28132 7871
rect 28356 7871 28408 7880
rect 28080 7828 28132 7837
rect 28356 7837 28365 7871
rect 28365 7837 28399 7871
rect 28399 7837 28408 7871
rect 28356 7828 28408 7837
rect 29644 7828 29696 7880
rect 29828 7871 29880 7880
rect 29828 7837 29862 7871
rect 29862 7837 29880 7871
rect 29828 7828 29880 7837
rect 16948 7760 17000 7812
rect 17500 7760 17552 7812
rect 19432 7760 19484 7812
rect 21824 7760 21876 7812
rect 26148 7760 26200 7812
rect 1952 7692 2004 7744
rect 6552 7692 6604 7744
rect 10416 7692 10468 7744
rect 12348 7735 12400 7744
rect 12348 7701 12357 7735
rect 12357 7701 12391 7735
rect 12391 7701 12400 7735
rect 12348 7692 12400 7701
rect 13544 7692 13596 7744
rect 16856 7692 16908 7744
rect 21088 7692 21140 7744
rect 23664 7692 23716 7744
rect 25780 7692 25832 7744
rect 26700 7735 26752 7744
rect 26700 7701 26709 7735
rect 26709 7701 26743 7735
rect 26743 7701 26752 7735
rect 26700 7692 26752 7701
rect 28080 7692 28132 7744
rect 29000 7735 29052 7744
rect 29000 7701 29009 7735
rect 29009 7701 29043 7735
rect 29043 7701 29052 7735
rect 29000 7692 29052 7701
rect 31208 7692 31260 7744
rect 7288 7590 7340 7642
rect 17592 7590 17644 7642
rect 27896 7590 27948 7642
rect 2044 7531 2096 7540
rect 2044 7497 2053 7531
rect 2053 7497 2087 7531
rect 2087 7497 2096 7531
rect 2044 7488 2096 7497
rect 3976 7488 4028 7540
rect 5264 7488 5316 7540
rect 5356 7488 5408 7540
rect 5632 7488 5684 7540
rect 6000 7488 6052 7540
rect 6276 7488 6328 7540
rect 8760 7531 8812 7540
rect 8760 7497 8769 7531
rect 8769 7497 8803 7531
rect 8803 7497 8812 7531
rect 8760 7488 8812 7497
rect 10048 7488 10100 7540
rect 10784 7488 10836 7540
rect 10968 7531 11020 7540
rect 10968 7497 10977 7531
rect 10977 7497 11011 7531
rect 11011 7497 11020 7531
rect 10968 7488 11020 7497
rect 12532 7488 12584 7540
rect 15660 7531 15712 7540
rect 15660 7497 15669 7531
rect 15669 7497 15703 7531
rect 15703 7497 15712 7531
rect 15660 7488 15712 7497
rect 16580 7488 16632 7540
rect 21824 7488 21876 7540
rect 1768 7352 1820 7404
rect 2228 7395 2280 7404
rect 2228 7361 2237 7395
rect 2237 7361 2271 7395
rect 2271 7361 2280 7395
rect 2228 7352 2280 7361
rect 2504 7395 2556 7404
rect 2504 7361 2513 7395
rect 2513 7361 2547 7395
rect 2547 7361 2556 7395
rect 2504 7352 2556 7361
rect 2688 7395 2740 7404
rect 2688 7361 2697 7395
rect 2697 7361 2731 7395
rect 2731 7361 2740 7395
rect 2688 7352 2740 7361
rect 2320 7284 2372 7336
rect 3608 7352 3660 7404
rect 4804 7420 4856 7472
rect 4528 7352 4580 7404
rect 4988 7284 5040 7336
rect 5448 7352 5500 7404
rect 5816 7395 5868 7404
rect 5816 7361 5825 7395
rect 5825 7361 5859 7395
rect 5859 7361 5868 7395
rect 5816 7352 5868 7361
rect 6552 7395 6604 7404
rect 6552 7361 6561 7395
rect 6561 7361 6595 7395
rect 6595 7361 6604 7395
rect 6552 7352 6604 7361
rect 6644 7352 6696 7404
rect 8116 7420 8168 7472
rect 9956 7420 10008 7472
rect 11336 7420 11388 7472
rect 6920 7284 6972 7336
rect 6000 7216 6052 7268
rect 7196 7216 7248 7268
rect 2228 7148 2280 7200
rect 3976 7148 4028 7200
rect 5172 7191 5224 7200
rect 5172 7157 5181 7191
rect 5181 7157 5215 7191
rect 5215 7157 5224 7191
rect 5172 7148 5224 7157
rect 5264 7148 5316 7200
rect 6092 7148 6144 7200
rect 9404 7148 9456 7200
rect 10232 7352 10284 7404
rect 10324 7352 10376 7404
rect 11520 7352 11572 7404
rect 12348 7420 12400 7472
rect 13820 7352 13872 7404
rect 14004 7420 14056 7472
rect 14280 7352 14332 7404
rect 14740 7395 14792 7404
rect 14740 7361 14749 7395
rect 14749 7361 14783 7395
rect 14783 7361 14792 7395
rect 14740 7352 14792 7361
rect 15016 7395 15068 7404
rect 15016 7361 15025 7395
rect 15025 7361 15059 7395
rect 15059 7361 15068 7395
rect 15016 7352 15068 7361
rect 15476 7352 15528 7404
rect 16028 7395 16080 7404
rect 16028 7361 16037 7395
rect 16037 7361 16071 7395
rect 16071 7361 16080 7395
rect 16028 7352 16080 7361
rect 15384 7284 15436 7336
rect 13820 7216 13872 7268
rect 15108 7216 15160 7268
rect 16948 7352 17000 7404
rect 17960 7420 18012 7472
rect 18696 7420 18748 7472
rect 17684 7352 17736 7404
rect 18144 7352 18196 7404
rect 18328 7395 18380 7404
rect 18328 7361 18362 7395
rect 18362 7361 18380 7395
rect 18328 7352 18380 7361
rect 20628 7352 20680 7404
rect 19616 7284 19668 7336
rect 19156 7216 19208 7268
rect 20996 7284 21048 7336
rect 21364 7420 21416 7472
rect 22836 7488 22888 7540
rect 26148 7488 26200 7540
rect 23388 7420 23440 7472
rect 26976 7463 27028 7472
rect 22652 7352 22704 7404
rect 23664 7395 23716 7404
rect 23664 7361 23673 7395
rect 23673 7361 23707 7395
rect 23707 7361 23716 7395
rect 23664 7352 23716 7361
rect 23756 7395 23808 7404
rect 23756 7361 23765 7395
rect 23765 7361 23799 7395
rect 23799 7361 23808 7395
rect 23756 7352 23808 7361
rect 21640 7284 21692 7336
rect 22192 7284 22244 7336
rect 22376 7284 22428 7336
rect 23296 7284 23348 7336
rect 25136 7352 25188 7404
rect 24492 7327 24544 7336
rect 24492 7293 24501 7327
rect 24501 7293 24535 7327
rect 24535 7293 24544 7327
rect 24492 7284 24544 7293
rect 26976 7429 26985 7463
rect 26985 7429 27019 7463
rect 27019 7429 27028 7463
rect 26976 7420 27028 7429
rect 26056 7395 26108 7404
rect 26056 7361 26065 7395
rect 26065 7361 26099 7395
rect 26099 7361 26108 7395
rect 26056 7352 26108 7361
rect 26424 7352 26476 7404
rect 27068 7284 27120 7336
rect 27436 7284 27488 7336
rect 28356 7488 28408 7540
rect 29276 7531 29328 7540
rect 29276 7497 29285 7531
rect 29285 7497 29319 7531
rect 29319 7497 29328 7531
rect 29276 7488 29328 7497
rect 30288 7488 30340 7540
rect 31208 7488 31260 7540
rect 29644 7420 29696 7472
rect 30196 7463 30248 7472
rect 30196 7429 30230 7463
rect 30230 7429 30248 7463
rect 30196 7420 30248 7429
rect 27988 7352 28040 7404
rect 29644 7284 29696 7336
rect 29920 7327 29972 7336
rect 29920 7293 29929 7327
rect 29929 7293 29963 7327
rect 29963 7293 29972 7327
rect 29920 7284 29972 7293
rect 10324 7148 10376 7200
rect 10600 7148 10652 7200
rect 12900 7148 12952 7200
rect 13452 7191 13504 7200
rect 13452 7157 13461 7191
rect 13461 7157 13495 7191
rect 13495 7157 13504 7191
rect 13452 7148 13504 7157
rect 14740 7148 14792 7200
rect 15936 7148 15988 7200
rect 16304 7148 16356 7200
rect 19248 7148 19300 7200
rect 19800 7148 19852 7200
rect 20904 7148 20956 7200
rect 21640 7148 21692 7200
rect 25504 7148 25556 7200
rect 27528 7148 27580 7200
rect 27620 7148 27672 7200
rect 28172 7148 28224 7200
rect 2136 7046 2188 7098
rect 12440 7046 12492 7098
rect 22744 7046 22796 7098
rect 1308 6944 1360 6996
rect 3608 6944 3660 6996
rect 4068 6944 4120 6996
rect 5540 6944 5592 6996
rect 8116 6987 8168 6996
rect 8116 6953 8125 6987
rect 8125 6953 8159 6987
rect 8159 6953 8168 6987
rect 8116 6944 8168 6953
rect 10232 6987 10284 6996
rect 10232 6953 10241 6987
rect 10241 6953 10275 6987
rect 10275 6953 10284 6987
rect 10232 6944 10284 6953
rect 12900 6944 12952 6996
rect 2412 6876 2464 6928
rect 4620 6876 4672 6928
rect 4804 6876 4856 6928
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 3976 6783 4028 6792
rect 3976 6749 3985 6783
rect 3985 6749 4019 6783
rect 4019 6749 4028 6783
rect 3976 6740 4028 6749
rect 4344 6808 4396 6860
rect 10600 6876 10652 6928
rect 12808 6876 12860 6928
rect 14280 6876 14332 6928
rect 17132 6944 17184 6996
rect 17776 6944 17828 6996
rect 19432 6944 19484 6996
rect 21640 6987 21692 6996
rect 21640 6953 21649 6987
rect 21649 6953 21683 6987
rect 21683 6953 21692 6987
rect 21640 6944 21692 6953
rect 22284 6944 22336 6996
rect 22652 6944 22704 6996
rect 23204 6944 23256 6996
rect 24492 6944 24544 6996
rect 25964 6944 26016 6996
rect 27344 6944 27396 6996
rect 8760 6808 8812 6860
rect 9772 6808 9824 6860
rect 11336 6851 11388 6860
rect 11336 6817 11345 6851
rect 11345 6817 11379 6851
rect 11379 6817 11388 6851
rect 11336 6808 11388 6817
rect 4620 6740 4672 6792
rect 5264 6740 5316 6792
rect 5448 6740 5500 6792
rect 1768 6672 1820 6724
rect 2320 6672 2372 6724
rect 10232 6740 10284 6792
rect 10416 6783 10468 6792
rect 10416 6749 10425 6783
rect 10425 6749 10459 6783
rect 10459 6749 10468 6783
rect 10416 6740 10468 6749
rect 10600 6783 10652 6792
rect 10600 6749 10609 6783
rect 10609 6749 10643 6783
rect 10643 6749 10652 6783
rect 10600 6740 10652 6749
rect 11980 6740 12032 6792
rect 13084 6740 13136 6792
rect 14464 6808 14516 6860
rect 14740 6808 14792 6860
rect 15016 6851 15068 6860
rect 15016 6817 15025 6851
rect 15025 6817 15059 6851
rect 15059 6817 15068 6851
rect 15016 6808 15068 6817
rect 15384 6851 15436 6860
rect 15384 6817 15418 6851
rect 15418 6817 15436 6851
rect 15384 6808 15436 6817
rect 15752 6808 15804 6860
rect 19708 6851 19760 6860
rect 19708 6817 19717 6851
rect 19717 6817 19751 6851
rect 19751 6817 19760 6851
rect 19708 6808 19760 6817
rect 22928 6808 22980 6860
rect 25504 6851 25556 6860
rect 14372 6783 14424 6792
rect 6644 6715 6696 6724
rect 3056 6604 3108 6656
rect 3884 6604 3936 6656
rect 6644 6681 6653 6715
rect 6653 6681 6687 6715
rect 6687 6681 6696 6715
rect 6644 6672 6696 6681
rect 4252 6604 4304 6656
rect 7380 6604 7432 6656
rect 12256 6672 12308 6724
rect 11888 6604 11940 6656
rect 14372 6749 14381 6783
rect 14381 6749 14415 6783
rect 14415 6749 14424 6783
rect 14372 6740 14424 6749
rect 16488 6740 16540 6792
rect 16948 6783 17000 6792
rect 16948 6749 16957 6783
rect 16957 6749 16991 6783
rect 16991 6749 17000 6783
rect 16948 6740 17000 6749
rect 17132 6783 17184 6792
rect 17132 6749 17141 6783
rect 17141 6749 17175 6783
rect 17175 6749 17184 6783
rect 17132 6740 17184 6749
rect 15844 6604 15896 6656
rect 16028 6604 16080 6656
rect 16580 6672 16632 6724
rect 17316 6740 17368 6792
rect 17684 6740 17736 6792
rect 17868 6783 17920 6792
rect 17868 6749 17877 6783
rect 17877 6749 17911 6783
rect 17911 6749 17920 6783
rect 17868 6740 17920 6749
rect 17960 6740 18012 6792
rect 19524 6783 19576 6792
rect 19524 6749 19533 6783
rect 19533 6749 19567 6783
rect 19567 6749 19576 6783
rect 19524 6740 19576 6749
rect 19800 6783 19852 6792
rect 19800 6749 19809 6783
rect 19809 6749 19843 6783
rect 19843 6749 19852 6783
rect 19800 6740 19852 6749
rect 22100 6740 22152 6792
rect 23296 6740 23348 6792
rect 24584 6783 24636 6792
rect 24584 6749 24593 6783
rect 24593 6749 24627 6783
rect 24627 6749 24636 6783
rect 24584 6740 24636 6749
rect 25504 6817 25513 6851
rect 25513 6817 25547 6851
rect 25547 6817 25556 6851
rect 25504 6808 25556 6817
rect 27068 6808 27120 6860
rect 28264 6808 28316 6860
rect 29736 6851 29788 6860
rect 29736 6817 29745 6851
rect 29745 6817 29779 6851
rect 29779 6817 29788 6851
rect 29736 6808 29788 6817
rect 27252 6740 27304 6792
rect 27988 6740 28040 6792
rect 30748 6808 30800 6860
rect 31116 6808 31168 6860
rect 19892 6672 19944 6724
rect 21824 6672 21876 6724
rect 21088 6604 21140 6656
rect 22836 6604 22888 6656
rect 25044 6647 25096 6656
rect 25044 6613 25053 6647
rect 25053 6613 25087 6647
rect 25087 6613 25096 6647
rect 25044 6604 25096 6613
rect 29000 6672 29052 6724
rect 30288 6740 30340 6792
rect 30564 6740 30616 6792
rect 31392 6740 31444 6792
rect 30472 6672 30524 6724
rect 27712 6604 27764 6656
rect 30196 6604 30248 6656
rect 7288 6502 7340 6554
rect 17592 6502 17644 6554
rect 27896 6502 27948 6554
rect 1768 6443 1820 6452
rect 1768 6409 1777 6443
rect 1777 6409 1811 6443
rect 1811 6409 1820 6443
rect 1768 6400 1820 6409
rect 2412 6400 2464 6452
rect 2872 6400 2924 6452
rect 4160 6400 4212 6452
rect 4620 6400 4672 6452
rect 10324 6443 10376 6452
rect 10324 6409 10333 6443
rect 10333 6409 10367 6443
rect 10367 6409 10376 6443
rect 10324 6400 10376 6409
rect 10416 6400 10468 6452
rect 12256 6443 12308 6452
rect 2504 6332 2556 6384
rect 6644 6332 6696 6384
rect 1216 6264 1268 6316
rect 1768 6264 1820 6316
rect 1952 6307 2004 6316
rect 1952 6273 1961 6307
rect 1961 6273 1995 6307
rect 1995 6273 2004 6307
rect 1952 6264 2004 6273
rect 2688 6264 2740 6316
rect 4436 6264 4488 6316
rect 1492 6196 1544 6248
rect 2320 6196 2372 6248
rect 2596 6196 2648 6248
rect 6000 6264 6052 6316
rect 9312 6264 9364 6316
rect 9680 6307 9732 6316
rect 9680 6273 9689 6307
rect 9689 6273 9723 6307
rect 9723 6273 9732 6307
rect 9680 6264 9732 6273
rect 9772 6264 9824 6316
rect 11520 6264 11572 6316
rect 6920 6239 6972 6248
rect 6920 6205 6929 6239
rect 6929 6205 6963 6239
rect 6963 6205 6972 6239
rect 6920 6196 6972 6205
rect 10416 6196 10468 6248
rect 8944 6128 8996 6180
rect 12256 6409 12265 6443
rect 12265 6409 12299 6443
rect 12299 6409 12308 6443
rect 12256 6400 12308 6409
rect 13084 6400 13136 6452
rect 14188 6400 14240 6452
rect 14924 6443 14976 6452
rect 14924 6409 14933 6443
rect 14933 6409 14967 6443
rect 14967 6409 14976 6443
rect 14924 6400 14976 6409
rect 15016 6400 15068 6452
rect 15384 6400 15436 6452
rect 13452 6264 13504 6316
rect 13820 6307 13872 6316
rect 13820 6273 13829 6307
rect 13829 6273 13863 6307
rect 13863 6273 13872 6307
rect 13820 6264 13872 6273
rect 14004 6264 14056 6316
rect 14372 6264 14424 6316
rect 14740 6307 14792 6316
rect 14740 6273 14749 6307
rect 14749 6273 14783 6307
rect 14783 6273 14792 6307
rect 14740 6264 14792 6273
rect 16120 6332 16172 6384
rect 12624 6239 12676 6248
rect 12624 6205 12633 6239
rect 12633 6205 12667 6239
rect 12667 6205 12676 6239
rect 12624 6196 12676 6205
rect 15476 6196 15528 6248
rect 16304 6264 16356 6316
rect 17960 6400 18012 6452
rect 18144 6400 18196 6452
rect 19892 6400 19944 6452
rect 22192 6400 22244 6452
rect 16488 6332 16540 6384
rect 16764 6264 16816 6316
rect 17224 6332 17276 6384
rect 17316 6307 17368 6316
rect 16028 6196 16080 6248
rect 17316 6273 17325 6307
rect 17325 6273 17359 6307
rect 17359 6273 17368 6307
rect 17316 6264 17368 6273
rect 17684 6264 17736 6316
rect 21732 6264 21784 6316
rect 17868 6239 17920 6248
rect 17868 6205 17877 6239
rect 17877 6205 17911 6239
rect 17911 6205 17920 6239
rect 17868 6196 17920 6205
rect 17960 6196 18012 6248
rect 27068 6400 27120 6452
rect 27436 6400 27488 6452
rect 29276 6400 29328 6452
rect 30380 6400 30432 6452
rect 26700 6332 26752 6384
rect 22468 6307 22520 6316
rect 22468 6273 22477 6307
rect 22477 6273 22511 6307
rect 22511 6273 22520 6307
rect 22468 6264 22520 6273
rect 24492 6264 24544 6316
rect 24860 6307 24912 6316
rect 24860 6273 24869 6307
rect 24869 6273 24903 6307
rect 24903 6273 24912 6307
rect 24860 6264 24912 6273
rect 24952 6264 25004 6316
rect 25596 6307 25648 6316
rect 25596 6273 25605 6307
rect 25605 6273 25639 6307
rect 25639 6273 25648 6307
rect 25596 6264 25648 6273
rect 25780 6307 25832 6316
rect 25780 6273 25789 6307
rect 25789 6273 25823 6307
rect 25823 6273 25832 6307
rect 25780 6264 25832 6273
rect 22836 6196 22888 6248
rect 25688 6196 25740 6248
rect 20904 6171 20956 6180
rect 20904 6137 20913 6171
rect 20913 6137 20947 6171
rect 20947 6137 20956 6171
rect 20904 6128 20956 6137
rect 24584 6128 24636 6180
rect 25964 6307 26016 6316
rect 25964 6273 25973 6307
rect 25973 6273 26007 6307
rect 26007 6273 26016 6307
rect 25964 6264 26016 6273
rect 26516 6264 26568 6316
rect 27344 6264 27396 6316
rect 27988 6264 28040 6316
rect 29184 6307 29236 6316
rect 29184 6273 29193 6307
rect 29193 6273 29227 6307
rect 29227 6273 29236 6307
rect 29184 6264 29236 6273
rect 30472 6264 30524 6316
rect 30748 6264 30800 6316
rect 31300 6264 31352 6316
rect 27620 6196 27672 6248
rect 29736 6128 29788 6180
rect 1492 6060 1544 6112
rect 4344 6060 4396 6112
rect 4712 6060 4764 6112
rect 10600 6060 10652 6112
rect 13820 6060 13872 6112
rect 15016 6060 15068 6112
rect 15936 6060 15988 6112
rect 16580 6060 16632 6112
rect 16856 6060 16908 6112
rect 17960 6060 18012 6112
rect 20720 6060 20772 6112
rect 22100 6060 22152 6112
rect 22652 6103 22704 6112
rect 22652 6069 22661 6103
rect 22661 6069 22695 6103
rect 22695 6069 22704 6103
rect 22652 6060 22704 6069
rect 23480 6103 23532 6112
rect 23480 6069 23489 6103
rect 23489 6069 23523 6103
rect 23523 6069 23532 6103
rect 23480 6060 23532 6069
rect 23756 6060 23808 6112
rect 25780 6060 25832 6112
rect 27068 6060 27120 6112
rect 28632 6060 28684 6112
rect 30656 6060 30708 6112
rect 2136 5958 2188 6010
rect 12440 5958 12492 6010
rect 22744 5958 22796 6010
rect 1492 5856 1544 5908
rect 2412 5788 2464 5840
rect 3608 5788 3660 5840
rect 3884 5788 3936 5840
rect 5080 5788 5132 5840
rect 6368 5788 6420 5840
rect 4344 5763 4396 5772
rect 4344 5729 4353 5763
rect 4353 5729 4387 5763
rect 4387 5729 4396 5763
rect 4344 5720 4396 5729
rect 6092 5720 6144 5772
rect 11704 5788 11756 5840
rect 12624 5788 12676 5840
rect 12900 5788 12952 5840
rect 7472 5763 7524 5772
rect 7472 5729 7481 5763
rect 7481 5729 7515 5763
rect 7515 5729 7524 5763
rect 7472 5720 7524 5729
rect 9496 5763 9548 5772
rect 9496 5729 9505 5763
rect 9505 5729 9539 5763
rect 9539 5729 9548 5763
rect 9496 5720 9548 5729
rect 9956 5720 10008 5772
rect 2688 5584 2740 5636
rect 4252 5652 4304 5704
rect 5632 5652 5684 5704
rect 8944 5652 8996 5704
rect 9404 5695 9456 5704
rect 9404 5661 9413 5695
rect 9413 5661 9447 5695
rect 9447 5661 9456 5695
rect 9404 5652 9456 5661
rect 11980 5695 12032 5704
rect 5356 5627 5408 5636
rect 5356 5593 5390 5627
rect 5390 5593 5408 5627
rect 5356 5584 5408 5593
rect 5540 5584 5592 5636
rect 7380 5627 7432 5636
rect 7380 5593 7389 5627
rect 7389 5593 7423 5627
rect 7423 5593 7432 5627
rect 7380 5584 7432 5593
rect 8668 5584 8720 5636
rect 11980 5661 11989 5695
rect 11989 5661 12023 5695
rect 12023 5661 12032 5695
rect 11980 5652 12032 5661
rect 13544 5720 13596 5772
rect 15016 5720 15068 5772
rect 12808 5695 12860 5704
rect 12808 5661 12817 5695
rect 12817 5661 12851 5695
rect 12851 5661 12860 5695
rect 12808 5652 12860 5661
rect 13084 5695 13136 5704
rect 13084 5661 13093 5695
rect 13093 5661 13127 5695
rect 13127 5661 13136 5695
rect 13084 5652 13136 5661
rect 10508 5584 10560 5636
rect 13176 5584 13228 5636
rect 14924 5695 14976 5704
rect 14924 5661 14933 5695
rect 14933 5661 14967 5695
rect 14967 5661 14976 5695
rect 15936 5720 15988 5772
rect 16948 5788 17000 5840
rect 19156 5788 19208 5840
rect 20628 5831 20680 5840
rect 20628 5797 20637 5831
rect 20637 5797 20671 5831
rect 20671 5797 20680 5831
rect 20628 5788 20680 5797
rect 17316 5720 17368 5772
rect 17960 5720 18012 5772
rect 24492 5856 24544 5908
rect 25688 5856 25740 5908
rect 27712 5899 27764 5908
rect 27712 5865 27721 5899
rect 27721 5865 27755 5899
rect 27755 5865 27764 5899
rect 27712 5856 27764 5865
rect 28080 5856 28132 5908
rect 31024 5856 31076 5908
rect 26332 5788 26384 5840
rect 14924 5652 14976 5661
rect 15660 5695 15712 5704
rect 15660 5661 15669 5695
rect 15669 5661 15703 5695
rect 15703 5661 15712 5695
rect 15660 5652 15712 5661
rect 15752 5652 15804 5704
rect 17040 5695 17092 5704
rect 16304 5584 16356 5636
rect 17040 5661 17049 5695
rect 17049 5661 17083 5695
rect 17083 5661 17092 5695
rect 17040 5652 17092 5661
rect 21916 5652 21968 5704
rect 22100 5695 22152 5704
rect 22100 5661 22134 5695
rect 22134 5661 22152 5695
rect 22100 5652 22152 5661
rect 24032 5652 24084 5704
rect 25412 5652 25464 5704
rect 26608 5695 26660 5704
rect 26608 5661 26617 5695
rect 26617 5661 26651 5695
rect 26651 5661 26660 5695
rect 26608 5652 26660 5661
rect 27068 5695 27120 5704
rect 29828 5788 29880 5840
rect 27068 5661 27084 5695
rect 27084 5661 27118 5695
rect 27118 5661 27120 5695
rect 27068 5652 27120 5661
rect 27528 5695 27580 5704
rect 27528 5661 27542 5695
rect 27542 5661 27576 5695
rect 27576 5661 27580 5695
rect 27528 5652 27580 5661
rect 17316 5584 17368 5636
rect 17868 5584 17920 5636
rect 19708 5584 19760 5636
rect 22560 5584 22612 5636
rect 23664 5584 23716 5636
rect 25872 5584 25924 5636
rect 26148 5584 26200 5636
rect 28724 5720 28776 5772
rect 29276 5652 29328 5704
rect 30472 5652 30524 5704
rect 30748 5652 30800 5704
rect 31116 5695 31168 5704
rect 31116 5661 31125 5695
rect 31125 5661 31159 5695
rect 31159 5661 31168 5695
rect 31116 5652 31168 5661
rect 3240 5559 3292 5568
rect 3240 5525 3249 5559
rect 3249 5525 3283 5559
rect 3283 5525 3292 5559
rect 3240 5516 3292 5525
rect 3792 5559 3844 5568
rect 3792 5525 3801 5559
rect 3801 5525 3835 5559
rect 3835 5525 3844 5559
rect 3792 5516 3844 5525
rect 4436 5516 4488 5568
rect 6920 5559 6972 5568
rect 6920 5525 6929 5559
rect 6929 5525 6963 5559
rect 6963 5525 6972 5559
rect 6920 5516 6972 5525
rect 8484 5516 8536 5568
rect 12164 5516 12216 5568
rect 15108 5516 15160 5568
rect 15384 5516 15436 5568
rect 15752 5516 15804 5568
rect 16028 5559 16080 5568
rect 16028 5525 16037 5559
rect 16037 5525 16071 5559
rect 16071 5525 16080 5559
rect 16028 5516 16080 5525
rect 17224 5516 17276 5568
rect 17960 5516 18012 5568
rect 20260 5516 20312 5568
rect 23204 5559 23256 5568
rect 23204 5525 23213 5559
rect 23213 5525 23247 5559
rect 23247 5525 23256 5559
rect 23204 5516 23256 5525
rect 28080 5516 28132 5568
rect 29460 5516 29512 5568
rect 30012 5584 30064 5636
rect 30472 5516 30524 5568
rect 7288 5414 7340 5466
rect 17592 5414 17644 5466
rect 27896 5414 27948 5466
rect 2688 5312 2740 5364
rect 5356 5355 5408 5364
rect 2044 5219 2096 5228
rect 2044 5185 2053 5219
rect 2053 5185 2087 5219
rect 2087 5185 2096 5219
rect 2044 5176 2096 5185
rect 2320 5244 2372 5296
rect 4160 5244 4212 5296
rect 4988 5244 5040 5296
rect 5356 5321 5365 5355
rect 5365 5321 5399 5355
rect 5399 5321 5408 5355
rect 5356 5312 5408 5321
rect 6920 5312 6972 5364
rect 5264 5244 5316 5296
rect 5448 5244 5500 5296
rect 3056 5219 3108 5228
rect 3056 5185 3090 5219
rect 3090 5185 3108 5219
rect 2596 5108 2648 5160
rect 1400 5040 1452 5092
rect 3056 5176 3108 5185
rect 6552 5219 6604 5228
rect 6552 5185 6561 5219
rect 6561 5185 6595 5219
rect 6595 5185 6604 5219
rect 6552 5176 6604 5185
rect 7840 5244 7892 5296
rect 8484 5287 8536 5296
rect 8484 5253 8493 5287
rect 8493 5253 8527 5287
rect 8527 5253 8536 5287
rect 8484 5244 8536 5253
rect 9404 5244 9456 5296
rect 16396 5312 16448 5364
rect 6460 5108 6512 5160
rect 7932 5176 7984 5228
rect 8576 5176 8628 5228
rect 10140 5176 10192 5228
rect 10508 5176 10560 5228
rect 14280 5176 14332 5228
rect 14372 5176 14424 5228
rect 3884 5040 3936 5092
rect 7656 5040 7708 5092
rect 9496 5108 9548 5160
rect 9956 5108 10008 5160
rect 12624 5108 12676 5160
rect 9772 5040 9824 5092
rect 12532 5040 12584 5092
rect 1676 4972 1728 5024
rect 4068 4972 4120 5024
rect 4528 4972 4580 5024
rect 6092 4972 6144 5024
rect 7104 4972 7156 5024
rect 11796 5015 11848 5024
rect 11796 4981 11805 5015
rect 11805 4981 11839 5015
rect 11839 4981 11848 5015
rect 11796 4972 11848 4981
rect 12900 5108 12952 5160
rect 13820 5108 13872 5160
rect 14832 5176 14884 5228
rect 16488 5176 16540 5228
rect 14924 5108 14976 5160
rect 15108 5151 15160 5160
rect 15108 5117 15117 5151
rect 15117 5117 15151 5151
rect 15151 5117 15160 5151
rect 15108 5108 15160 5117
rect 14004 5040 14056 5092
rect 15016 5040 15068 5092
rect 15384 5151 15436 5160
rect 15384 5117 15393 5151
rect 15393 5117 15427 5151
rect 15427 5117 15436 5151
rect 15384 5108 15436 5117
rect 15660 5108 15712 5160
rect 16396 5108 16448 5160
rect 18236 5244 18288 5296
rect 18420 5287 18472 5296
rect 18420 5253 18454 5287
rect 18454 5253 18472 5287
rect 18420 5244 18472 5253
rect 19800 5244 19852 5296
rect 21088 5287 21140 5296
rect 21088 5253 21113 5287
rect 21113 5253 21140 5287
rect 21088 5244 21140 5253
rect 16856 5176 16908 5228
rect 17316 5176 17368 5228
rect 19340 5176 19392 5228
rect 19892 5176 19944 5228
rect 22376 5244 22428 5296
rect 23480 5244 23532 5296
rect 25688 5244 25740 5296
rect 18144 5151 18196 5160
rect 18144 5117 18153 5151
rect 18153 5117 18187 5151
rect 18187 5117 18196 5151
rect 18144 5108 18196 5117
rect 20444 5151 20496 5160
rect 20444 5117 20453 5151
rect 20453 5117 20487 5151
rect 20487 5117 20496 5151
rect 20444 5108 20496 5117
rect 15752 5040 15804 5092
rect 15568 4972 15620 5024
rect 16948 4972 17000 5024
rect 18788 4972 18840 5024
rect 19984 5015 20036 5024
rect 19984 4981 19993 5015
rect 19993 4981 20027 5015
rect 20027 4981 20036 5015
rect 19984 4972 20036 4981
rect 20260 4972 20312 5024
rect 21272 5108 21324 5160
rect 24032 5176 24084 5228
rect 25780 5219 25832 5228
rect 25780 5185 25789 5219
rect 25789 5185 25823 5219
rect 25823 5185 25832 5219
rect 25780 5176 25832 5185
rect 22008 5151 22060 5160
rect 22008 5117 22017 5151
rect 22017 5117 22051 5151
rect 22051 5117 22060 5151
rect 22008 5108 22060 5117
rect 26700 5176 26752 5228
rect 30380 5244 30432 5296
rect 30196 5219 30248 5228
rect 23296 5040 23348 5092
rect 22008 4972 22060 5024
rect 22192 4972 22244 5024
rect 24952 4972 25004 5024
rect 26424 5083 26476 5092
rect 26424 5049 26433 5083
rect 26433 5049 26467 5083
rect 26467 5049 26476 5083
rect 26424 5040 26476 5049
rect 27620 5108 27672 5160
rect 27252 5040 27304 5092
rect 25412 4972 25464 5024
rect 28632 4972 28684 5024
rect 29092 5015 29144 5024
rect 29092 4981 29101 5015
rect 29101 4981 29135 5015
rect 29135 4981 29144 5015
rect 29092 4972 29144 4981
rect 30196 5185 30230 5219
rect 30230 5185 30248 5219
rect 30196 5176 30248 5185
rect 29552 5108 29604 5160
rect 29920 5151 29972 5160
rect 29920 5117 29929 5151
rect 29929 5117 29963 5151
rect 29963 5117 29972 5151
rect 29920 5108 29972 5117
rect 30656 4972 30708 5024
rect 31300 5015 31352 5024
rect 31300 4981 31309 5015
rect 31309 4981 31343 5015
rect 31343 4981 31352 5015
rect 31300 4972 31352 4981
rect 2136 4870 2188 4922
rect 12440 4870 12492 4922
rect 22744 4870 22796 4922
rect 1584 4768 1636 4820
rect 1400 4675 1452 4684
rect 1400 4641 1409 4675
rect 1409 4641 1443 4675
rect 1443 4641 1452 4675
rect 1400 4632 1452 4641
rect 1676 4607 1728 4616
rect 1676 4573 1710 4607
rect 1710 4573 1728 4607
rect 1676 4564 1728 4573
rect 5264 4768 5316 4820
rect 7564 4768 7616 4820
rect 7932 4811 7984 4820
rect 7932 4777 7941 4811
rect 7941 4777 7975 4811
rect 7975 4777 7984 4811
rect 7932 4768 7984 4777
rect 9680 4768 9732 4820
rect 14740 4768 14792 4820
rect 15016 4768 15068 4820
rect 18052 4768 18104 4820
rect 21272 4768 21324 4820
rect 6184 4700 6236 4752
rect 6644 4700 6696 4752
rect 7656 4700 7708 4752
rect 8024 4700 8076 4752
rect 12624 4700 12676 4752
rect 2596 4632 2648 4684
rect 2688 4564 2740 4616
rect 9312 4632 9364 4684
rect 11336 4632 11388 4684
rect 14372 4675 14424 4684
rect 14372 4641 14381 4675
rect 14381 4641 14415 4675
rect 14415 4641 14424 4675
rect 14372 4632 14424 4641
rect 6644 4607 6696 4616
rect 3792 4496 3844 4548
rect 4712 4539 4764 4548
rect 3240 4428 3292 4480
rect 4712 4505 4721 4539
rect 4721 4505 4755 4539
rect 4755 4505 4764 4539
rect 4712 4496 4764 4505
rect 6644 4573 6653 4607
rect 6653 4573 6687 4607
rect 6687 4573 6696 4607
rect 6644 4564 6696 4573
rect 9588 4564 9640 4616
rect 12164 4564 12216 4616
rect 13544 4607 13596 4616
rect 6736 4496 6788 4548
rect 7472 4539 7524 4548
rect 7472 4505 7481 4539
rect 7481 4505 7515 4539
rect 7515 4505 7524 4539
rect 7472 4496 7524 4505
rect 10324 4496 10376 4548
rect 13544 4573 13553 4607
rect 13553 4573 13587 4607
rect 13587 4573 13596 4607
rect 13544 4564 13596 4573
rect 14096 4607 14148 4616
rect 14096 4573 14105 4607
rect 14105 4573 14139 4607
rect 14139 4573 14148 4607
rect 15108 4632 15160 4684
rect 14096 4564 14148 4573
rect 15016 4564 15068 4616
rect 15844 4700 15896 4752
rect 16028 4700 16080 4752
rect 16304 4700 16356 4752
rect 17316 4700 17368 4752
rect 22100 4700 22152 4752
rect 23112 4700 23164 4752
rect 16396 4632 16448 4684
rect 18328 4632 18380 4684
rect 18604 4675 18656 4684
rect 18604 4641 18613 4675
rect 18613 4641 18647 4675
rect 18647 4641 18656 4675
rect 20260 4675 20312 4684
rect 18604 4632 18656 4641
rect 20260 4641 20269 4675
rect 20269 4641 20303 4675
rect 20303 4641 20312 4675
rect 20260 4632 20312 4641
rect 20628 4632 20680 4684
rect 23204 4632 23256 4684
rect 23572 4632 23624 4684
rect 23848 4632 23900 4684
rect 26240 4700 26292 4752
rect 24860 4675 24912 4684
rect 24860 4641 24869 4675
rect 24869 4641 24903 4675
rect 24903 4641 24912 4675
rect 24860 4632 24912 4641
rect 16856 4564 16908 4616
rect 15200 4496 15252 4548
rect 15568 4539 15620 4548
rect 15568 4505 15577 4539
rect 15577 4505 15611 4539
rect 15611 4505 15620 4539
rect 15568 4496 15620 4505
rect 15936 4496 15988 4548
rect 17316 4564 17368 4616
rect 20076 4607 20128 4616
rect 17132 4496 17184 4548
rect 17684 4496 17736 4548
rect 18328 4496 18380 4548
rect 20076 4573 20085 4607
rect 20085 4573 20119 4607
rect 20119 4573 20128 4607
rect 20076 4564 20128 4573
rect 20996 4607 21048 4616
rect 20996 4573 21005 4607
rect 21005 4573 21039 4607
rect 21039 4573 21048 4607
rect 20996 4564 21048 4573
rect 21180 4607 21232 4616
rect 21180 4573 21189 4607
rect 21189 4573 21223 4607
rect 21223 4573 21232 4607
rect 21180 4564 21232 4573
rect 21732 4607 21784 4616
rect 21732 4573 21741 4607
rect 21741 4573 21775 4607
rect 21775 4573 21784 4607
rect 21732 4564 21784 4573
rect 19156 4496 19208 4548
rect 20628 4496 20680 4548
rect 22560 4564 22612 4616
rect 27988 4632 28040 4684
rect 29184 4632 29236 4684
rect 29552 4675 29604 4684
rect 29552 4641 29561 4675
rect 29561 4641 29595 4675
rect 29595 4641 29604 4675
rect 29552 4632 29604 4641
rect 28080 4564 28132 4616
rect 28540 4564 28592 4616
rect 26976 4496 27028 4548
rect 27804 4496 27856 4548
rect 29368 4496 29420 4548
rect 5080 4471 5132 4480
rect 5080 4437 5089 4471
rect 5089 4437 5123 4471
rect 5123 4437 5132 4471
rect 5080 4428 5132 4437
rect 5264 4471 5316 4480
rect 5264 4437 5273 4471
rect 5273 4437 5307 4471
rect 5307 4437 5316 4471
rect 5264 4428 5316 4437
rect 6368 4428 6420 4480
rect 9496 4428 9548 4480
rect 13544 4428 13596 4480
rect 15752 4428 15804 4480
rect 20168 4428 20220 4480
rect 28264 4428 28316 4480
rect 28356 4428 28408 4480
rect 30012 4428 30064 4480
rect 31116 4428 31168 4480
rect 7288 4326 7340 4378
rect 17592 4326 17644 4378
rect 27896 4326 27948 4378
rect 2044 4224 2096 4276
rect 4712 4224 4764 4276
rect 4988 4224 5040 4276
rect 7472 4224 7524 4276
rect 9956 4224 10008 4276
rect 10324 4267 10376 4276
rect 10324 4233 10333 4267
rect 10333 4233 10367 4267
rect 10367 4233 10376 4267
rect 10324 4224 10376 4233
rect 2228 4088 2280 4140
rect 2412 4131 2464 4140
rect 2412 4097 2421 4131
rect 2421 4097 2455 4131
rect 2455 4097 2464 4131
rect 2412 4088 2464 4097
rect 2688 4088 2740 4140
rect 2872 4088 2924 4140
rect 3976 4156 4028 4208
rect 5264 4156 5316 4208
rect 14004 4224 14056 4276
rect 14280 4224 14332 4276
rect 15200 4224 15252 4276
rect 15936 4224 15988 4276
rect 16488 4224 16540 4276
rect 11888 4199 11940 4208
rect 11888 4165 11897 4199
rect 11897 4165 11931 4199
rect 11931 4165 11940 4199
rect 11888 4156 11940 4165
rect 13084 4156 13136 4208
rect 3792 4088 3844 4140
rect 4252 4131 4304 4140
rect 4252 4097 4261 4131
rect 4261 4097 4295 4131
rect 4295 4097 4304 4131
rect 4252 4088 4304 4097
rect 5448 4088 5500 4140
rect 7380 4088 7432 4140
rect 7656 4088 7708 4140
rect 8576 4131 8628 4140
rect 8576 4097 8585 4131
rect 8585 4097 8619 4131
rect 8619 4097 8628 4131
rect 8576 4088 8628 4097
rect 9312 4088 9364 4140
rect 3700 4063 3752 4072
rect 3700 4029 3709 4063
rect 3709 4029 3743 4063
rect 3743 4029 3752 4063
rect 3700 4020 3752 4029
rect 7104 4020 7156 4072
rect 2412 3952 2464 4004
rect 3516 3952 3568 4004
rect 5816 3952 5868 4004
rect 6736 3952 6788 4004
rect 9496 4020 9548 4072
rect 9956 4088 10008 4140
rect 11704 4088 11756 4140
rect 14280 4131 14332 4140
rect 14280 4097 14289 4131
rect 14289 4097 14323 4131
rect 14323 4097 14332 4131
rect 14280 4088 14332 4097
rect 14372 4088 14424 4140
rect 15016 4156 15068 4208
rect 17224 4199 17276 4208
rect 17224 4165 17233 4199
rect 17233 4165 17267 4199
rect 17267 4165 17276 4199
rect 17224 4156 17276 4165
rect 15844 4131 15896 4140
rect 15844 4097 15853 4131
rect 15853 4097 15887 4131
rect 15887 4097 15896 4131
rect 15844 4088 15896 4097
rect 16948 4131 17000 4140
rect 17684 4224 17736 4276
rect 18328 4224 18380 4276
rect 18972 4156 19024 4208
rect 20444 4224 20496 4276
rect 29368 4267 29420 4276
rect 29368 4233 29377 4267
rect 29377 4233 29411 4267
rect 29411 4233 29420 4267
rect 29368 4224 29420 4233
rect 16948 4097 16964 4131
rect 16964 4097 16998 4131
rect 16998 4097 17000 4131
rect 16948 4088 17000 4097
rect 7932 3995 7984 4004
rect 7932 3961 7941 3995
rect 7941 3961 7975 3995
rect 7975 3961 7984 3995
rect 7932 3952 7984 3961
rect 3148 3884 3200 3936
rect 5724 3884 5776 3936
rect 6644 3884 6696 3936
rect 6920 3884 6972 3936
rect 12808 3952 12860 4004
rect 16948 3952 17000 4004
rect 17868 4088 17920 4140
rect 18604 4131 18656 4140
rect 18604 4097 18613 4131
rect 18613 4097 18647 4131
rect 18647 4097 18656 4131
rect 18604 4088 18656 4097
rect 18788 4131 18840 4140
rect 18788 4097 18797 4131
rect 18797 4097 18831 4131
rect 18831 4097 18840 4131
rect 18788 4088 18840 4097
rect 19340 4088 19392 4140
rect 22100 4156 22152 4208
rect 24860 4156 24912 4208
rect 25228 4156 25280 4208
rect 20168 4131 20220 4140
rect 20168 4097 20202 4131
rect 20202 4097 20220 4131
rect 22008 4131 22060 4140
rect 20168 4088 20220 4097
rect 22008 4097 22017 4131
rect 22017 4097 22051 4131
rect 22051 4097 22060 4131
rect 22008 4088 22060 4097
rect 22560 4131 22612 4140
rect 22560 4097 22569 4131
rect 22569 4097 22603 4131
rect 22603 4097 22612 4131
rect 22560 4088 22612 4097
rect 23848 4131 23900 4140
rect 23848 4097 23857 4131
rect 23857 4097 23891 4131
rect 23891 4097 23900 4131
rect 23848 4088 23900 4097
rect 27344 4199 27396 4208
rect 27344 4165 27353 4199
rect 27353 4165 27387 4199
rect 27387 4165 27396 4199
rect 27344 4156 27396 4165
rect 19156 4020 19208 4072
rect 19248 4020 19300 4072
rect 10600 3884 10652 3936
rect 12900 3884 12952 3936
rect 13268 3884 13320 3936
rect 16764 3884 16816 3936
rect 17684 3884 17736 3936
rect 19248 3927 19300 3936
rect 19248 3893 19257 3927
rect 19257 3893 19291 3927
rect 19291 3893 19300 3927
rect 19248 3884 19300 3893
rect 21180 4020 21232 4072
rect 22652 4020 22704 4072
rect 23204 4020 23256 4072
rect 24124 4063 24176 4072
rect 24124 4029 24133 4063
rect 24133 4029 24167 4063
rect 24167 4029 24176 4063
rect 24124 4020 24176 4029
rect 25044 4020 25096 4072
rect 25688 4088 25740 4140
rect 26424 4131 26476 4140
rect 26424 4097 26433 4131
rect 26433 4097 26467 4131
rect 26467 4097 26476 4131
rect 26424 4088 26476 4097
rect 26608 4088 26660 4140
rect 27068 4131 27120 4140
rect 27068 4097 27078 4131
rect 27078 4097 27112 4131
rect 27112 4097 27120 4131
rect 27252 4131 27304 4140
rect 27068 4088 27120 4097
rect 27252 4097 27261 4131
rect 27261 4097 27295 4131
rect 27295 4097 27304 4131
rect 27252 4088 27304 4097
rect 28264 4131 28316 4140
rect 26332 4020 26384 4072
rect 26700 4020 26752 4072
rect 28264 4097 28273 4131
rect 28273 4097 28307 4131
rect 28307 4097 28316 4131
rect 28264 4088 28316 4097
rect 28540 4131 28592 4140
rect 28540 4097 28549 4131
rect 28549 4097 28583 4131
rect 28583 4097 28592 4131
rect 28540 4088 28592 4097
rect 29460 4088 29512 4140
rect 29828 4131 29880 4140
rect 29828 4097 29837 4131
rect 29837 4097 29871 4131
rect 29871 4097 29880 4131
rect 30472 4131 30524 4140
rect 29828 4088 29880 4097
rect 30472 4097 30481 4131
rect 30481 4097 30515 4131
rect 30515 4097 30524 4131
rect 30472 4088 30524 4097
rect 30748 4131 30800 4140
rect 30748 4097 30757 4131
rect 30757 4097 30791 4131
rect 30791 4097 30800 4131
rect 30748 4088 30800 4097
rect 31300 4156 31352 4208
rect 29092 4020 29144 4072
rect 30104 4020 30156 4072
rect 30564 4020 30616 4072
rect 29736 3995 29788 4004
rect 29736 3961 29745 3995
rect 29745 3961 29779 3995
rect 29779 3961 29788 3995
rect 29736 3952 29788 3961
rect 21824 3927 21876 3936
rect 21824 3893 21833 3927
rect 21833 3893 21867 3927
rect 21867 3893 21876 3927
rect 21824 3884 21876 3893
rect 23572 3884 23624 3936
rect 26056 3884 26108 3936
rect 28632 3884 28684 3936
rect 2136 3782 2188 3834
rect 12440 3782 12492 3834
rect 22744 3782 22796 3834
rect 5080 3680 5132 3732
rect 5448 3723 5500 3732
rect 5448 3689 5457 3723
rect 5457 3689 5491 3723
rect 5491 3689 5500 3723
rect 5448 3680 5500 3689
rect 5724 3680 5776 3732
rect 6092 3680 6144 3732
rect 12716 3680 12768 3732
rect 13820 3680 13872 3732
rect 17040 3680 17092 3732
rect 3148 3655 3200 3664
rect 3148 3621 3157 3655
rect 3157 3621 3191 3655
rect 3191 3621 3200 3655
rect 3148 3612 3200 3621
rect 2688 3544 2740 3596
rect 2412 3476 2464 3528
rect 3700 3544 3752 3596
rect 4528 3544 4580 3596
rect 6276 3544 6328 3596
rect 4344 3476 4396 3528
rect 5172 3476 5224 3528
rect 4712 3340 4764 3392
rect 6092 3408 6144 3460
rect 9220 3612 9272 3664
rect 6828 3544 6880 3596
rect 6920 3519 6972 3528
rect 6460 3408 6512 3460
rect 6644 3451 6696 3460
rect 6644 3417 6653 3451
rect 6653 3417 6687 3451
rect 6687 3417 6696 3451
rect 6644 3408 6696 3417
rect 6920 3485 6929 3519
rect 6929 3485 6963 3519
rect 6963 3485 6972 3519
rect 6920 3476 6972 3485
rect 9220 3519 9272 3528
rect 9220 3485 9229 3519
rect 9229 3485 9263 3519
rect 9263 3485 9272 3519
rect 9220 3476 9272 3485
rect 9496 3519 9548 3528
rect 9496 3485 9505 3519
rect 9505 3485 9539 3519
rect 9539 3485 9548 3519
rect 9496 3476 9548 3485
rect 9772 3476 9824 3528
rect 10692 3612 10744 3664
rect 10416 3476 10468 3528
rect 10692 3476 10744 3528
rect 7564 3408 7616 3460
rect 7840 3408 7892 3460
rect 10968 3408 11020 3460
rect 16856 3612 16908 3664
rect 11336 3544 11388 3596
rect 13176 3544 13228 3596
rect 11796 3519 11848 3528
rect 11796 3485 11830 3519
rect 11830 3485 11848 3519
rect 11796 3476 11848 3485
rect 15292 3544 15344 3596
rect 15476 3544 15528 3596
rect 15568 3544 15620 3596
rect 16488 3544 16540 3596
rect 13544 3519 13596 3528
rect 13544 3485 13553 3519
rect 13553 3485 13587 3519
rect 13587 3485 13596 3519
rect 13544 3476 13596 3485
rect 14280 3519 14332 3528
rect 14280 3485 14289 3519
rect 14289 3485 14323 3519
rect 14323 3485 14332 3519
rect 14280 3476 14332 3485
rect 14372 3476 14424 3528
rect 14832 3476 14884 3528
rect 16028 3476 16080 3528
rect 16580 3476 16632 3528
rect 16764 3519 16816 3528
rect 16764 3485 16774 3519
rect 16774 3485 16808 3519
rect 16808 3485 16816 3519
rect 16764 3476 16816 3485
rect 17868 3476 17920 3528
rect 19892 3723 19944 3732
rect 19892 3689 19901 3723
rect 19901 3689 19935 3723
rect 19935 3689 19944 3723
rect 19892 3680 19944 3689
rect 20996 3723 21048 3732
rect 20996 3689 21005 3723
rect 21005 3689 21039 3723
rect 21039 3689 21048 3723
rect 20996 3680 21048 3689
rect 23664 3680 23716 3732
rect 23756 3723 23808 3732
rect 23756 3689 23765 3723
rect 23765 3689 23799 3723
rect 23799 3689 23808 3723
rect 23756 3680 23808 3689
rect 26240 3680 26292 3732
rect 26608 3680 26660 3732
rect 30656 3723 30708 3732
rect 30656 3689 30665 3723
rect 30665 3689 30699 3723
rect 30699 3689 30708 3723
rect 30656 3680 30708 3689
rect 20904 3612 20956 3664
rect 18328 3544 18380 3596
rect 19248 3544 19300 3596
rect 21548 3612 21600 3664
rect 26424 3612 26476 3664
rect 29736 3612 29788 3664
rect 31024 3655 31076 3664
rect 31024 3621 31033 3655
rect 31033 3621 31067 3655
rect 31067 3621 31076 3655
rect 31024 3612 31076 3621
rect 16488 3408 16540 3460
rect 17040 3451 17092 3460
rect 17040 3417 17049 3451
rect 17049 3417 17083 3451
rect 17083 3417 17092 3451
rect 17040 3408 17092 3417
rect 17224 3408 17276 3460
rect 18696 3519 18748 3528
rect 18696 3485 18705 3519
rect 18705 3485 18739 3519
rect 18739 3485 18748 3519
rect 18696 3476 18748 3485
rect 19340 3476 19392 3528
rect 20260 3476 20312 3528
rect 18604 3408 18656 3460
rect 20628 3476 20680 3528
rect 24124 3544 24176 3596
rect 20904 3408 20956 3460
rect 22192 3476 22244 3528
rect 22284 3519 22336 3528
rect 22284 3485 22293 3519
rect 22293 3485 22327 3519
rect 22327 3485 22336 3519
rect 22560 3519 22612 3528
rect 22284 3476 22336 3485
rect 22560 3485 22569 3519
rect 22569 3485 22603 3519
rect 22603 3485 22612 3519
rect 22560 3476 22612 3485
rect 22836 3476 22888 3528
rect 23572 3519 23624 3528
rect 23572 3485 23581 3519
rect 23581 3485 23615 3519
rect 23615 3485 23624 3519
rect 23572 3476 23624 3485
rect 25044 3476 25096 3528
rect 25228 3519 25280 3528
rect 25228 3485 25237 3519
rect 25237 3485 25271 3519
rect 25271 3485 25280 3519
rect 25228 3476 25280 3485
rect 25596 3476 25648 3528
rect 28356 3544 28408 3596
rect 28632 3544 28684 3596
rect 31116 3587 31168 3596
rect 26148 3519 26200 3528
rect 26148 3485 26157 3519
rect 26157 3485 26191 3519
rect 26191 3485 26200 3519
rect 26148 3476 26200 3485
rect 26516 3476 26568 3528
rect 26976 3519 27028 3528
rect 26976 3485 26985 3519
rect 26985 3485 27019 3519
rect 27019 3485 27028 3519
rect 26976 3476 27028 3485
rect 27712 3476 27764 3528
rect 29736 3519 29788 3528
rect 28724 3451 28776 3460
rect 7104 3340 7156 3392
rect 7748 3383 7800 3392
rect 7748 3349 7757 3383
rect 7757 3349 7791 3383
rect 7791 3349 7800 3383
rect 7748 3340 7800 3349
rect 10048 3340 10100 3392
rect 11612 3340 11664 3392
rect 13544 3340 13596 3392
rect 18420 3340 18472 3392
rect 19800 3340 19852 3392
rect 24860 3340 24912 3392
rect 25872 3340 25924 3392
rect 28724 3417 28733 3451
rect 28733 3417 28767 3451
rect 28767 3417 28776 3451
rect 28724 3408 28776 3417
rect 29736 3485 29745 3519
rect 29745 3485 29779 3519
rect 29779 3485 29788 3519
rect 29736 3476 29788 3485
rect 30012 3519 30064 3528
rect 30012 3485 30021 3519
rect 30021 3485 30055 3519
rect 30055 3485 30064 3519
rect 30012 3476 30064 3485
rect 31116 3553 31125 3587
rect 31125 3553 31159 3587
rect 31159 3553 31168 3587
rect 31116 3544 31168 3553
rect 30748 3408 30800 3460
rect 30564 3340 30616 3392
rect 7288 3238 7340 3290
rect 17592 3238 17644 3290
rect 27896 3238 27948 3290
rect 2780 3136 2832 3188
rect 9680 3136 9732 3188
rect 2228 3068 2280 3120
rect 2320 3000 2372 3052
rect 2596 3043 2648 3052
rect 2596 3009 2605 3043
rect 2605 3009 2639 3043
rect 2639 3009 2648 3043
rect 2596 3000 2648 3009
rect 4344 3068 4396 3120
rect 4160 3000 4212 3052
rect 3976 2932 4028 2984
rect 6092 3068 6144 3120
rect 7748 3068 7800 3120
rect 11704 3136 11756 3188
rect 13820 3136 13872 3188
rect 14832 3136 14884 3188
rect 15568 3136 15620 3188
rect 17684 3136 17736 3188
rect 20076 3136 20128 3188
rect 6276 3000 6328 3052
rect 6552 3043 6604 3052
rect 6552 3009 6561 3043
rect 6561 3009 6595 3043
rect 6595 3009 6604 3043
rect 6552 3000 6604 3009
rect 6736 3000 6788 3052
rect 6920 3000 6972 3052
rect 8668 3000 8720 3052
rect 8944 3043 8996 3052
rect 8944 3009 8953 3043
rect 8953 3009 8987 3043
rect 8987 3009 8996 3043
rect 10600 3068 10652 3120
rect 11336 3068 11388 3120
rect 9588 3043 9640 3052
rect 8944 3000 8996 3009
rect 9588 3009 9597 3043
rect 9597 3009 9631 3043
rect 9631 3009 9640 3043
rect 9588 3000 9640 3009
rect 3516 2864 3568 2916
rect 4436 2864 4488 2916
rect 2320 2796 2372 2848
rect 3332 2796 3384 2848
rect 3792 2796 3844 2848
rect 4804 2796 4856 2848
rect 8208 2975 8260 2984
rect 8208 2941 8217 2975
rect 8217 2941 8251 2975
rect 8251 2941 8260 2975
rect 8208 2932 8260 2941
rect 11612 3000 11664 3052
rect 12716 3068 12768 3120
rect 12900 3000 12952 3052
rect 13360 3000 13412 3052
rect 6184 2864 6236 2916
rect 6460 2864 6512 2916
rect 7564 2907 7616 2916
rect 7564 2873 7573 2907
rect 7573 2873 7607 2907
rect 7607 2873 7616 2907
rect 7564 2864 7616 2873
rect 10968 2907 11020 2916
rect 10968 2873 10977 2907
rect 10977 2873 11011 2907
rect 11011 2873 11020 2907
rect 10968 2864 11020 2873
rect 11060 2864 11112 2916
rect 14372 3068 14424 3120
rect 14280 3000 14332 3052
rect 15660 3068 15712 3120
rect 16120 3068 16172 3120
rect 16488 3068 16540 3120
rect 30748 3179 30800 3188
rect 30748 3145 30757 3179
rect 30757 3145 30791 3179
rect 30791 3145 30800 3179
rect 30748 3136 30800 3145
rect 31116 3136 31168 3188
rect 25228 3068 25280 3120
rect 15752 3043 15804 3052
rect 15752 3009 15761 3043
rect 15761 3009 15795 3043
rect 15795 3009 15804 3043
rect 15752 3000 15804 3009
rect 16856 3043 16908 3052
rect 14188 2932 14240 2984
rect 16856 3009 16865 3043
rect 16865 3009 16899 3043
rect 16899 3009 16908 3043
rect 16856 3000 16908 3009
rect 17132 3043 17184 3052
rect 17132 3009 17141 3043
rect 17141 3009 17175 3043
rect 17175 3009 17184 3043
rect 17132 3000 17184 3009
rect 17316 3043 17368 3052
rect 17316 3009 17325 3043
rect 17325 3009 17359 3043
rect 17359 3009 17368 3043
rect 17316 3000 17368 3009
rect 18604 3043 18656 3052
rect 18604 3009 18613 3043
rect 18613 3009 18647 3043
rect 18647 3009 18656 3043
rect 18604 3000 18656 3009
rect 19800 3000 19852 3052
rect 20260 3000 20312 3052
rect 20904 3043 20956 3052
rect 20904 3009 20913 3043
rect 20913 3009 20947 3043
rect 20947 3009 20956 3043
rect 20904 3000 20956 3009
rect 22284 3043 22336 3052
rect 22284 3009 22293 3043
rect 22293 3009 22327 3043
rect 22327 3009 22336 3043
rect 22284 3000 22336 3009
rect 22560 3043 22612 3052
rect 22560 3009 22569 3043
rect 22569 3009 22603 3043
rect 22603 3009 22612 3043
rect 22560 3000 22612 3009
rect 23020 3000 23072 3052
rect 23112 3000 23164 3052
rect 23296 3000 23348 3052
rect 24492 3000 24544 3052
rect 25044 3000 25096 3052
rect 25872 3000 25924 3052
rect 28264 3068 28316 3120
rect 16948 2932 17000 2984
rect 18972 2932 19024 2984
rect 27988 3000 28040 3052
rect 31208 3068 31260 3120
rect 30656 3000 30708 3052
rect 7104 2796 7156 2848
rect 8116 2796 8168 2848
rect 14924 2796 14976 2848
rect 15844 2796 15896 2848
rect 16856 2864 16908 2916
rect 17868 2864 17920 2916
rect 21272 2864 21324 2916
rect 28540 2932 28592 2984
rect 28724 2932 28776 2984
rect 23020 2864 23072 2916
rect 24584 2907 24636 2916
rect 24584 2873 24593 2907
rect 24593 2873 24627 2907
rect 24627 2873 24636 2907
rect 24584 2864 24636 2873
rect 28908 2864 28960 2916
rect 17776 2796 17828 2848
rect 18236 2796 18288 2848
rect 19800 2796 19852 2848
rect 20444 2796 20496 2848
rect 22652 2796 22704 2848
rect 25320 2839 25372 2848
rect 25320 2805 25329 2839
rect 25329 2805 25363 2839
rect 25363 2805 25372 2839
rect 25320 2796 25372 2805
rect 26148 2796 26200 2848
rect 2136 2694 2188 2746
rect 12440 2694 12492 2746
rect 22744 2694 22796 2746
rect 2596 2592 2648 2644
rect 1400 2456 1452 2508
rect 4160 2592 4212 2644
rect 4528 2592 4580 2644
rect 8944 2592 8996 2644
rect 9864 2592 9916 2644
rect 10692 2592 10744 2644
rect 13084 2592 13136 2644
rect 14280 2592 14332 2644
rect 16212 2592 16264 2644
rect 10876 2524 10928 2576
rect 18696 2592 18748 2644
rect 22836 2592 22888 2644
rect 25228 2592 25280 2644
rect 27344 2592 27396 2644
rect 29092 2592 29144 2644
rect 30656 2635 30708 2644
rect 19248 2524 19300 2576
rect 6552 2388 6604 2440
rect 6736 2388 6788 2440
rect 8116 2456 8168 2508
rect 11336 2456 11388 2508
rect 12808 2456 12860 2508
rect 14556 2499 14608 2508
rect 14556 2465 14565 2499
rect 14565 2465 14599 2499
rect 14599 2465 14608 2499
rect 14556 2456 14608 2465
rect 18788 2456 18840 2508
rect 7564 2431 7616 2440
rect 7564 2397 7573 2431
rect 7573 2397 7607 2431
rect 7607 2397 7616 2431
rect 7564 2388 7616 2397
rect 9588 2388 9640 2440
rect 10508 2388 10560 2440
rect 16212 2388 16264 2440
rect 18144 2388 18196 2440
rect 18420 2431 18472 2440
rect 18420 2397 18429 2431
rect 18429 2397 18463 2431
rect 18463 2397 18472 2431
rect 18420 2388 18472 2397
rect 18604 2431 18656 2440
rect 18604 2397 18613 2431
rect 18613 2397 18647 2431
rect 18647 2397 18656 2431
rect 18604 2388 18656 2397
rect 21916 2388 21968 2440
rect 23112 2388 23164 2440
rect 24492 2524 24544 2576
rect 28356 2524 28408 2576
rect 30656 2601 30665 2635
rect 30665 2601 30699 2635
rect 30699 2601 30708 2635
rect 30656 2592 30708 2601
rect 2044 2320 2096 2372
rect 3148 2320 3200 2372
rect 3516 2252 3568 2304
rect 4436 2252 4488 2304
rect 7380 2252 7432 2304
rect 10232 2320 10284 2372
rect 13084 2320 13136 2372
rect 15660 2320 15712 2372
rect 16672 2363 16724 2372
rect 16672 2329 16706 2363
rect 16706 2329 16724 2363
rect 16672 2320 16724 2329
rect 19800 2320 19852 2372
rect 22928 2320 22980 2372
rect 24032 2388 24084 2440
rect 27620 2388 27672 2440
rect 28264 2388 28316 2440
rect 28540 2388 28592 2440
rect 24584 2320 24636 2372
rect 25780 2320 25832 2372
rect 25964 2320 26016 2372
rect 28816 2431 28868 2440
rect 28816 2397 28825 2431
rect 28825 2397 28859 2431
rect 28859 2397 28868 2431
rect 28816 2388 28868 2397
rect 30104 2456 30156 2508
rect 29736 2431 29788 2440
rect 29736 2397 29738 2431
rect 29738 2397 29772 2431
rect 29772 2397 29788 2431
rect 29736 2388 29788 2397
rect 30012 2431 30064 2440
rect 30012 2397 30021 2431
rect 30021 2397 30055 2431
rect 30055 2397 30064 2431
rect 30012 2388 30064 2397
rect 30288 2431 30340 2440
rect 30288 2397 30297 2431
rect 30297 2397 30331 2431
rect 30331 2397 30340 2431
rect 30288 2388 30340 2397
rect 30564 2388 30616 2440
rect 31024 2431 31076 2440
rect 31024 2397 31033 2431
rect 31033 2397 31067 2431
rect 31067 2397 31076 2431
rect 31024 2388 31076 2397
rect 11060 2252 11112 2304
rect 12072 2252 12124 2304
rect 14096 2252 14148 2304
rect 15936 2295 15988 2304
rect 15936 2261 15945 2295
rect 15945 2261 15979 2295
rect 15979 2261 15988 2295
rect 15936 2252 15988 2261
rect 17040 2252 17092 2304
rect 17316 2252 17368 2304
rect 17776 2295 17828 2304
rect 17776 2261 17785 2295
rect 17785 2261 17819 2295
rect 17819 2261 17828 2295
rect 17776 2252 17828 2261
rect 17868 2252 17920 2304
rect 21456 2252 21508 2304
rect 23572 2252 23624 2304
rect 25136 2252 25188 2304
rect 25872 2295 25924 2304
rect 25872 2261 25881 2295
rect 25881 2261 25915 2295
rect 25915 2261 25924 2295
rect 25872 2252 25924 2261
rect 26240 2252 26292 2304
rect 27068 2252 27120 2304
rect 27988 2252 28040 2304
rect 28080 2252 28132 2304
rect 30840 2252 30892 2304
rect 7288 2150 7340 2202
rect 17592 2150 17644 2202
rect 27896 2150 27948 2202
rect 2044 2048 2096 2100
rect 3148 2091 3200 2100
rect 3148 2057 3157 2091
rect 3157 2057 3191 2091
rect 3191 2057 3200 2091
rect 3148 2048 3200 2057
rect 6828 2048 6880 2100
rect 7564 2048 7616 2100
rect 8208 2048 8260 2100
rect 4712 2023 4764 2032
rect 4712 1989 4746 2023
rect 4746 1989 4764 2023
rect 4712 1980 4764 1989
rect 2320 1955 2372 1964
rect 2320 1921 2329 1955
rect 2329 1921 2363 1955
rect 2363 1921 2372 1955
rect 2320 1912 2372 1921
rect 3332 1955 3384 1964
rect 2688 1844 2740 1896
rect 3332 1921 3341 1955
rect 3341 1921 3375 1955
rect 3375 1921 3384 1955
rect 3332 1912 3384 1921
rect 4068 1912 4120 1964
rect 4160 1912 4212 1964
rect 3056 1844 3108 1896
rect 7012 1980 7064 2032
rect 11060 2048 11112 2100
rect 13360 2023 13412 2032
rect 13360 1989 13369 2023
rect 13369 1989 13403 2023
rect 13403 1989 13412 2023
rect 13360 1980 13412 1989
rect 7196 1955 7248 1964
rect 6552 1751 6604 1760
rect 6552 1717 6561 1751
rect 6561 1717 6595 1751
rect 6595 1717 6604 1751
rect 6552 1708 6604 1717
rect 7196 1921 7205 1955
rect 7205 1921 7239 1955
rect 7239 1921 7248 1955
rect 7196 1912 7248 1921
rect 7472 1955 7524 1964
rect 7472 1921 7506 1955
rect 7506 1921 7524 1955
rect 9588 1955 9640 1964
rect 7472 1912 7524 1921
rect 9588 1921 9597 1955
rect 9597 1921 9631 1955
rect 9631 1921 9640 1955
rect 9588 1912 9640 1921
rect 9680 1912 9732 1964
rect 11336 1912 11388 1964
rect 13544 1955 13596 1964
rect 13544 1921 13553 1955
rect 13553 1921 13587 1955
rect 13587 1921 13596 1955
rect 13544 1912 13596 1921
rect 12900 1819 12952 1828
rect 12900 1785 12909 1819
rect 12909 1785 12943 1819
rect 12943 1785 12952 1819
rect 12900 1776 12952 1785
rect 17868 1980 17920 2032
rect 14556 1955 14608 1964
rect 14556 1921 14565 1955
rect 14565 1921 14599 1955
rect 14599 1921 14608 1955
rect 14556 1912 14608 1921
rect 14832 1955 14884 1964
rect 14832 1921 14866 1955
rect 14866 1921 14884 1955
rect 14832 1912 14884 1921
rect 16856 1912 16908 1964
rect 17132 1912 17184 1964
rect 13544 1708 13596 1760
rect 16580 1844 16632 1896
rect 16764 1844 16816 1896
rect 17776 1912 17828 1964
rect 18144 1980 18196 2032
rect 20628 2048 20680 2100
rect 23020 2048 23072 2100
rect 25596 2048 25648 2100
rect 25964 2091 26016 2100
rect 25964 2057 25973 2091
rect 25973 2057 26007 2091
rect 26007 2057 26016 2091
rect 25964 2048 26016 2057
rect 18328 1955 18380 1964
rect 18328 1921 18362 1955
rect 18362 1921 18380 1955
rect 18328 1912 18380 1921
rect 19984 1912 20036 1964
rect 21916 1955 21968 1964
rect 21916 1921 21925 1955
rect 21925 1921 21959 1955
rect 21959 1921 21968 1955
rect 21916 1912 21968 1921
rect 22468 1912 22520 1964
rect 24032 1955 24084 1964
rect 24032 1921 24041 1955
rect 24041 1921 24075 1955
rect 24075 1921 24084 1955
rect 24032 1912 24084 1921
rect 24676 1912 24728 1964
rect 26148 1955 26200 1964
rect 26148 1921 26157 1955
rect 26157 1921 26191 1955
rect 26191 1921 26200 1955
rect 26148 1912 26200 1921
rect 26332 1955 26384 1964
rect 26332 1921 26341 1955
rect 26341 1921 26375 1955
rect 26375 1921 26384 1955
rect 26332 1912 26384 1921
rect 27344 1912 27396 1964
rect 27620 1980 27672 2032
rect 28908 1980 28960 2032
rect 27712 1955 27764 1964
rect 27712 1921 27746 1955
rect 27746 1921 27764 1955
rect 27712 1912 27764 1921
rect 30656 1912 30708 1964
rect 31300 1955 31352 1964
rect 31300 1921 31309 1955
rect 31309 1921 31343 1955
rect 31343 1921 31352 1955
rect 31300 1912 31352 1921
rect 28816 1819 28868 1828
rect 28816 1785 28825 1819
rect 28825 1785 28859 1819
rect 28859 1785 28868 1819
rect 28816 1776 28868 1785
rect 30288 1776 30340 1828
rect 15752 1708 15804 1760
rect 16856 1751 16908 1760
rect 16856 1717 16865 1751
rect 16865 1717 16899 1751
rect 16899 1717 16908 1751
rect 16856 1708 16908 1717
rect 17684 1708 17736 1760
rect 2136 1606 2188 1658
rect 12440 1606 12492 1658
rect 22744 1606 22796 1658
rect 1860 1504 1912 1556
rect 2872 1504 2924 1556
rect 6276 1504 6328 1556
rect 7472 1504 7524 1556
rect 10232 1547 10284 1556
rect 10232 1513 10241 1547
rect 10241 1513 10275 1547
rect 10275 1513 10284 1547
rect 10232 1504 10284 1513
rect 13084 1547 13136 1556
rect 13084 1513 13093 1547
rect 13093 1513 13127 1547
rect 13127 1513 13136 1547
rect 13084 1504 13136 1513
rect 13544 1504 13596 1556
rect 14832 1504 14884 1556
rect 15660 1547 15712 1556
rect 15660 1513 15669 1547
rect 15669 1513 15703 1547
rect 15703 1513 15712 1547
rect 15660 1504 15712 1513
rect 16672 1547 16724 1556
rect 16672 1513 16681 1547
rect 16681 1513 16715 1547
rect 16715 1513 16724 1547
rect 16672 1504 16724 1513
rect 18328 1504 18380 1556
rect 18604 1547 18656 1556
rect 18604 1513 18613 1547
rect 18613 1513 18647 1547
rect 18647 1513 18656 1547
rect 18604 1504 18656 1513
rect 22468 1547 22520 1556
rect 22468 1513 22477 1547
rect 22477 1513 22511 1547
rect 22511 1513 22520 1547
rect 22468 1504 22520 1513
rect 24676 1547 24728 1556
rect 2964 1436 3016 1488
rect 6552 1436 6604 1488
rect 24676 1513 24685 1547
rect 24685 1513 24719 1547
rect 24719 1513 24728 1547
rect 24676 1504 24728 1513
rect 25780 1547 25832 1556
rect 25780 1513 25789 1547
rect 25789 1513 25823 1547
rect 25823 1513 25832 1547
rect 25780 1504 25832 1513
rect 26332 1504 26384 1556
rect 27712 1504 27764 1556
rect 28816 1547 28868 1556
rect 28816 1513 28825 1547
rect 28825 1513 28859 1547
rect 28859 1513 28868 1547
rect 28816 1504 28868 1513
rect 30656 1547 30708 1556
rect 30656 1513 30665 1547
rect 30665 1513 30699 1547
rect 30699 1513 30708 1547
rect 30656 1504 30708 1513
rect 29644 1436 29696 1488
rect 6828 1411 6880 1420
rect 6828 1377 6837 1411
rect 6837 1377 6871 1411
rect 6871 1377 6880 1411
rect 6828 1368 6880 1377
rect 9956 1368 10008 1420
rect 2504 1343 2556 1352
rect 2504 1309 2513 1343
rect 2513 1309 2547 1343
rect 2547 1309 2556 1343
rect 2504 1300 2556 1309
rect 3884 1343 3936 1352
rect 3884 1309 3893 1343
rect 3893 1309 3927 1343
rect 3927 1309 3936 1343
rect 3884 1300 3936 1309
rect 4896 1300 4948 1352
rect 5816 1343 5868 1352
rect 5816 1309 5825 1343
rect 5825 1309 5859 1343
rect 5859 1309 5868 1343
rect 5816 1300 5868 1309
rect 6368 1300 6420 1352
rect 5724 1232 5776 1284
rect 7380 1300 7432 1352
rect 7840 1300 7892 1352
rect 8392 1343 8444 1352
rect 8392 1309 8401 1343
rect 8401 1309 8435 1343
rect 8435 1309 8444 1343
rect 8392 1300 8444 1309
rect 9220 1343 9272 1352
rect 8300 1232 8352 1284
rect 9220 1309 9229 1343
rect 9229 1309 9263 1343
rect 9263 1309 9272 1343
rect 9220 1300 9272 1309
rect 10048 1300 10100 1352
rect 10600 1343 10652 1352
rect 10600 1309 10609 1343
rect 10609 1309 10643 1343
rect 10643 1309 10652 1343
rect 10600 1300 10652 1309
rect 11704 1343 11756 1352
rect 11704 1309 11713 1343
rect 11713 1309 11747 1343
rect 11747 1309 11756 1343
rect 11704 1300 11756 1309
rect 13268 1343 13320 1352
rect 13268 1309 13277 1343
rect 13277 1309 13311 1343
rect 13311 1309 13320 1343
rect 13268 1300 13320 1309
rect 13820 1368 13872 1420
rect 15936 1368 15988 1420
rect 17684 1368 17736 1420
rect 21548 1368 21600 1420
rect 23204 1368 23256 1420
rect 13636 1300 13688 1352
rect 14924 1343 14976 1352
rect 14924 1309 14933 1343
rect 14933 1309 14967 1343
rect 14967 1309 14976 1343
rect 14924 1300 14976 1309
rect 15844 1343 15896 1352
rect 15844 1309 15853 1343
rect 15853 1309 15887 1343
rect 15887 1309 15896 1343
rect 15844 1300 15896 1309
rect 16028 1343 16080 1352
rect 16028 1309 16037 1343
rect 16037 1309 16071 1343
rect 16071 1309 16080 1343
rect 16028 1300 16080 1309
rect 16580 1300 16632 1352
rect 16856 1343 16908 1352
rect 16856 1309 16865 1343
rect 16865 1309 16899 1343
rect 16899 1309 16908 1343
rect 16856 1300 16908 1309
rect 17960 1300 18012 1352
rect 18236 1300 18288 1352
rect 18696 1343 18748 1352
rect 18696 1309 18705 1343
rect 18705 1309 18739 1343
rect 18739 1309 18748 1343
rect 18696 1300 18748 1309
rect 19340 1300 19392 1352
rect 20720 1300 20772 1352
rect 22008 1343 22060 1352
rect 22008 1309 22017 1343
rect 22017 1309 22051 1343
rect 22051 1309 22060 1343
rect 22008 1300 22060 1309
rect 22652 1343 22704 1352
rect 22652 1309 22661 1343
rect 22661 1309 22695 1343
rect 22695 1309 22704 1343
rect 22652 1300 22704 1309
rect 22928 1343 22980 1352
rect 22928 1309 22937 1343
rect 22937 1309 22971 1343
rect 22971 1309 22980 1343
rect 22928 1300 22980 1309
rect 23572 1343 23624 1352
rect 23572 1309 23581 1343
rect 23581 1309 23615 1343
rect 23615 1309 23624 1343
rect 23572 1300 23624 1309
rect 24952 1368 25004 1420
rect 25136 1411 25188 1420
rect 25136 1377 25145 1411
rect 25145 1377 25179 1411
rect 25179 1377 25188 1411
rect 25136 1368 25188 1377
rect 26240 1411 26292 1420
rect 26240 1377 26249 1411
rect 26249 1377 26283 1411
rect 26283 1377 26292 1411
rect 26240 1368 26292 1377
rect 31024 1411 31076 1420
rect 24860 1343 24912 1352
rect 24860 1309 24869 1343
rect 24869 1309 24903 1343
rect 24903 1309 24912 1343
rect 24860 1300 24912 1309
rect 25320 1300 25372 1352
rect 27436 1343 27488 1352
rect 27436 1309 27445 1343
rect 27445 1309 27479 1343
rect 27479 1309 27488 1343
rect 28080 1343 28132 1352
rect 27436 1300 27488 1309
rect 28080 1309 28089 1343
rect 28089 1309 28123 1343
rect 28123 1309 28132 1343
rect 28080 1300 28132 1309
rect 9404 1232 9456 1284
rect 11980 1232 12032 1284
rect 3240 1164 3292 1216
rect 5632 1207 5684 1216
rect 5632 1173 5641 1207
rect 5641 1173 5675 1207
rect 5675 1173 5684 1207
rect 5632 1164 5684 1173
rect 9680 1164 9732 1216
rect 12348 1207 12400 1216
rect 12348 1173 12357 1207
rect 12357 1173 12391 1207
rect 12391 1173 12400 1207
rect 12348 1164 12400 1173
rect 13728 1164 13780 1216
rect 14096 1207 14148 1216
rect 14096 1173 14105 1207
rect 14105 1173 14139 1207
rect 14139 1173 14148 1207
rect 14096 1164 14148 1173
rect 16028 1164 16080 1216
rect 17500 1164 17552 1216
rect 19064 1164 19116 1216
rect 19708 1164 19760 1216
rect 20904 1164 20956 1216
rect 23296 1164 23348 1216
rect 26332 1164 26384 1216
rect 28172 1232 28224 1284
rect 28356 1343 28408 1352
rect 28356 1309 28365 1343
rect 28365 1309 28399 1343
rect 28399 1309 28408 1343
rect 28356 1300 28408 1309
rect 29000 1343 29052 1352
rect 29000 1309 29009 1343
rect 29009 1309 29043 1343
rect 29043 1309 29052 1343
rect 29736 1343 29788 1352
rect 29000 1300 29052 1309
rect 29736 1309 29745 1343
rect 29745 1309 29779 1343
rect 29779 1309 29788 1343
rect 29736 1300 29788 1309
rect 31024 1377 31033 1411
rect 31033 1377 31067 1411
rect 31067 1377 31076 1411
rect 31024 1368 31076 1377
rect 30840 1343 30892 1352
rect 30840 1309 30849 1343
rect 30849 1309 30883 1343
rect 30883 1309 30892 1343
rect 30840 1300 30892 1309
rect 31116 1343 31168 1352
rect 31116 1309 31125 1343
rect 31125 1309 31159 1343
rect 31159 1309 31168 1343
rect 31116 1300 31168 1309
rect 28816 1232 28868 1284
rect 7288 1062 7340 1114
rect 17592 1062 17644 1114
rect 27896 1062 27948 1114
rect 5816 960 5868 1012
rect 17408 960 17460 1012
rect 29736 960 29788 1012
rect 8392 892 8444 944
rect 13820 892 13872 944
rect 22008 892 22060 944
rect 24860 892 24912 944
rect 9220 824 9272 876
rect 19616 824 19668 876
rect 24768 824 24820 876
rect 29000 824 29052 876
rect 5632 756 5684 808
rect 6276 688 6328 740
rect 11980 688 12032 740
rect 24308 756 24360 808
rect 27436 756 27488 808
rect 31300 756 31352 808
rect 29092 688 29144 740
rect 28448 620 28500 672
<< metal2 >>
rect 8298 42720 8354 43520
rect 24858 42720 24914 43520
rect 1216 42356 1268 42362
rect 1216 42298 1268 42304
rect 1228 35894 1256 42298
rect 1492 42220 1544 42226
rect 1492 42162 1544 42168
rect 1400 41608 1452 41614
rect 1400 41550 1452 41556
rect 1412 41138 1440 41550
rect 1400 41132 1452 41138
rect 1400 41074 1452 41080
rect 1504 40730 1532 42162
rect 1584 42016 1636 42022
rect 1584 41958 1636 41964
rect 1492 40724 1544 40730
rect 1492 40666 1544 40672
rect 1400 39976 1452 39982
rect 1400 39918 1452 39924
rect 1412 38350 1440 39918
rect 1400 38344 1452 38350
rect 1400 38286 1452 38292
rect 1308 37868 1360 37874
rect 1308 37810 1360 37816
rect 1320 37194 1348 37810
rect 1412 37262 1440 38286
rect 1400 37256 1452 37262
rect 1400 37198 1452 37204
rect 1308 37188 1360 37194
rect 1308 37130 1360 37136
rect 1044 35866 1256 35894
rect 1044 19334 1072 35866
rect 1412 35698 1440 37198
rect 1492 37188 1544 37194
rect 1492 37130 1544 37136
rect 1504 36922 1532 37130
rect 1492 36916 1544 36922
rect 1492 36858 1544 36864
rect 1596 35894 1624 41958
rect 2134 41914 2190 42480
rect 7286 42458 7342 42480
rect 7286 42406 7288 42458
rect 7340 42406 7342 42458
rect 2872 42220 2924 42226
rect 2872 42162 2924 42168
rect 2596 42084 2648 42090
rect 2596 42026 2648 42032
rect 2134 41862 2136 41914
rect 2188 41862 2190 41914
rect 1676 41132 1728 41138
rect 1676 41074 1728 41080
rect 1688 40730 1716 41074
rect 2134 40826 2190 41862
rect 2608 41426 2636 42026
rect 2688 42016 2740 42022
rect 2688 41958 2740 41964
rect 2700 41614 2728 41958
rect 2688 41608 2740 41614
rect 2688 41550 2740 41556
rect 2688 41472 2740 41478
rect 2608 41420 2688 41426
rect 2608 41414 2740 41420
rect 2608 41398 2728 41414
rect 2134 40774 2136 40826
rect 2188 40774 2190 40826
rect 1676 40724 1728 40730
rect 1676 40666 1728 40672
rect 2134 39738 2190 40774
rect 2700 40526 2728 41398
rect 2884 40730 2912 42162
rect 3240 42152 3292 42158
rect 3240 42094 3292 42100
rect 3252 40934 3280 42094
rect 5264 41676 5316 41682
rect 5264 41618 5316 41624
rect 3976 41608 4028 41614
rect 3976 41550 4028 41556
rect 4344 41608 4396 41614
rect 4344 41550 4396 41556
rect 4988 41608 5040 41614
rect 4988 41550 5040 41556
rect 3884 41472 3936 41478
rect 3884 41414 3936 41420
rect 3896 41138 3924 41414
rect 3884 41132 3936 41138
rect 3884 41074 3936 41080
rect 3240 40928 3292 40934
rect 3240 40870 3292 40876
rect 2872 40724 2924 40730
rect 2872 40666 2924 40672
rect 2872 40588 2924 40594
rect 2872 40530 2924 40536
rect 2688 40520 2740 40526
rect 2688 40462 2740 40468
rect 2596 40044 2648 40050
rect 2596 39986 2648 39992
rect 2134 39686 2136 39738
rect 2188 39686 2190 39738
rect 1860 39296 1912 39302
rect 1860 39238 1912 39244
rect 1596 35866 1808 35894
rect 1400 35692 1452 35698
rect 1400 35634 1452 35640
rect 1676 35692 1728 35698
rect 1676 35634 1728 35640
rect 1412 33522 1440 35634
rect 1688 35290 1716 35634
rect 1676 35284 1728 35290
rect 1676 35226 1728 35232
rect 1584 34400 1636 34406
rect 1584 34342 1636 34348
rect 1400 33516 1452 33522
rect 1400 33458 1452 33464
rect 1412 32434 1440 33458
rect 1400 32428 1452 32434
rect 1400 32370 1452 32376
rect 1400 30728 1452 30734
rect 1400 30670 1452 30676
rect 1412 29646 1440 30670
rect 1400 29640 1452 29646
rect 1400 29582 1452 29588
rect 1412 28558 1440 29582
rect 1400 28552 1452 28558
rect 1400 28494 1452 28500
rect 1596 27962 1624 34342
rect 1676 33516 1728 33522
rect 1676 33458 1728 33464
rect 1688 33114 1716 33458
rect 1676 33108 1728 33114
rect 1676 33050 1728 33056
rect 1780 31278 1808 35866
rect 1768 31272 1820 31278
rect 1768 31214 1820 31220
rect 1768 31136 1820 31142
rect 1768 31078 1820 31084
rect 1780 30734 1808 31078
rect 1768 30728 1820 30734
rect 1768 30670 1820 30676
rect 1596 27934 1808 27962
rect 1400 27872 1452 27878
rect 1400 27814 1452 27820
rect 1412 27010 1440 27814
rect 1584 27532 1636 27538
rect 1584 27474 1636 27480
rect 1320 26982 1440 27010
rect 1320 25974 1348 26982
rect 1400 26920 1452 26926
rect 1400 26862 1452 26868
rect 1308 25968 1360 25974
rect 1308 25910 1360 25916
rect 1412 25770 1440 26862
rect 1492 26308 1544 26314
rect 1492 26250 1544 26256
rect 1400 25764 1452 25770
rect 1400 25706 1452 25712
rect 1308 23860 1360 23866
rect 1308 23802 1360 23808
rect 1320 23610 1348 23802
rect 1412 23730 1440 25706
rect 1504 25294 1532 26250
rect 1596 25702 1624 27474
rect 1676 26988 1728 26994
rect 1676 26930 1728 26936
rect 1688 26042 1716 26930
rect 1780 26790 1808 27934
rect 1872 27130 1900 39238
rect 2134 38650 2190 39686
rect 2608 39642 2636 39986
rect 2596 39636 2648 39642
rect 2596 39578 2648 39584
rect 2700 39506 2728 40462
rect 2884 39846 2912 40530
rect 3252 40526 3280 40870
rect 3240 40520 3292 40526
rect 3240 40462 3292 40468
rect 3516 40520 3568 40526
rect 3516 40462 3568 40468
rect 2872 39840 2924 39846
rect 2872 39782 2924 39788
rect 3252 39506 3280 40462
rect 3528 40050 3556 40462
rect 3988 40186 4016 41550
rect 4068 41472 4120 41478
rect 4068 41414 4120 41420
rect 4080 40526 4108 41414
rect 4356 40526 4384 41550
rect 4436 41200 4488 41206
rect 4436 41142 4488 41148
rect 4068 40520 4120 40526
rect 4068 40462 4120 40468
rect 4344 40520 4396 40526
rect 4344 40462 4396 40468
rect 3976 40180 4028 40186
rect 3976 40122 4028 40128
rect 4448 40050 4476 41142
rect 5000 40594 5028 41550
rect 5276 40934 5304 41618
rect 5356 41608 5408 41614
rect 5356 41550 5408 41556
rect 7012 41608 7064 41614
rect 7012 41550 7064 41556
rect 5264 40928 5316 40934
rect 5264 40870 5316 40876
rect 4620 40588 4672 40594
rect 4620 40530 4672 40536
rect 4988 40588 5040 40594
rect 4988 40530 5040 40536
rect 3516 40044 3568 40050
rect 3516 39986 3568 39992
rect 4436 40044 4488 40050
rect 4436 39986 4488 39992
rect 4528 40044 4580 40050
rect 4632 40032 4660 40530
rect 5172 40520 5224 40526
rect 5172 40462 5224 40468
rect 4580 40004 4660 40032
rect 4528 39986 4580 39992
rect 2688 39500 2740 39506
rect 2688 39442 2740 39448
rect 3240 39500 3292 39506
rect 3240 39442 3292 39448
rect 2412 38956 2464 38962
rect 2412 38898 2464 38904
rect 2228 38752 2280 38758
rect 2228 38694 2280 38700
rect 2134 38598 2136 38650
rect 2188 38598 2190 38650
rect 2134 37562 2190 38598
rect 2240 38282 2268 38694
rect 2228 38276 2280 38282
rect 2228 38218 2280 38224
rect 2424 38010 2452 38898
rect 2700 38758 2728 39442
rect 2780 39432 2832 39438
rect 2780 39374 2832 39380
rect 3056 39432 3108 39438
rect 3056 39374 3108 39380
rect 2792 39098 2820 39374
rect 2780 39092 2832 39098
rect 2780 39034 2832 39040
rect 2780 38888 2832 38894
rect 2780 38830 2832 38836
rect 2688 38752 2740 38758
rect 2688 38694 2740 38700
rect 2792 38332 2820 38830
rect 3068 38554 3096 39374
rect 3528 39098 3556 39986
rect 3792 39840 3844 39846
rect 3792 39782 3844 39788
rect 3804 39370 3832 39782
rect 4252 39432 4304 39438
rect 4252 39374 4304 39380
rect 3792 39364 3844 39370
rect 3792 39306 3844 39312
rect 3516 39092 3568 39098
rect 3516 39034 3568 39040
rect 3804 38962 3832 39306
rect 3792 38956 3844 38962
rect 3792 38898 3844 38904
rect 3056 38548 3108 38554
rect 3056 38490 3108 38496
rect 2872 38344 2924 38350
rect 2792 38304 2872 38332
rect 2412 38004 2464 38010
rect 2412 37946 2464 37952
rect 2320 37664 2372 37670
rect 2320 37606 2372 37612
rect 2134 37510 2136 37562
rect 2188 37510 2190 37562
rect 2134 36474 2190 37510
rect 2228 36576 2280 36582
rect 2228 36518 2280 36524
rect 2134 36422 2136 36474
rect 2188 36422 2190 36474
rect 2044 36032 2096 36038
rect 2044 35974 2096 35980
rect 2056 35086 2084 35974
rect 2134 35386 2190 36422
rect 2240 35766 2268 36518
rect 2228 35760 2280 35766
rect 2228 35702 2280 35708
rect 2134 35334 2136 35386
rect 2188 35334 2190 35386
rect 2044 35080 2096 35086
rect 2044 35022 2096 35028
rect 1952 35012 2004 35018
rect 1952 34954 2004 34960
rect 1964 34202 1992 34954
rect 2134 34298 2190 35334
rect 2240 35290 2268 35702
rect 2228 35284 2280 35290
rect 2228 35226 2280 35232
rect 2134 34246 2136 34298
rect 2188 34246 2190 34298
rect 1952 34196 2004 34202
rect 1952 34138 2004 34144
rect 2134 33210 2190 34246
rect 2240 34202 2268 35226
rect 2228 34196 2280 34202
rect 2228 34138 2280 34144
rect 2134 33158 2136 33210
rect 2188 33158 2190 33210
rect 2134 32122 2190 33158
rect 2134 32070 2136 32122
rect 2188 32070 2190 32122
rect 2044 31816 2096 31822
rect 2044 31758 2096 31764
rect 2056 31414 2084 31758
rect 2044 31408 2096 31414
rect 2044 31350 2096 31356
rect 2044 31272 2096 31278
rect 2044 31214 2096 31220
rect 1952 28212 2004 28218
rect 1952 28154 2004 28160
rect 1860 27124 1912 27130
rect 1860 27066 1912 27072
rect 1768 26784 1820 26790
rect 1768 26726 1820 26732
rect 1860 26376 1912 26382
rect 1860 26318 1912 26324
rect 1768 26240 1820 26246
rect 1768 26182 1820 26188
rect 1676 26036 1728 26042
rect 1676 25978 1728 25984
rect 1780 25906 1808 26182
rect 1872 25906 1900 26318
rect 1768 25900 1820 25906
rect 1768 25842 1820 25848
rect 1860 25900 1912 25906
rect 1860 25842 1912 25848
rect 1676 25832 1728 25838
rect 1676 25774 1728 25780
rect 1584 25696 1636 25702
rect 1584 25638 1636 25644
rect 1492 25288 1544 25294
rect 1492 25230 1544 25236
rect 1492 25152 1544 25158
rect 1492 25094 1544 25100
rect 1504 23866 1532 25094
rect 1596 24154 1624 25638
rect 1688 24886 1716 25774
rect 1768 25152 1820 25158
rect 1768 25094 1820 25100
rect 1676 24880 1728 24886
rect 1676 24822 1728 24828
rect 1688 24274 1716 24822
rect 1676 24268 1728 24274
rect 1676 24210 1728 24216
rect 1596 24126 1716 24154
rect 1584 24064 1636 24070
rect 1584 24006 1636 24012
rect 1492 23860 1544 23866
rect 1492 23802 1544 23808
rect 1400 23724 1452 23730
rect 1400 23666 1452 23672
rect 1492 23724 1544 23730
rect 1492 23666 1544 23672
rect 1320 23582 1440 23610
rect 1412 21842 1440 23582
rect 1504 22778 1532 23666
rect 1492 22772 1544 22778
rect 1492 22714 1544 22720
rect 1412 21814 1532 21842
rect 1400 21684 1452 21690
rect 1400 21626 1452 21632
rect 1308 19848 1360 19854
rect 1308 19790 1360 19796
rect 1124 19780 1176 19786
rect 1124 19722 1176 19728
rect 952 19306 1072 19334
rect 952 17814 980 19306
rect 1136 18714 1164 19722
rect 1320 19174 1348 19790
rect 1308 19168 1360 19174
rect 1308 19110 1360 19116
rect 1044 18686 1164 18714
rect 940 17808 992 17814
rect 940 17750 992 17756
rect 1044 15026 1072 18686
rect 1412 16130 1440 21626
rect 1504 17610 1532 21814
rect 1596 19718 1624 24006
rect 1688 22778 1716 24126
rect 1676 22772 1728 22778
rect 1676 22714 1728 22720
rect 1676 22636 1728 22642
rect 1676 22578 1728 22584
rect 1688 22234 1716 22578
rect 1676 22228 1728 22234
rect 1676 22170 1728 22176
rect 1676 21344 1728 21350
rect 1676 21286 1728 21292
rect 1688 20534 1716 21286
rect 1676 20528 1728 20534
rect 1676 20470 1728 20476
rect 1688 19786 1716 20470
rect 1676 19780 1728 19786
rect 1676 19722 1728 19728
rect 1584 19712 1636 19718
rect 1584 19654 1636 19660
rect 1584 19440 1636 19446
rect 1584 19382 1636 19388
rect 1492 17604 1544 17610
rect 1492 17546 1544 17552
rect 1492 16448 1544 16454
rect 1492 16390 1544 16396
rect 1136 16102 1440 16130
rect 1032 15020 1084 15026
rect 1032 14962 1084 14968
rect 1136 10266 1164 16102
rect 1400 16040 1452 16046
rect 1400 15982 1452 15988
rect 1412 14414 1440 15982
rect 1504 15706 1532 16390
rect 1492 15700 1544 15706
rect 1492 15642 1544 15648
rect 1492 15428 1544 15434
rect 1492 15370 1544 15376
rect 1504 15094 1532 15370
rect 1492 15088 1544 15094
rect 1492 15030 1544 15036
rect 1400 14408 1452 14414
rect 1400 14350 1452 14356
rect 1308 13932 1360 13938
rect 1308 13874 1360 13880
rect 1320 12782 1348 13874
rect 1308 12776 1360 12782
rect 1308 12718 1360 12724
rect 1320 11914 1348 12718
rect 1412 12238 1440 14350
rect 1492 13388 1544 13394
rect 1492 13330 1544 13336
rect 1504 12918 1532 13330
rect 1492 12912 1544 12918
rect 1492 12854 1544 12860
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1228 11886 1348 11914
rect 1124 10260 1176 10266
rect 1124 10202 1176 10208
rect 1228 6322 1256 11886
rect 1596 11778 1624 19382
rect 1676 19372 1728 19378
rect 1676 19314 1728 19320
rect 1688 18426 1716 19314
rect 1676 18420 1728 18426
rect 1676 18362 1728 18368
rect 1780 17082 1808 25094
rect 1872 22030 1900 25842
rect 1964 24682 1992 28154
rect 1952 24676 2004 24682
rect 1952 24618 2004 24624
rect 1860 22024 1912 22030
rect 1860 21966 1912 21972
rect 1860 20868 1912 20874
rect 1860 20810 1912 20816
rect 1872 20602 1900 20810
rect 1860 20596 1912 20602
rect 1860 20538 1912 20544
rect 1964 19530 1992 24618
rect 2056 20602 2084 31214
rect 2134 31034 2190 32070
rect 2134 30982 2136 31034
rect 2188 30982 2190 31034
rect 2134 29946 2190 30982
rect 2134 29894 2136 29946
rect 2188 29894 2190 29946
rect 2134 28858 2190 29894
rect 2228 28960 2280 28966
rect 2228 28902 2280 28908
rect 2134 28806 2136 28858
rect 2188 28806 2190 28858
rect 2134 27770 2190 28806
rect 2240 28490 2268 28902
rect 2228 28484 2280 28490
rect 2228 28426 2280 28432
rect 2332 28014 2360 37606
rect 2792 37466 2820 38304
rect 2872 38286 2924 38292
rect 3068 37942 3096 38490
rect 3056 37936 3108 37942
rect 3056 37878 3108 37884
rect 4264 37874 4292 39374
rect 4448 38486 4476 39986
rect 4632 39506 4660 40004
rect 4620 39500 4672 39506
rect 4620 39442 4672 39448
rect 4632 39030 4660 39442
rect 4620 39024 4672 39030
rect 4620 38966 4672 38972
rect 5184 38962 5212 40462
rect 5276 40118 5304 40870
rect 5368 40594 5396 41550
rect 5816 41472 5868 41478
rect 5816 41414 5868 41420
rect 5356 40588 5408 40594
rect 5356 40530 5408 40536
rect 5368 40186 5396 40530
rect 5356 40180 5408 40186
rect 5356 40122 5408 40128
rect 5264 40112 5316 40118
rect 5264 40054 5316 40060
rect 5172 38956 5224 38962
rect 5172 38898 5224 38904
rect 5276 38894 5304 40054
rect 5828 40050 5856 41414
rect 7024 41206 7052 41550
rect 7286 41370 7342 42406
rect 8312 42378 8340 42720
rect 8220 42362 8340 42378
rect 8208 42356 8340 42362
rect 8260 42350 8340 42356
rect 8208 42298 8260 42304
rect 7656 42220 7708 42226
rect 7656 42162 7708 42168
rect 8116 42220 8168 42226
rect 8116 42162 8168 42168
rect 9128 42220 9180 42226
rect 9128 42162 9180 42168
rect 10232 42220 10284 42226
rect 10232 42162 10284 42168
rect 7668 41414 7696 42162
rect 7286 41318 7288 41370
rect 7340 41318 7342 41370
rect 7012 41200 7064 41206
rect 7012 41142 7064 41148
rect 6920 41132 6972 41138
rect 6920 41074 6972 41080
rect 6932 40662 6960 41074
rect 7024 40730 7052 41142
rect 7012 40724 7064 40730
rect 7012 40666 7064 40672
rect 6920 40656 6972 40662
rect 6920 40598 6972 40604
rect 7286 40282 7342 41318
rect 7286 40230 7288 40282
rect 7340 40230 7342 40282
rect 5816 40044 5868 40050
rect 5816 39986 5868 39992
rect 6736 40044 6788 40050
rect 7104 40044 7156 40050
rect 6788 40004 6868 40032
rect 6736 39986 6788 39992
rect 5908 39840 5960 39846
rect 5908 39782 5960 39788
rect 5448 39296 5500 39302
rect 5448 39238 5500 39244
rect 5356 38956 5408 38962
rect 5356 38898 5408 38904
rect 5264 38888 5316 38894
rect 5264 38830 5316 38836
rect 5368 38486 5396 38898
rect 5460 38554 5488 39238
rect 5920 39030 5948 39782
rect 6840 39386 6868 40004
rect 7104 39986 7156 39992
rect 7116 39438 7144 39986
rect 7196 39840 7248 39846
rect 7196 39782 7248 39788
rect 7208 39642 7236 39782
rect 7196 39636 7248 39642
rect 7196 39578 7248 39584
rect 6656 39370 6868 39386
rect 7104 39432 7156 39438
rect 7104 39374 7156 39380
rect 6644 39364 6880 39370
rect 6696 39358 6828 39364
rect 6644 39306 6696 39312
rect 6828 39306 6880 39312
rect 5908 39024 5960 39030
rect 5908 38966 5960 38972
rect 5632 38956 5684 38962
rect 5632 38898 5684 38904
rect 6552 38956 6604 38962
rect 6552 38898 6604 38904
rect 5448 38548 5500 38554
rect 5448 38490 5500 38496
rect 4436 38480 4488 38486
rect 4436 38422 4488 38428
rect 4528 38480 4580 38486
rect 4528 38422 4580 38428
rect 5356 38480 5408 38486
rect 5356 38422 5408 38428
rect 4436 38344 4488 38350
rect 4436 38286 4488 38292
rect 4448 37942 4476 38286
rect 4540 38282 4568 38422
rect 4528 38276 4580 38282
rect 4528 38218 4580 38224
rect 4436 37936 4488 37942
rect 4436 37878 4488 37884
rect 4252 37868 4304 37874
rect 4252 37810 4304 37816
rect 4160 37800 4212 37806
rect 4160 37742 4212 37748
rect 3792 37664 3844 37670
rect 3792 37606 3844 37612
rect 2780 37460 2832 37466
rect 2780 37402 2832 37408
rect 2792 36768 2820 37402
rect 3240 37188 3292 37194
rect 3240 37130 3292 37136
rect 2872 36780 2924 36786
rect 2792 36740 2872 36768
rect 2872 36722 2924 36728
rect 3252 36718 3280 37130
rect 3804 36922 3832 37606
rect 3792 36916 3844 36922
rect 3792 36858 3844 36864
rect 3804 36786 3832 36858
rect 4172 36786 4200 37742
rect 4344 37256 4396 37262
rect 4344 37198 4396 37204
rect 4356 36922 4384 37198
rect 4712 37188 4764 37194
rect 4712 37130 4764 37136
rect 4344 36916 4396 36922
rect 4344 36858 4396 36864
rect 3792 36780 3844 36786
rect 3792 36722 3844 36728
rect 4160 36780 4212 36786
rect 4160 36722 4212 36728
rect 4344 36780 4396 36786
rect 4344 36722 4396 36728
rect 4620 36780 4672 36786
rect 4620 36722 4672 36728
rect 3240 36712 3292 36718
rect 3240 36654 3292 36660
rect 2412 36576 2464 36582
rect 2412 36518 2464 36524
rect 2424 33930 2452 36518
rect 2504 36372 2556 36378
rect 2504 36314 2556 36320
rect 2516 34066 2544 36314
rect 2596 36304 2648 36310
rect 2596 36246 2648 36252
rect 2504 34060 2556 34066
rect 2504 34002 2556 34008
rect 2412 33924 2464 33930
rect 2412 33866 2464 33872
rect 2504 32904 2556 32910
rect 2504 32846 2556 32852
rect 2412 32428 2464 32434
rect 2412 32370 2464 32376
rect 2424 32026 2452 32370
rect 2516 32298 2544 32846
rect 2504 32292 2556 32298
rect 2504 32234 2556 32240
rect 2412 32020 2464 32026
rect 2412 31962 2464 31968
rect 2608 31754 2636 36246
rect 3252 36174 3280 36654
rect 3332 36644 3384 36650
rect 3332 36586 3384 36592
rect 3240 36168 3292 36174
rect 3240 36110 3292 36116
rect 2964 36032 3016 36038
rect 2964 35974 3016 35980
rect 2688 35148 2740 35154
rect 2688 35090 2740 35096
rect 2700 34474 2728 35090
rect 2976 35086 3004 35974
rect 3252 35834 3280 36110
rect 3240 35828 3292 35834
rect 3240 35770 3292 35776
rect 3344 35766 3372 36586
rect 3804 36174 3832 36722
rect 4172 36174 4200 36722
rect 3792 36168 3844 36174
rect 3792 36110 3844 36116
rect 4160 36168 4212 36174
rect 4160 36110 4212 36116
rect 3332 35760 3384 35766
rect 3332 35702 3384 35708
rect 3792 35488 3844 35494
rect 3792 35430 3844 35436
rect 3804 35154 3832 35430
rect 3792 35148 3844 35154
rect 3792 35090 3844 35096
rect 4356 35086 4384 36722
rect 4632 36378 4660 36722
rect 4620 36372 4672 36378
rect 4620 36314 4672 36320
rect 4632 36038 4660 36314
rect 4724 36174 4752 37130
rect 5368 36718 5396 38422
rect 5448 38412 5500 38418
rect 5448 38354 5500 38360
rect 5460 37806 5488 38354
rect 5540 38344 5592 38350
rect 5540 38286 5592 38292
rect 5552 38010 5580 38286
rect 5540 38004 5592 38010
rect 5540 37946 5592 37952
rect 5644 37942 5672 38898
rect 5724 38752 5776 38758
rect 5724 38694 5776 38700
rect 5632 37936 5684 37942
rect 5632 37878 5684 37884
rect 5540 37868 5592 37874
rect 5540 37810 5592 37816
rect 5448 37800 5500 37806
rect 5448 37742 5500 37748
rect 5356 36712 5408 36718
rect 5356 36654 5408 36660
rect 5460 36242 5488 37742
rect 5552 37738 5580 37810
rect 5540 37732 5592 37738
rect 5540 37674 5592 37680
rect 5644 36786 5672 37878
rect 5736 37262 5764 38694
rect 6564 38554 6592 38898
rect 6552 38548 6604 38554
rect 6552 38490 6604 38496
rect 6564 37874 6592 38490
rect 5816 37868 5868 37874
rect 5816 37810 5868 37816
rect 6552 37868 6604 37874
rect 6552 37810 6604 37816
rect 5724 37256 5776 37262
rect 5724 37198 5776 37204
rect 5632 36780 5684 36786
rect 5632 36722 5684 36728
rect 5448 36236 5500 36242
rect 5448 36178 5500 36184
rect 4712 36168 4764 36174
rect 4712 36110 4764 36116
rect 5172 36168 5224 36174
rect 5172 36110 5224 36116
rect 4620 36032 4672 36038
rect 4620 35974 4672 35980
rect 5184 35306 5212 36110
rect 5092 35290 5212 35306
rect 5080 35284 5212 35290
rect 5132 35278 5212 35284
rect 5080 35226 5132 35232
rect 2964 35080 3016 35086
rect 2964 35022 3016 35028
rect 4344 35080 4396 35086
rect 4344 35022 4396 35028
rect 2780 34944 2832 34950
rect 2780 34886 2832 34892
rect 2792 34678 2820 34886
rect 5184 34746 5212 35278
rect 5172 34740 5224 34746
rect 5172 34682 5224 34688
rect 2780 34672 2832 34678
rect 2780 34614 2832 34620
rect 5828 34610 5856 37810
rect 6092 37732 6144 37738
rect 6092 37674 6144 37680
rect 6104 37330 6132 37674
rect 6840 37398 6868 39306
rect 6828 37392 6880 37398
rect 6828 37334 6880 37340
rect 6092 37324 6144 37330
rect 6092 37266 6144 37272
rect 6104 36258 6132 37266
rect 6460 37256 6512 37262
rect 6460 37198 6512 37204
rect 6276 37120 6328 37126
rect 6276 37062 6328 37068
rect 6288 36378 6316 37062
rect 6368 36576 6420 36582
rect 6368 36518 6420 36524
rect 6276 36372 6328 36378
rect 6276 36314 6328 36320
rect 6104 36230 6224 36258
rect 5080 34604 5132 34610
rect 5080 34546 5132 34552
rect 5632 34604 5684 34610
rect 5632 34546 5684 34552
rect 5816 34604 5868 34610
rect 5816 34546 5868 34552
rect 2688 34468 2740 34474
rect 2688 34410 2740 34416
rect 2700 33590 2728 34410
rect 2872 34400 2924 34406
rect 2872 34342 2924 34348
rect 3148 34400 3200 34406
rect 3148 34342 3200 34348
rect 2780 34060 2832 34066
rect 2780 34002 2832 34008
rect 2688 33584 2740 33590
rect 2688 33526 2740 33532
rect 2792 33046 2820 34002
rect 2884 33930 2912 34342
rect 3160 34066 3188 34342
rect 3148 34060 3200 34066
rect 3148 34002 3200 34008
rect 2964 33992 3016 33998
rect 2964 33934 3016 33940
rect 3240 33992 3292 33998
rect 3240 33934 3292 33940
rect 4436 33992 4488 33998
rect 4436 33934 4488 33940
rect 2872 33924 2924 33930
rect 2872 33866 2924 33872
rect 2872 33312 2924 33318
rect 2872 33254 2924 33260
rect 2884 33114 2912 33254
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2780 33040 2832 33046
rect 2780 32982 2832 32988
rect 2688 32224 2740 32230
rect 2688 32166 2740 32172
rect 2700 31822 2728 32166
rect 2792 31958 2820 32982
rect 2976 32026 3004 33934
rect 3252 33114 3280 33934
rect 3332 33856 3384 33862
rect 3332 33798 3384 33804
rect 3344 33522 3372 33798
rect 4448 33590 4476 33934
rect 5092 33658 5120 34546
rect 5080 33652 5132 33658
rect 5080 33594 5132 33600
rect 4436 33584 4488 33590
rect 4436 33526 4488 33532
rect 5448 33584 5500 33590
rect 5448 33526 5500 33532
rect 3332 33516 3384 33522
rect 3332 33458 3384 33464
rect 3240 33108 3292 33114
rect 3240 33050 3292 33056
rect 4160 33040 4212 33046
rect 4160 32982 4212 32988
rect 3424 32972 3476 32978
rect 3424 32914 3476 32920
rect 3056 32904 3108 32910
rect 3056 32846 3108 32852
rect 3068 32502 3096 32846
rect 3056 32496 3108 32502
rect 3056 32438 3108 32444
rect 3436 32434 3464 32914
rect 3976 32904 4028 32910
rect 3976 32846 4028 32852
rect 3988 32774 4016 32846
rect 3976 32768 4028 32774
rect 3976 32710 4028 32716
rect 3424 32428 3476 32434
rect 3424 32370 3476 32376
rect 2964 32020 3016 32026
rect 2964 31962 3016 31968
rect 2780 31952 2832 31958
rect 2780 31894 2832 31900
rect 2688 31816 2740 31822
rect 2688 31758 2740 31764
rect 2872 31816 2924 31822
rect 2872 31758 2924 31764
rect 2424 31726 2636 31754
rect 2424 28218 2452 31726
rect 2504 31408 2556 31414
rect 2504 31350 2556 31356
rect 2412 28212 2464 28218
rect 2412 28154 2464 28160
rect 2412 28076 2464 28082
rect 2412 28018 2464 28024
rect 2320 28008 2372 28014
rect 2320 27950 2372 27956
rect 2320 27872 2372 27878
rect 2320 27814 2372 27820
rect 2134 27718 2136 27770
rect 2188 27718 2190 27770
rect 2134 26682 2190 27718
rect 2134 26630 2136 26682
rect 2188 26630 2190 26682
rect 2134 25594 2190 26630
rect 2228 26036 2280 26042
rect 2228 25978 2280 25984
rect 2134 25542 2136 25594
rect 2188 25542 2190 25594
rect 2134 24506 2190 25542
rect 2240 25362 2268 25978
rect 2228 25356 2280 25362
rect 2228 25298 2280 25304
rect 2228 25220 2280 25226
rect 2228 25162 2280 25168
rect 2240 24954 2268 25162
rect 2228 24948 2280 24954
rect 2228 24890 2280 24896
rect 2228 24812 2280 24818
rect 2228 24754 2280 24760
rect 2134 24454 2136 24506
rect 2188 24454 2190 24506
rect 2134 23418 2190 24454
rect 2240 23730 2268 24754
rect 2228 23724 2280 23730
rect 2228 23666 2280 23672
rect 2134 23366 2136 23418
rect 2188 23366 2190 23418
rect 2134 22330 2190 23366
rect 2228 23044 2280 23050
rect 2228 22986 2280 22992
rect 2240 22506 2268 22986
rect 2228 22500 2280 22506
rect 2228 22442 2280 22448
rect 2134 22278 2136 22330
rect 2188 22278 2190 22330
rect 2134 21242 2190 22278
rect 2228 22024 2280 22030
rect 2228 21966 2280 21972
rect 2134 21190 2136 21242
rect 2188 21190 2190 21242
rect 2044 20596 2096 20602
rect 2044 20538 2096 20544
rect 2044 20460 2096 20466
rect 2044 20402 2096 20408
rect 2056 20058 2084 20402
rect 2134 20154 2190 21190
rect 2240 20466 2268 21966
rect 2332 21690 2360 27814
rect 2320 21684 2372 21690
rect 2320 21626 2372 21632
rect 2320 21344 2372 21350
rect 2320 21286 2372 21292
rect 2228 20460 2280 20466
rect 2228 20402 2280 20408
rect 2228 20256 2280 20262
rect 2228 20198 2280 20204
rect 2134 20102 2136 20154
rect 2188 20102 2190 20154
rect 2044 20052 2096 20058
rect 2044 19994 2096 20000
rect 1872 19502 1992 19530
rect 1872 19446 1900 19502
rect 1860 19440 1912 19446
rect 1860 19382 1912 19388
rect 1952 19372 2004 19378
rect 1952 19314 2004 19320
rect 1964 18834 1992 19314
rect 2134 19066 2190 20102
rect 2134 19014 2136 19066
rect 2188 19014 2190 19066
rect 1952 18828 2004 18834
rect 1952 18770 2004 18776
rect 1952 18624 2004 18630
rect 1952 18566 2004 18572
rect 1964 18290 1992 18566
rect 1952 18284 2004 18290
rect 1952 18226 2004 18232
rect 2134 17978 2190 19014
rect 2240 18358 2268 20198
rect 2228 18352 2280 18358
rect 2228 18294 2280 18300
rect 2228 18080 2280 18086
rect 2228 18022 2280 18028
rect 2134 17926 2136 17978
rect 2188 17926 2190 17978
rect 2044 17536 2096 17542
rect 2044 17478 2096 17484
rect 1688 17054 1808 17082
rect 1860 17060 1912 17066
rect 1688 15162 1716 17054
rect 1860 17002 1912 17008
rect 1768 16992 1820 16998
rect 1768 16934 1820 16940
rect 1676 15156 1728 15162
rect 1676 15098 1728 15104
rect 1676 15020 1728 15026
rect 1676 14962 1728 14968
rect 1504 11750 1624 11778
rect 1504 10690 1532 11750
rect 1584 11688 1636 11694
rect 1584 11630 1636 11636
rect 1320 10662 1532 10690
rect 1320 9738 1348 10662
rect 1492 10600 1544 10606
rect 1492 10542 1544 10548
rect 1320 9710 1440 9738
rect 1412 9674 1440 9710
rect 1320 9646 1440 9674
rect 1320 7002 1348 9646
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1412 7954 1440 9522
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 1308 6996 1360 7002
rect 1308 6938 1360 6944
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1216 6316 1268 6322
rect 1216 6258 1268 6264
rect 1412 5098 1440 6734
rect 1504 6254 1532 10542
rect 1492 6248 1544 6254
rect 1492 6190 1544 6196
rect 1492 6112 1544 6118
rect 1492 6054 1544 6060
rect 1504 5914 1532 6054
rect 1492 5908 1544 5914
rect 1492 5850 1544 5856
rect 1400 5092 1452 5098
rect 1400 5034 1452 5040
rect 1412 4690 1440 5034
rect 1596 4826 1624 11630
rect 1688 8974 1716 14962
rect 1780 11626 1808 16934
rect 1872 16046 1900 17002
rect 2056 16590 2084 17478
rect 2134 16890 2190 17926
rect 2134 16838 2136 16890
rect 2188 16838 2190 16890
rect 2044 16584 2096 16590
rect 2044 16526 2096 16532
rect 2044 16448 2096 16454
rect 2044 16390 2096 16396
rect 1860 16040 1912 16046
rect 1860 15982 1912 15988
rect 1860 15904 1912 15910
rect 1860 15846 1912 15852
rect 1872 15502 1900 15846
rect 1860 15496 1912 15502
rect 1860 15438 1912 15444
rect 1952 14952 2004 14958
rect 1952 14894 2004 14900
rect 1860 14816 1912 14822
rect 1860 14758 1912 14764
rect 1872 14074 1900 14758
rect 1860 14068 1912 14074
rect 1860 14010 1912 14016
rect 1860 12708 1912 12714
rect 1860 12650 1912 12656
rect 1768 11620 1820 11626
rect 1768 11562 1820 11568
rect 1872 11150 1900 12650
rect 1964 11762 1992 14894
rect 1952 11756 2004 11762
rect 1952 11698 2004 11704
rect 2056 11234 2084 16390
rect 1964 11206 2084 11234
rect 2134 15802 2190 16838
rect 2240 16182 2268 18022
rect 2332 16266 2360 21286
rect 2424 16454 2452 28018
rect 2516 26450 2544 31350
rect 2596 31340 2648 31346
rect 2596 31282 2648 31288
rect 2608 30394 2636 31282
rect 2884 30870 2912 31758
rect 3884 31476 3936 31482
rect 3884 31418 3936 31424
rect 3608 31272 3660 31278
rect 3608 31214 3660 31220
rect 2872 30864 2924 30870
rect 2872 30806 2924 30812
rect 2596 30388 2648 30394
rect 2596 30330 2648 30336
rect 2884 30258 2912 30806
rect 3620 30258 3648 31214
rect 3700 31136 3752 31142
rect 3700 31078 3752 31084
rect 3712 30734 3740 31078
rect 3700 30728 3752 30734
rect 3700 30670 3752 30676
rect 3712 30326 3740 30670
rect 3700 30320 3752 30326
rect 3700 30262 3752 30268
rect 2872 30252 2924 30258
rect 2872 30194 2924 30200
rect 3608 30252 3660 30258
rect 3608 30194 3660 30200
rect 2780 30048 2832 30054
rect 2780 29990 2832 29996
rect 2596 29572 2648 29578
rect 2596 29514 2648 29520
rect 2608 27606 2636 29514
rect 2688 28552 2740 28558
rect 2688 28494 2740 28500
rect 2700 27878 2728 28494
rect 2688 27872 2740 27878
rect 2688 27814 2740 27820
rect 2596 27600 2648 27606
rect 2596 27542 2648 27548
rect 2596 27124 2648 27130
rect 2596 27066 2648 27072
rect 2504 26444 2556 26450
rect 2504 26386 2556 26392
rect 2608 24886 2636 27066
rect 2700 27062 2728 27814
rect 2792 27470 2820 29990
rect 3620 29850 3648 30194
rect 3608 29844 3660 29850
rect 3608 29786 3660 29792
rect 3148 29708 3200 29714
rect 3148 29650 3200 29656
rect 3160 29306 3188 29650
rect 3712 29646 3740 30262
rect 3700 29640 3752 29646
rect 3700 29582 3752 29588
rect 3148 29300 3200 29306
rect 3148 29242 3200 29248
rect 3712 29238 3740 29582
rect 3700 29232 3752 29238
rect 3700 29174 3752 29180
rect 3792 29164 3844 29170
rect 3792 29106 3844 29112
rect 3804 28694 3832 29106
rect 3056 28688 3108 28694
rect 3056 28630 3108 28636
rect 3792 28688 3844 28694
rect 3792 28630 3844 28636
rect 3068 27538 3096 28630
rect 3896 27554 3924 31418
rect 3988 31346 4016 32710
rect 4068 31952 4120 31958
rect 4068 31894 4120 31900
rect 3976 31340 4028 31346
rect 3976 31282 4028 31288
rect 4080 31278 4108 31894
rect 4172 31822 4200 32982
rect 4252 32496 4304 32502
rect 4252 32438 4304 32444
rect 4264 31822 4292 32438
rect 4448 32434 4476 33526
rect 5356 33516 5408 33522
rect 5356 33458 5408 33464
rect 4712 33380 4764 33386
rect 4712 33322 4764 33328
rect 4620 33312 4672 33318
rect 4620 33254 4672 33260
rect 4632 32978 4660 33254
rect 4620 32972 4672 32978
rect 4620 32914 4672 32920
rect 4528 32904 4580 32910
rect 4528 32846 4580 32852
rect 4540 32502 4568 32846
rect 4528 32496 4580 32502
rect 4528 32438 4580 32444
rect 4436 32428 4488 32434
rect 4436 32370 4488 32376
rect 4632 31822 4660 32914
rect 4724 32910 4752 33322
rect 5368 33046 5396 33458
rect 5356 33040 5408 33046
rect 5356 32982 5408 32988
rect 4712 32904 4764 32910
rect 4712 32846 4764 32852
rect 5368 32858 5396 32982
rect 5460 32978 5488 33526
rect 5448 32972 5500 32978
rect 5448 32914 5500 32920
rect 5368 32830 5488 32858
rect 4988 32428 5040 32434
rect 4988 32370 5040 32376
rect 5000 31890 5028 32370
rect 5460 32366 5488 32830
rect 5644 32570 5672 34546
rect 5724 34196 5776 34202
rect 5724 34138 5776 34144
rect 5736 33522 5764 34138
rect 5724 33516 5776 33522
rect 5724 33458 5776 33464
rect 5828 32842 5856 34546
rect 5908 32904 5960 32910
rect 5908 32846 5960 32852
rect 6092 32904 6144 32910
rect 6092 32846 6144 32852
rect 5816 32836 5868 32842
rect 5816 32778 5868 32784
rect 5724 32768 5776 32774
rect 5724 32710 5776 32716
rect 5632 32564 5684 32570
rect 5632 32506 5684 32512
rect 5448 32360 5500 32366
rect 5448 32302 5500 32308
rect 5644 32230 5672 32506
rect 5736 32502 5764 32710
rect 5920 32570 5948 32846
rect 5908 32564 5960 32570
rect 5908 32506 5960 32512
rect 5724 32496 5776 32502
rect 5724 32438 5776 32444
rect 5632 32224 5684 32230
rect 5632 32166 5684 32172
rect 6104 31890 6132 32846
rect 4988 31884 5040 31890
rect 4988 31826 5040 31832
rect 6092 31884 6144 31890
rect 6092 31826 6144 31832
rect 4160 31816 4212 31822
rect 4160 31758 4212 31764
rect 4252 31816 4304 31822
rect 4252 31758 4304 31764
rect 4620 31816 4672 31822
rect 4620 31758 4672 31764
rect 4252 31340 4304 31346
rect 4252 31282 4304 31288
rect 4068 31272 4120 31278
rect 4068 31214 4120 31220
rect 4264 30938 4292 31282
rect 4804 31272 4856 31278
rect 4804 31214 4856 31220
rect 4344 31136 4396 31142
rect 4344 31078 4396 31084
rect 4252 30932 4304 30938
rect 4252 30874 4304 30880
rect 4160 30660 4212 30666
rect 4160 30602 4212 30608
rect 4172 30122 4200 30602
rect 4356 30326 4384 31078
rect 4344 30320 4396 30326
rect 4344 30262 4396 30268
rect 4252 30184 4304 30190
rect 4252 30126 4304 30132
rect 4160 30116 4212 30122
rect 4160 30058 4212 30064
rect 4172 29578 4200 30058
rect 4264 29782 4292 30126
rect 4252 29776 4304 29782
rect 4252 29718 4304 29724
rect 4160 29572 4212 29578
rect 4160 29514 4212 29520
rect 4172 29102 4200 29514
rect 4264 29170 4292 29718
rect 4816 29646 4844 31214
rect 4896 30728 4948 30734
rect 4896 30670 4948 30676
rect 4908 30054 4936 30670
rect 4896 30048 4948 30054
rect 4896 29990 4948 29996
rect 4804 29640 4856 29646
rect 4804 29582 4856 29588
rect 4344 29504 4396 29510
rect 4344 29446 4396 29452
rect 4252 29164 4304 29170
rect 4252 29106 4304 29112
rect 4160 29096 4212 29102
rect 4160 29038 4212 29044
rect 4356 28558 4384 29446
rect 4816 29306 4844 29582
rect 4804 29300 4856 29306
rect 4804 29242 4856 29248
rect 4908 29238 4936 29990
rect 5000 29646 5028 31826
rect 6196 31754 6224 36230
rect 6380 34678 6408 36518
rect 6472 35766 6500 37198
rect 6644 37120 6696 37126
rect 6644 37062 6696 37068
rect 6552 36780 6604 36786
rect 6552 36722 6604 36728
rect 6460 35760 6512 35766
rect 6460 35702 6512 35708
rect 6564 35290 6592 36722
rect 6656 36174 6684 37062
rect 6840 36854 6868 37334
rect 7012 37256 7064 37262
rect 7012 37198 7064 37204
rect 6828 36848 6880 36854
rect 6828 36790 6880 36796
rect 6828 36712 6880 36718
rect 6828 36654 6880 36660
rect 6644 36168 6696 36174
rect 6644 36110 6696 36116
rect 6552 35284 6604 35290
rect 6552 35226 6604 35232
rect 6368 34672 6420 34678
rect 6368 34614 6420 34620
rect 6368 34536 6420 34542
rect 6368 34478 6420 34484
rect 6380 34066 6408 34478
rect 6840 34202 6868 36654
rect 7024 36650 7052 37198
rect 7116 37126 7144 39374
rect 7286 39194 7342 40230
rect 7286 39142 7288 39194
rect 7340 39142 7342 39194
rect 7286 38106 7342 39142
rect 7286 38054 7288 38106
rect 7340 38054 7342 38106
rect 7104 37120 7156 37126
rect 7104 37062 7156 37068
rect 7286 37018 7342 38054
rect 7286 36966 7288 37018
rect 7340 36966 7342 37018
rect 7012 36644 7064 36650
rect 7012 36586 7064 36592
rect 7012 36032 7064 36038
rect 7012 35974 7064 35980
rect 7024 35698 7052 35974
rect 7286 35930 7342 36966
rect 7286 35878 7288 35930
rect 7340 35878 7342 35930
rect 7012 35692 7064 35698
rect 7012 35634 7064 35640
rect 6920 35624 6972 35630
rect 6920 35566 6972 35572
rect 6932 35086 6960 35566
rect 7012 35556 7064 35562
rect 7012 35498 7064 35504
rect 7024 35154 7052 35498
rect 7012 35148 7064 35154
rect 7012 35090 7064 35096
rect 6920 35080 6972 35086
rect 6920 35022 6972 35028
rect 6920 34944 6972 34950
rect 6920 34886 6972 34892
rect 6828 34196 6880 34202
rect 6828 34138 6880 34144
rect 6368 34060 6420 34066
rect 6368 34002 6420 34008
rect 6736 33516 6788 33522
rect 6736 33458 6788 33464
rect 6552 33380 6604 33386
rect 6552 33322 6604 33328
rect 6368 32836 6420 32842
rect 6368 32778 6420 32784
rect 6380 31890 6408 32778
rect 6564 32416 6592 33322
rect 6644 32428 6696 32434
rect 6564 32388 6644 32416
rect 6644 32370 6696 32376
rect 6552 32292 6604 32298
rect 6552 32234 6604 32240
rect 6368 31884 6420 31890
rect 6368 31826 6420 31832
rect 6564 31822 6592 32234
rect 6644 32224 6696 32230
rect 6644 32166 6696 32172
rect 6460 31816 6512 31822
rect 6460 31758 6512 31764
rect 6552 31816 6604 31822
rect 6552 31758 6604 31764
rect 6196 31726 6316 31754
rect 5172 31204 5224 31210
rect 5172 31146 5224 31152
rect 5184 29714 5212 31146
rect 5816 31136 5868 31142
rect 5816 31078 5868 31084
rect 5172 29708 5224 29714
rect 5172 29650 5224 29656
rect 4988 29640 5040 29646
rect 4988 29582 5040 29588
rect 4896 29232 4948 29238
rect 4896 29174 4948 29180
rect 4528 29164 4580 29170
rect 4528 29106 4580 29112
rect 4436 28960 4488 28966
rect 4436 28902 4488 28908
rect 4448 28626 4476 28902
rect 4540 28762 4568 29106
rect 5184 28966 5212 29650
rect 5356 29572 5408 29578
rect 5356 29514 5408 29520
rect 5172 28960 5224 28966
rect 5172 28902 5224 28908
rect 4528 28756 4580 28762
rect 4528 28698 4580 28704
rect 5368 28626 5396 29514
rect 4436 28620 4488 28626
rect 4436 28562 4488 28568
rect 5356 28620 5408 28626
rect 5356 28562 5408 28568
rect 4344 28552 4396 28558
rect 4344 28494 4396 28500
rect 4344 27940 4396 27946
rect 4344 27882 4396 27888
rect 4252 27872 4304 27878
rect 4252 27814 4304 27820
rect 2872 27532 2924 27538
rect 2872 27474 2924 27480
rect 3056 27532 3108 27538
rect 3896 27526 4016 27554
rect 4264 27538 4292 27814
rect 4356 27606 4384 27882
rect 4448 27674 4476 28562
rect 5540 28076 5592 28082
rect 5540 28018 5592 28024
rect 5448 28008 5500 28014
rect 5448 27950 5500 27956
rect 5356 27940 5408 27946
rect 5356 27882 5408 27888
rect 5172 27872 5224 27878
rect 5172 27814 5224 27820
rect 4436 27668 4488 27674
rect 4436 27610 4488 27616
rect 4344 27600 4396 27606
rect 4344 27542 4396 27548
rect 3056 27474 3108 27480
rect 2780 27464 2832 27470
rect 2780 27406 2832 27412
rect 2780 27328 2832 27334
rect 2780 27270 2832 27276
rect 2688 27056 2740 27062
rect 2688 26998 2740 27004
rect 2688 26784 2740 26790
rect 2688 26726 2740 26732
rect 2596 24880 2648 24886
rect 2596 24822 2648 24828
rect 2596 24744 2648 24750
rect 2596 24686 2648 24692
rect 2608 23322 2636 24686
rect 2700 24410 2728 26726
rect 2792 25974 2820 27270
rect 2884 26790 2912 27474
rect 2872 26784 2924 26790
rect 2872 26726 2924 26732
rect 3148 26784 3200 26790
rect 3148 26726 3200 26732
rect 2884 26382 2912 26726
rect 2872 26376 2924 26382
rect 2872 26318 2924 26324
rect 2780 25968 2832 25974
rect 2780 25910 2832 25916
rect 2884 25362 2912 26318
rect 2964 25424 3016 25430
rect 2964 25366 3016 25372
rect 2872 25356 2924 25362
rect 2872 25298 2924 25304
rect 2884 24698 2912 25298
rect 2976 24818 3004 25366
rect 2964 24812 3016 24818
rect 2964 24754 3016 24760
rect 2884 24670 3004 24698
rect 2688 24404 2740 24410
rect 2688 24346 2740 24352
rect 2780 24268 2832 24274
rect 2780 24210 2832 24216
rect 2688 24200 2740 24206
rect 2688 24142 2740 24148
rect 2700 23526 2728 24142
rect 2792 23866 2820 24210
rect 2780 23860 2832 23866
rect 2780 23802 2832 23808
rect 2976 23594 3004 24670
rect 2964 23588 3016 23594
rect 2964 23530 3016 23536
rect 2688 23520 2740 23526
rect 2688 23462 2740 23468
rect 2596 23316 2648 23322
rect 2596 23258 2648 23264
rect 2700 22794 2728 23462
rect 2976 23050 3004 23530
rect 3056 23112 3108 23118
rect 3056 23054 3108 23060
rect 2964 23044 3016 23050
rect 2964 22986 3016 22992
rect 2700 22766 3004 22794
rect 3068 22778 3096 23054
rect 2596 22568 2648 22574
rect 2596 22510 2648 22516
rect 2504 21548 2556 21554
rect 2504 21490 2556 21496
rect 2412 16448 2464 16454
rect 2412 16390 2464 16396
rect 2332 16238 2452 16266
rect 2228 16176 2280 16182
rect 2228 16118 2280 16124
rect 2134 15750 2136 15802
rect 2188 15750 2190 15802
rect 2134 14714 2190 15750
rect 2424 15502 2452 16238
rect 2516 15586 2544 21490
rect 2608 21146 2636 22510
rect 2700 22030 2728 22766
rect 2976 22658 3004 22766
rect 3056 22772 3108 22778
rect 3056 22714 3108 22720
rect 2976 22630 3096 22658
rect 3068 22574 3096 22630
rect 3056 22568 3108 22574
rect 3056 22510 3108 22516
rect 2688 22024 2740 22030
rect 2688 21966 2740 21972
rect 3160 21894 3188 26726
rect 3332 26512 3384 26518
rect 3332 26454 3384 26460
rect 3240 26376 3292 26382
rect 3240 26318 3292 26324
rect 3148 21888 3200 21894
rect 3148 21830 3200 21836
rect 2780 21480 2832 21486
rect 2780 21422 2832 21428
rect 2596 21140 2648 21146
rect 2596 21082 2648 21088
rect 2792 20942 2820 21422
rect 3056 21344 3108 21350
rect 3056 21286 3108 21292
rect 2872 21140 2924 21146
rect 2872 21082 2924 21088
rect 2780 20936 2832 20942
rect 2780 20878 2832 20884
rect 2688 20460 2740 20466
rect 2688 20402 2740 20408
rect 2596 20392 2648 20398
rect 2596 20334 2648 20340
rect 2608 19174 2636 20334
rect 2700 19378 2728 20402
rect 2792 19514 2820 20878
rect 2884 19854 2912 21082
rect 3068 20398 3096 21286
rect 3056 20392 3108 20398
rect 3056 20334 3108 20340
rect 2872 19848 2924 19854
rect 2872 19790 2924 19796
rect 2780 19508 2832 19514
rect 2780 19450 2832 19456
rect 2688 19372 2740 19378
rect 2884 19334 2912 19790
rect 3056 19780 3108 19786
rect 3056 19722 3108 19728
rect 2688 19314 2740 19320
rect 2792 19306 2912 19334
rect 2596 19168 2648 19174
rect 2596 19110 2648 19116
rect 2608 18698 2636 19110
rect 2596 18692 2648 18698
rect 2596 18634 2648 18640
rect 2608 16658 2636 18634
rect 2688 18216 2740 18222
rect 2688 18158 2740 18164
rect 2700 17746 2728 18158
rect 2688 17740 2740 17746
rect 2688 17682 2740 17688
rect 2688 17196 2740 17202
rect 2688 17138 2740 17144
rect 2596 16652 2648 16658
rect 2596 16594 2648 16600
rect 2596 16516 2648 16522
rect 2596 16458 2648 16464
rect 2608 15706 2636 16458
rect 2596 15700 2648 15706
rect 2596 15642 2648 15648
rect 2516 15558 2636 15586
rect 2412 15496 2464 15502
rect 2412 15438 2464 15444
rect 2320 15428 2372 15434
rect 2320 15370 2372 15376
rect 2228 15156 2280 15162
rect 2228 15098 2280 15104
rect 2134 14662 2136 14714
rect 2188 14662 2190 14714
rect 2134 13626 2190 14662
rect 2134 13574 2136 13626
rect 2188 13574 2190 13626
rect 2134 12538 2190 13574
rect 2240 12730 2268 15098
rect 2332 15094 2360 15370
rect 2412 15360 2464 15366
rect 2412 15302 2464 15308
rect 2504 15360 2556 15366
rect 2504 15302 2556 15308
rect 2320 15088 2372 15094
rect 2320 15030 2372 15036
rect 2332 13870 2360 15030
rect 2424 14550 2452 15302
rect 2516 15026 2544 15302
rect 2504 15020 2556 15026
rect 2504 14962 2556 14968
rect 2412 14544 2464 14550
rect 2412 14486 2464 14492
rect 2320 13864 2372 13870
rect 2320 13806 2372 13812
rect 2320 13456 2372 13462
rect 2320 13398 2372 13404
rect 2332 12850 2360 13398
rect 2516 13326 2544 14962
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 2320 12844 2372 12850
rect 2320 12786 2372 12792
rect 2412 12776 2464 12782
rect 2240 12702 2360 12730
rect 2412 12718 2464 12724
rect 2228 12640 2280 12646
rect 2228 12582 2280 12588
rect 2134 12486 2136 12538
rect 2188 12486 2190 12538
rect 2134 11450 2190 12486
rect 2240 12170 2268 12582
rect 2332 12170 2360 12702
rect 2228 12164 2280 12170
rect 2228 12106 2280 12112
rect 2320 12164 2372 12170
rect 2320 12106 2372 12112
rect 2134 11398 2136 11450
rect 2188 11398 2190 11450
rect 1860 11144 1912 11150
rect 1780 11104 1860 11132
rect 1780 10606 1808 11104
rect 1860 11086 1912 11092
rect 1860 10736 1912 10742
rect 1860 10678 1912 10684
rect 1768 10600 1820 10606
rect 1768 10542 1820 10548
rect 1768 10464 1820 10470
rect 1768 10406 1820 10412
rect 1780 9994 1808 10406
rect 1768 9988 1820 9994
rect 1768 9930 1820 9936
rect 1768 9648 1820 9654
rect 1768 9590 1820 9596
rect 1676 8968 1728 8974
rect 1676 8910 1728 8916
rect 1780 8498 1808 9590
rect 1768 8492 1820 8498
rect 1768 8434 1820 8440
rect 1768 7880 1820 7886
rect 1872 7868 1900 10678
rect 1964 9382 1992 11206
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 1952 9376 2004 9382
rect 1952 9318 2004 9324
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 1964 8566 1992 8774
rect 1952 8560 2004 8566
rect 1952 8502 2004 8508
rect 1820 7840 1900 7868
rect 1768 7822 1820 7828
rect 1780 7410 1808 7822
rect 1952 7744 2004 7750
rect 1952 7686 2004 7692
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 1768 6724 1820 6730
rect 1768 6666 1820 6672
rect 1780 6458 1808 6666
rect 1768 6452 1820 6458
rect 1768 6394 1820 6400
rect 1964 6322 1992 7686
rect 2056 7546 2084 10610
rect 2134 10362 2190 11398
rect 2424 11354 2452 12718
rect 2516 11898 2544 13262
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2228 11008 2280 11014
rect 2228 10950 2280 10956
rect 2240 10674 2268 10950
rect 2228 10668 2280 10674
rect 2228 10610 2280 10616
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2134 10310 2136 10362
rect 2188 10310 2190 10362
rect 2134 9274 2190 10310
rect 2228 9920 2280 9926
rect 2228 9862 2280 9868
rect 2240 9586 2268 9862
rect 2332 9654 2360 10610
rect 2320 9648 2372 9654
rect 2320 9590 2372 9596
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2134 9222 2136 9274
rect 2188 9222 2190 9274
rect 2134 8186 2190 9222
rect 2240 9042 2268 9522
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 2228 9036 2280 9042
rect 2228 8978 2280 8984
rect 2332 8430 2360 9454
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2134 8134 2136 8186
rect 2188 8134 2190 8186
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 2134 7098 2190 8134
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2240 7410 2268 7822
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2240 7206 2268 7346
rect 2332 7342 2360 8366
rect 2424 8362 2452 9454
rect 2608 9110 2636 15558
rect 2700 14618 2728 17138
rect 2792 16590 2820 19306
rect 2964 19168 3016 19174
rect 2964 19110 3016 19116
rect 2872 18692 2924 18698
rect 2872 18634 2924 18640
rect 2884 17678 2912 18634
rect 2976 18290 3004 19110
rect 2964 18284 3016 18290
rect 2964 18226 3016 18232
rect 3068 17882 3096 19722
rect 3148 18284 3200 18290
rect 3148 18226 3200 18232
rect 3160 18154 3188 18226
rect 3148 18148 3200 18154
rect 3148 18090 3200 18096
rect 3160 17882 3188 18090
rect 3056 17876 3108 17882
rect 3056 17818 3108 17824
rect 3148 17876 3200 17882
rect 3148 17818 3200 17824
rect 3056 17740 3108 17746
rect 3056 17682 3108 17688
rect 2872 17672 2924 17678
rect 2872 17614 2924 17620
rect 2872 17536 2924 17542
rect 2872 17478 2924 17484
rect 2780 16584 2832 16590
rect 2780 16526 2832 16532
rect 2884 15638 2912 17478
rect 2872 15632 2924 15638
rect 2872 15574 2924 15580
rect 2884 15162 2912 15574
rect 3068 15450 3096 17682
rect 3148 16448 3200 16454
rect 3148 16390 3200 16396
rect 3160 16182 3188 16390
rect 3148 16176 3200 16182
rect 3148 16118 3200 16124
rect 3068 15422 3188 15450
rect 3056 15360 3108 15366
rect 3056 15302 3108 15308
rect 2872 15156 2924 15162
rect 2872 15098 2924 15104
rect 2688 14612 2740 14618
rect 2688 14554 2740 14560
rect 2688 14340 2740 14346
rect 2688 14282 2740 14288
rect 2700 13530 2728 14282
rect 2780 14272 2832 14278
rect 2780 14214 2832 14220
rect 2792 13870 2820 14214
rect 3068 14006 3096 15302
rect 3160 14006 3188 15422
rect 3056 14000 3108 14006
rect 3056 13942 3108 13948
rect 3148 14000 3200 14006
rect 3148 13942 3200 13948
rect 2780 13864 2832 13870
rect 3160 13852 3188 13942
rect 2780 13806 2832 13812
rect 2976 13824 3188 13852
rect 2688 13524 2740 13530
rect 2688 13466 2740 13472
rect 2792 12850 2820 13806
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 2780 12844 2832 12850
rect 2780 12786 2832 12792
rect 2884 12186 2912 12854
rect 2976 12442 3004 13824
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 3148 13524 3200 13530
rect 3148 13466 3200 13472
rect 2964 12436 3016 12442
rect 2964 12378 3016 12384
rect 2792 12158 2912 12186
rect 2688 11688 2740 11694
rect 2688 11630 2740 11636
rect 2700 10062 2728 11630
rect 2792 11150 2820 12158
rect 2976 11150 3004 12378
rect 3068 12306 3096 13466
rect 3056 12300 3108 12306
rect 3056 12242 3108 12248
rect 3068 11558 3096 12242
rect 3056 11552 3108 11558
rect 3056 11494 3108 11500
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 3068 11098 3096 11494
rect 3160 11218 3188 13466
rect 3148 11212 3200 11218
rect 3148 11154 3200 11160
rect 2792 10690 2820 11086
rect 2872 11076 2924 11082
rect 3068 11070 3188 11098
rect 2872 11018 2924 11024
rect 2884 10810 2912 11018
rect 2872 10804 2924 10810
rect 2872 10746 2924 10752
rect 2792 10662 2912 10690
rect 2780 10532 2832 10538
rect 2780 10474 2832 10480
rect 2688 10056 2740 10062
rect 2688 9998 2740 10004
rect 2792 9602 2820 10474
rect 2700 9586 2820 9602
rect 2688 9580 2820 9586
rect 2740 9574 2820 9580
rect 2688 9522 2740 9528
rect 2596 9104 2648 9110
rect 2596 9046 2648 9052
rect 2412 8356 2464 8362
rect 2412 8298 2464 8304
rect 2596 8288 2648 8294
rect 2596 8230 2648 8236
rect 2688 8288 2740 8294
rect 2688 8230 2740 8236
rect 2412 7948 2464 7954
rect 2412 7890 2464 7896
rect 2320 7336 2372 7342
rect 2320 7278 2372 7284
rect 2228 7200 2280 7206
rect 2228 7142 2280 7148
rect 2134 7046 2136 7098
rect 2188 7046 2190 7098
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 1584 4820 1636 4826
rect 1584 4762 1636 4768
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 1412 2514 1440 4626
rect 1688 4622 1716 4966
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1780 2774 1808 6258
rect 2134 6010 2190 7046
rect 2134 5958 2136 6010
rect 2188 5958 2190 6010
rect 2044 5228 2096 5234
rect 2044 5170 2096 5176
rect 2056 4282 2084 5170
rect 2134 4922 2190 5958
rect 2134 4870 2136 4922
rect 2188 4870 2190 4922
rect 2044 4276 2096 4282
rect 2044 4218 2096 4224
rect 2134 3834 2190 4870
rect 2240 4146 2268 7142
rect 2424 6934 2452 7890
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2516 7410 2544 7822
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2412 6928 2464 6934
rect 2412 6870 2464 6876
rect 2320 6724 2372 6730
rect 2320 6666 2372 6672
rect 2332 6254 2360 6666
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 2320 6248 2372 6254
rect 2320 6190 2372 6196
rect 2332 5302 2360 6190
rect 2424 5846 2452 6394
rect 2504 6384 2556 6390
rect 2504 6326 2556 6332
rect 2412 5840 2464 5846
rect 2412 5782 2464 5788
rect 2320 5296 2372 5302
rect 2320 5238 2372 5244
rect 2424 4146 2452 5782
rect 2228 4140 2280 4146
rect 2412 4140 2464 4146
rect 2228 4082 2280 4088
rect 2332 4100 2412 4128
rect 2134 3782 2136 3834
rect 2188 3782 2190 3834
rect 1780 2746 1900 2774
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1872 1562 1900 2746
rect 2134 2746 2190 3782
rect 2240 3126 2268 4082
rect 2228 3120 2280 3126
rect 2228 3062 2280 3068
rect 2332 3058 2360 4100
rect 2412 4082 2464 4088
rect 2412 4004 2464 4010
rect 2412 3946 2464 3952
rect 2424 3534 2452 3946
rect 2412 3528 2464 3534
rect 2412 3470 2464 3476
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 2320 2848 2372 2854
rect 2320 2790 2372 2796
rect 2134 2694 2136 2746
rect 2188 2694 2190 2746
rect 2044 2372 2096 2378
rect 2044 2314 2096 2320
rect 2056 2106 2084 2314
rect 2044 2100 2096 2106
rect 2044 2042 2096 2048
rect 2134 1658 2190 2694
rect 2332 1970 2360 2790
rect 2320 1964 2372 1970
rect 2320 1906 2372 1912
rect 2134 1606 2136 1658
rect 2188 1606 2190 1658
rect 1860 1556 1912 1562
rect 1860 1498 1912 1504
rect 2134 1040 2190 1606
rect 2516 1358 2544 6326
rect 2608 6254 2636 8230
rect 2700 8090 2728 8230
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 2700 6322 2728 7346
rect 2884 6458 2912 10662
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 3068 10266 3096 10542
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 3068 9674 3096 10202
rect 2976 9646 3096 9674
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 2688 5636 2740 5642
rect 2688 5578 2740 5584
rect 2700 5370 2728 5578
rect 2688 5364 2740 5370
rect 2688 5306 2740 5312
rect 2596 5160 2648 5166
rect 2596 5102 2648 5108
rect 2608 4690 2636 5102
rect 2596 4684 2648 4690
rect 2596 4626 2648 4632
rect 2608 3058 2636 4626
rect 2688 4616 2740 4622
rect 2688 4558 2740 4564
rect 2700 4146 2728 4558
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2688 3596 2740 3602
rect 2688 3538 2740 3544
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 2608 2650 2636 2994
rect 2596 2644 2648 2650
rect 2596 2586 2648 2592
rect 2700 1902 2728 3538
rect 2780 3188 2832 3194
rect 2780 3130 2832 3136
rect 2688 1896 2740 1902
rect 2688 1838 2740 1844
rect 2504 1352 2556 1358
rect 2504 1294 2556 1300
rect 2792 800 2820 3130
rect 2884 1562 2912 4082
rect 2872 1556 2924 1562
rect 2872 1498 2924 1504
rect 2976 1494 3004 9646
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 3068 7954 3096 8774
rect 3056 7948 3108 7954
rect 3056 7890 3108 7896
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 3068 5234 3096 6598
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 3160 5114 3188 11070
rect 3252 9058 3280 26318
rect 3344 9178 3372 26454
rect 3792 26240 3844 26246
rect 3792 26182 3844 26188
rect 3804 25242 3832 26182
rect 3988 25498 4016 27526
rect 4252 27532 4304 27538
rect 4252 27474 4304 27480
rect 5184 27470 5212 27814
rect 4160 27464 4212 27470
rect 4160 27406 4212 27412
rect 5172 27464 5224 27470
rect 5172 27406 5224 27412
rect 4068 27328 4120 27334
rect 4068 27270 4120 27276
rect 4080 26994 4108 27270
rect 4068 26988 4120 26994
rect 4068 26930 4120 26936
rect 4172 26586 4200 27406
rect 4344 27396 4396 27402
rect 4344 27338 4396 27344
rect 5080 27396 5132 27402
rect 5080 27338 5132 27344
rect 4160 26580 4212 26586
rect 4160 26522 4212 26528
rect 4068 26376 4120 26382
rect 4068 26318 4120 26324
rect 3976 25492 4028 25498
rect 3976 25434 4028 25440
rect 4080 25378 4108 26318
rect 4356 25974 4384 27338
rect 4528 26444 4580 26450
rect 4528 26386 4580 26392
rect 4344 25968 4396 25974
rect 4344 25910 4396 25916
rect 4436 25696 4488 25702
rect 4436 25638 4488 25644
rect 3988 25350 4108 25378
rect 3804 25214 3924 25242
rect 3988 25226 4016 25350
rect 3792 25152 3844 25158
rect 3792 25094 3844 25100
rect 3516 24744 3568 24750
rect 3516 24686 3568 24692
rect 3424 22636 3476 22642
rect 3424 22578 3476 22584
rect 3436 9926 3464 22578
rect 3528 21146 3556 24686
rect 3804 24410 3832 25094
rect 3792 24404 3844 24410
rect 3792 24346 3844 24352
rect 3700 23792 3752 23798
rect 3700 23734 3752 23740
rect 3608 22432 3660 22438
rect 3608 22374 3660 22380
rect 3620 21622 3648 22374
rect 3608 21616 3660 21622
rect 3608 21558 3660 21564
rect 3516 21140 3568 21146
rect 3516 21082 3568 21088
rect 3516 19916 3568 19922
rect 3516 19858 3568 19864
rect 3528 19378 3556 19858
rect 3608 19712 3660 19718
rect 3608 19654 3660 19660
rect 3516 19372 3568 19378
rect 3516 19314 3568 19320
rect 3620 17678 3648 19654
rect 3608 17672 3660 17678
rect 3608 17614 3660 17620
rect 3516 17536 3568 17542
rect 3516 17478 3568 17484
rect 3528 17270 3556 17478
rect 3516 17264 3568 17270
rect 3516 17206 3568 17212
rect 3620 15026 3648 17614
rect 3608 15020 3660 15026
rect 3608 14962 3660 14968
rect 3516 14816 3568 14822
rect 3516 14758 3568 14764
rect 3528 14618 3556 14758
rect 3516 14612 3568 14618
rect 3516 14554 3568 14560
rect 3516 14272 3568 14278
rect 3516 14214 3568 14220
rect 3528 14006 3556 14214
rect 3516 14000 3568 14006
rect 3516 13942 3568 13948
rect 3620 13462 3648 14962
rect 3608 13456 3660 13462
rect 3608 13398 3660 13404
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 3528 12986 3556 13126
rect 3516 12980 3568 12986
rect 3516 12922 3568 12928
rect 3608 12640 3660 12646
rect 3608 12582 3660 12588
rect 3620 12306 3648 12582
rect 3608 12300 3660 12306
rect 3608 12242 3660 12248
rect 3712 12186 3740 23734
rect 3792 23520 3844 23526
rect 3792 23462 3844 23468
rect 3804 23186 3832 23462
rect 3792 23180 3844 23186
rect 3792 23122 3844 23128
rect 3792 22636 3844 22642
rect 3792 22578 3844 22584
rect 3804 22234 3832 22578
rect 3896 22234 3924 25214
rect 3976 25220 4028 25226
rect 3976 25162 4028 25168
rect 3988 23254 4016 25162
rect 4448 24886 4476 25638
rect 4436 24880 4488 24886
rect 4436 24822 4488 24828
rect 4068 23792 4120 23798
rect 4068 23734 4120 23740
rect 3976 23248 4028 23254
rect 3976 23190 4028 23196
rect 4080 22642 4108 23734
rect 4160 23520 4212 23526
rect 4160 23462 4212 23468
rect 4172 23118 4200 23462
rect 4448 23186 4476 24822
rect 4540 24274 4568 26386
rect 4712 26376 4764 26382
rect 4712 26318 4764 26324
rect 4988 26376 5040 26382
rect 4988 26318 5040 26324
rect 4724 25294 4752 26318
rect 4804 26308 4856 26314
rect 4804 26250 4856 26256
rect 4816 25906 4844 26250
rect 4804 25900 4856 25906
rect 4804 25842 4856 25848
rect 4712 25288 4764 25294
rect 4712 25230 4764 25236
rect 4528 24268 4580 24274
rect 4528 24210 4580 24216
rect 4528 24064 4580 24070
rect 4528 24006 4580 24012
rect 4436 23180 4488 23186
rect 4436 23122 4488 23128
rect 4160 23112 4212 23118
rect 4160 23054 4212 23060
rect 4160 22976 4212 22982
rect 4160 22918 4212 22924
rect 4068 22636 4120 22642
rect 4068 22578 4120 22584
rect 3792 22228 3844 22234
rect 3792 22170 3844 22176
rect 3884 22228 3936 22234
rect 3884 22170 3936 22176
rect 3792 22024 3844 22030
rect 3792 21966 3844 21972
rect 3804 21622 3832 21966
rect 3792 21616 3844 21622
rect 3792 21558 3844 21564
rect 3884 19848 3936 19854
rect 3884 19790 3936 19796
rect 3896 19514 3924 19790
rect 3884 19508 3936 19514
rect 3884 19450 3936 19456
rect 3792 19372 3844 19378
rect 3792 19314 3844 19320
rect 3804 18358 3832 19314
rect 3792 18352 3844 18358
rect 3792 18294 3844 18300
rect 3804 16658 3832 18294
rect 3896 18222 3924 19450
rect 3976 19304 4028 19310
rect 3976 19246 4028 19252
rect 3988 18834 4016 19246
rect 3976 18828 4028 18834
rect 3976 18770 4028 18776
rect 3884 18216 3936 18222
rect 3884 18158 3936 18164
rect 3896 17338 3924 18158
rect 3988 17660 4016 18770
rect 4080 17882 4108 22578
rect 4172 18358 4200 22918
rect 4252 22568 4304 22574
rect 4252 22510 4304 22516
rect 4264 21894 4292 22510
rect 4436 22024 4488 22030
rect 4436 21966 4488 21972
rect 4252 21888 4304 21894
rect 4252 21830 4304 21836
rect 4448 21486 4476 21966
rect 4436 21480 4488 21486
rect 4436 21422 4488 21428
rect 4252 20392 4304 20398
rect 4252 20334 4304 20340
rect 4160 18352 4212 18358
rect 4160 18294 4212 18300
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 4068 17672 4120 17678
rect 3988 17632 4068 17660
rect 3884 17332 3936 17338
rect 3884 17274 3936 17280
rect 3896 17066 3924 17274
rect 3884 17060 3936 17066
rect 3884 17002 3936 17008
rect 3792 16652 3844 16658
rect 3792 16594 3844 16600
rect 3804 16096 3832 16594
rect 3884 16108 3936 16114
rect 3804 16068 3884 16096
rect 3804 15570 3832 16068
rect 3884 16050 3936 16056
rect 3792 15564 3844 15570
rect 3792 15506 3844 15512
rect 3988 15162 4016 17632
rect 4068 17614 4120 17620
rect 4264 16776 4292 20334
rect 4344 19712 4396 19718
rect 4344 19654 4396 19660
rect 4356 19514 4384 19654
rect 4344 19508 4396 19514
rect 4344 19450 4396 19456
rect 4436 19304 4488 19310
rect 4436 19246 4488 19252
rect 4448 17678 4476 19246
rect 4436 17672 4488 17678
rect 4436 17614 4488 17620
rect 4172 16748 4292 16776
rect 3884 15156 3936 15162
rect 3884 15098 3936 15104
rect 3976 15156 4028 15162
rect 3976 15098 4028 15104
rect 3792 13320 3844 13326
rect 3792 13262 3844 13268
rect 3528 12158 3740 12186
rect 3804 12170 3832 13262
rect 3896 12442 3924 15098
rect 3976 15020 4028 15026
rect 3976 14962 4028 14968
rect 3988 13938 4016 14962
rect 4068 14544 4120 14550
rect 4172 14532 4200 16748
rect 4252 16584 4304 16590
rect 4252 16526 4304 16532
rect 4120 14504 4200 14532
rect 4068 14486 4120 14492
rect 3976 13932 4028 13938
rect 3976 13874 4028 13880
rect 3988 13394 4016 13874
rect 3976 13388 4028 13394
rect 3976 13330 4028 13336
rect 3976 13252 4028 13258
rect 3976 13194 4028 13200
rect 3988 12782 4016 13194
rect 4080 12918 4108 14486
rect 4160 14408 4212 14414
rect 4264 14396 4292 16526
rect 4436 16108 4488 16114
rect 4436 16050 4488 16056
rect 4344 15972 4396 15978
rect 4344 15914 4396 15920
rect 4356 15570 4384 15914
rect 4344 15564 4396 15570
rect 4344 15506 4396 15512
rect 4448 15042 4476 16050
rect 4212 14368 4292 14396
rect 4356 15014 4476 15042
rect 4160 14350 4212 14356
rect 4068 12912 4120 12918
rect 4068 12854 4120 12860
rect 3976 12776 4028 12782
rect 3976 12718 4028 12724
rect 3884 12436 3936 12442
rect 3884 12378 3936 12384
rect 3792 12164 3844 12170
rect 3424 9920 3476 9926
rect 3424 9862 3476 9868
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3252 9030 3464 9058
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3252 8430 3280 8910
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3240 8424 3292 8430
rect 3240 8366 3292 8372
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 3068 5086 3188 5114
rect 3068 1902 3096 5086
rect 3252 4486 3280 5510
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3344 4298 3372 8434
rect 3252 4270 3372 4298
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 3160 3670 3188 3878
rect 3148 3664 3200 3670
rect 3148 3606 3200 3612
rect 3148 2372 3200 2378
rect 3148 2314 3200 2320
rect 3160 2106 3188 2314
rect 3148 2100 3200 2106
rect 3148 2042 3200 2048
rect 3056 1896 3108 1902
rect 3056 1838 3108 1844
rect 2964 1488 3016 1494
rect 2964 1430 3016 1436
rect 3252 1222 3280 4270
rect 3332 2848 3384 2854
rect 3332 2790 3384 2796
rect 3344 1970 3372 2790
rect 3436 2774 3464 9030
rect 3528 4010 3556 12158
rect 3792 12106 3844 12112
rect 3700 12096 3752 12102
rect 3700 12038 3752 12044
rect 3712 11830 3740 12038
rect 3700 11824 3752 11830
rect 3700 11766 3752 11772
rect 4172 11354 4200 14350
rect 4356 14278 4384 15014
rect 4436 14952 4488 14958
rect 4436 14894 4488 14900
rect 4344 14272 4396 14278
rect 4344 14214 4396 14220
rect 4252 14000 4304 14006
rect 4252 13942 4304 13948
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 3620 10538 3648 11290
rect 4264 11234 4292 13942
rect 4344 13728 4396 13734
rect 4344 13670 4396 13676
rect 4356 12850 4384 13670
rect 4344 12844 4396 12850
rect 4344 12786 4396 12792
rect 4448 12238 4476 14894
rect 4436 12232 4488 12238
rect 4436 12174 4488 12180
rect 4540 11880 4568 24006
rect 4724 23594 4752 25230
rect 4712 23588 4764 23594
rect 4712 23530 4764 23536
rect 4620 22636 4672 22642
rect 4620 22578 4672 22584
rect 4632 20448 4660 22578
rect 4724 22030 4752 23530
rect 4816 23526 4844 25842
rect 5000 25294 5028 26318
rect 5092 26246 5120 27338
rect 5080 26240 5132 26246
rect 5080 26182 5132 26188
rect 5092 25294 5120 26182
rect 4988 25288 5040 25294
rect 4988 25230 5040 25236
rect 5080 25288 5132 25294
rect 5080 25230 5132 25236
rect 4896 24812 4948 24818
rect 4896 24754 4948 24760
rect 4908 24410 4936 24754
rect 4896 24404 4948 24410
rect 4896 24346 4948 24352
rect 5000 23662 5028 25230
rect 5092 24954 5120 25230
rect 5172 25152 5224 25158
rect 5172 25094 5224 25100
rect 5080 24948 5132 24954
rect 5080 24890 5132 24896
rect 5092 24070 5120 24890
rect 5184 24206 5212 25094
rect 5368 24410 5396 27882
rect 5356 24404 5408 24410
rect 5356 24346 5408 24352
rect 5172 24200 5224 24206
rect 5172 24142 5224 24148
rect 5080 24064 5132 24070
rect 5080 24006 5132 24012
rect 4988 23656 5040 23662
rect 4988 23598 5040 23604
rect 5264 23656 5316 23662
rect 5264 23598 5316 23604
rect 4804 23520 4856 23526
rect 4804 23462 4856 23468
rect 5172 23520 5224 23526
rect 5172 23462 5224 23468
rect 4804 23316 4856 23322
rect 4804 23258 4856 23264
rect 4816 22710 4844 23258
rect 4804 22704 4856 22710
rect 4804 22646 4856 22652
rect 4988 22500 5040 22506
rect 4988 22442 5040 22448
rect 4896 22160 4948 22166
rect 4896 22102 4948 22108
rect 4712 22024 4764 22030
rect 4712 21966 4764 21972
rect 4908 21554 4936 22102
rect 4896 21548 4948 21554
rect 4896 21490 4948 21496
rect 5000 21350 5028 22442
rect 5184 22098 5212 23462
rect 5276 23186 5304 23598
rect 5368 23322 5396 24346
rect 5460 23594 5488 27950
rect 5552 26586 5580 28018
rect 5724 28008 5776 28014
rect 5724 27950 5776 27956
rect 5736 26858 5764 27950
rect 5724 26852 5776 26858
rect 5724 26794 5776 26800
rect 5632 26784 5684 26790
rect 5632 26726 5684 26732
rect 5540 26580 5592 26586
rect 5540 26522 5592 26528
rect 5540 24404 5592 24410
rect 5540 24346 5592 24352
rect 5552 23866 5580 24346
rect 5540 23860 5592 23866
rect 5540 23802 5592 23808
rect 5448 23588 5500 23594
rect 5448 23530 5500 23536
rect 5356 23316 5408 23322
rect 5356 23258 5408 23264
rect 5264 23180 5316 23186
rect 5264 23122 5316 23128
rect 5276 22166 5304 23122
rect 5356 23112 5408 23118
rect 5356 23054 5408 23060
rect 5264 22160 5316 22166
rect 5264 22102 5316 22108
rect 5172 22092 5224 22098
rect 5172 22034 5224 22040
rect 5080 22024 5132 22030
rect 5080 21966 5132 21972
rect 5092 21690 5120 21966
rect 5080 21684 5132 21690
rect 5080 21626 5132 21632
rect 5264 21480 5316 21486
rect 5264 21422 5316 21428
rect 4712 21344 4764 21350
rect 4712 21286 4764 21292
rect 4988 21344 5040 21350
rect 4988 21286 5040 21292
rect 4724 20874 4752 21286
rect 4712 20868 4764 20874
rect 4712 20810 4764 20816
rect 5000 20534 5028 21286
rect 5080 20868 5132 20874
rect 5080 20810 5132 20816
rect 5092 20602 5120 20810
rect 5080 20596 5132 20602
rect 5080 20538 5132 20544
rect 4988 20528 5040 20534
rect 4988 20470 5040 20476
rect 4712 20460 4764 20466
rect 4632 20420 4712 20448
rect 4712 20402 4764 20408
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 4632 17814 4660 19110
rect 4724 18766 4752 20402
rect 5172 20324 5224 20330
rect 5172 20266 5224 20272
rect 5184 20058 5212 20266
rect 5172 20052 5224 20058
rect 5172 19994 5224 20000
rect 5184 19378 5212 19994
rect 5172 19372 5224 19378
rect 5172 19314 5224 19320
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4896 18760 4948 18766
rect 4896 18702 4948 18708
rect 4620 17808 4672 17814
rect 4620 17750 4672 17756
rect 4632 15416 4660 17750
rect 4724 15484 4752 18702
rect 4908 18222 4936 18702
rect 5172 18692 5224 18698
rect 5172 18634 5224 18640
rect 4896 18216 4948 18222
rect 4896 18158 4948 18164
rect 5080 18080 5132 18086
rect 5080 18022 5132 18028
rect 4988 17876 5040 17882
rect 4988 17818 5040 17824
rect 5000 17270 5028 17818
rect 5092 17610 5120 18022
rect 5080 17604 5132 17610
rect 5080 17546 5132 17552
rect 4988 17264 5040 17270
rect 4988 17206 5040 17212
rect 4804 16448 4856 16454
rect 4804 16390 4856 16396
rect 4816 15706 4844 16390
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 5000 15620 5028 17206
rect 5092 15978 5120 17546
rect 5184 17066 5212 18634
rect 5172 17060 5224 17066
rect 5172 17002 5224 17008
rect 5080 15972 5132 15978
rect 5080 15914 5132 15920
rect 5080 15632 5132 15638
rect 5000 15592 5080 15620
rect 5080 15574 5132 15580
rect 4724 15456 4936 15484
rect 4908 15450 4936 15456
rect 4908 15422 5028 15450
rect 4632 15388 4844 15416
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 4632 13870 4660 14418
rect 4620 13864 4672 13870
rect 4620 13806 4672 13812
rect 3988 11206 4292 11234
rect 4448 11852 4568 11880
rect 3608 10532 3660 10538
rect 3608 10474 3660 10480
rect 3884 10260 3936 10266
rect 3884 10202 3936 10208
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3700 9716 3752 9722
rect 3700 9658 3752 9664
rect 3608 9444 3660 9450
rect 3608 9386 3660 9392
rect 3620 8566 3648 9386
rect 3608 8560 3660 8566
rect 3608 8502 3660 8508
rect 3608 7812 3660 7818
rect 3608 7754 3660 7760
rect 3620 7410 3648 7754
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3620 5846 3648 6938
rect 3608 5840 3660 5846
rect 3608 5782 3660 5788
rect 3712 4434 3740 9658
rect 3804 5930 3832 9862
rect 3896 9722 3924 10202
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3988 9450 4016 11206
rect 4448 11150 4476 11852
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4436 11144 4488 11150
rect 4436 11086 4488 11092
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 3976 9444 4028 9450
rect 3976 9386 4028 9392
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 3896 6662 3924 9114
rect 3988 8498 4016 9386
rect 4068 8900 4120 8906
rect 4068 8842 4120 8848
rect 3976 8492 4028 8498
rect 3976 8434 4028 8440
rect 3976 8356 4028 8362
rect 3976 8298 4028 8304
rect 3988 7546 4016 8298
rect 3976 7540 4028 7546
rect 3976 7482 4028 7488
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 3988 6798 4016 7142
rect 4080 7002 4108 8842
rect 4172 8498 4200 9998
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 4172 6458 4200 8434
rect 4264 6662 4292 11086
rect 4540 10742 4568 11698
rect 4632 11694 4660 13806
rect 4712 13456 4764 13462
rect 4816 13444 4844 15388
rect 4896 15156 4948 15162
rect 4896 15098 4948 15104
rect 4764 13416 4844 13444
rect 4712 13398 4764 13404
rect 4724 12102 4752 13398
rect 4804 13184 4856 13190
rect 4804 13126 4856 13132
rect 4816 12986 4844 13126
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4908 12288 4936 15098
rect 5000 13326 5028 15422
rect 5080 15020 5132 15026
rect 5080 14962 5132 14968
rect 4988 13320 5040 13326
rect 4988 13262 5040 13268
rect 4816 12260 4936 12288
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4528 10736 4580 10742
rect 4816 10690 4844 12260
rect 4896 12164 4948 12170
rect 4896 12106 4948 12112
rect 4528 10678 4580 10684
rect 4632 10662 4844 10690
rect 4528 10600 4580 10606
rect 4528 10542 4580 10548
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 4356 8634 4384 8774
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 3804 5902 4016 5930
rect 3884 5840 3936 5846
rect 3884 5782 3936 5788
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3804 4554 3832 5510
rect 3896 5098 3924 5782
rect 3884 5092 3936 5098
rect 3884 5034 3936 5040
rect 3792 4548 3844 4554
rect 3792 4490 3844 4496
rect 3712 4406 3924 4434
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 3516 4004 3568 4010
rect 3516 3946 3568 3952
rect 3528 2922 3556 3946
rect 3712 3602 3740 4014
rect 3700 3596 3752 3602
rect 3700 3538 3752 3544
rect 3516 2916 3568 2922
rect 3516 2858 3568 2864
rect 3804 2854 3832 4082
rect 3792 2848 3844 2854
rect 3792 2790 3844 2796
rect 3436 2746 3556 2774
rect 3528 2310 3556 2746
rect 3516 2304 3568 2310
rect 3516 2246 3568 2252
rect 3332 1964 3384 1970
rect 3332 1906 3384 1912
rect 3896 1358 3924 4406
rect 3988 4214 4016 5902
rect 4172 5302 4200 6394
rect 4264 5930 4292 6598
rect 4356 6118 4384 6802
rect 4448 6322 4476 10406
rect 4540 9586 4568 10542
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 4540 7410 4568 9522
rect 4528 7404 4580 7410
rect 4528 7346 4580 7352
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4264 5902 4476 5930
rect 4344 5772 4396 5778
rect 4344 5714 4396 5720
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 4160 5296 4212 5302
rect 4160 5238 4212 5244
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 3976 4208 4028 4214
rect 3976 4150 4028 4156
rect 3988 2990 4016 4150
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 4080 1970 4108 4966
rect 4172 3058 4200 5238
rect 4264 4146 4292 5646
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 4356 3534 4384 5714
rect 4448 5574 4476 5902
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4540 5030 4568 7346
rect 4632 6934 4660 10662
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4712 9648 4764 9654
rect 4712 9590 4764 9596
rect 4620 6928 4672 6934
rect 4620 6870 4672 6876
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4632 6458 4660 6734
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4724 6118 4752 9590
rect 4816 8956 4844 10542
rect 4908 9654 4936 12106
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 5000 10674 5028 11698
rect 5092 11354 5120 14962
rect 5184 14498 5212 17002
rect 5276 16658 5304 21422
rect 5368 20618 5396 23054
rect 5448 22976 5500 22982
rect 5448 22918 5500 22924
rect 5460 22642 5488 22918
rect 5448 22636 5500 22642
rect 5448 22578 5500 22584
rect 5368 20590 5488 20618
rect 5356 20460 5408 20466
rect 5356 20402 5408 20408
rect 5368 20262 5396 20402
rect 5356 20256 5408 20262
rect 5356 20198 5408 20204
rect 5264 16652 5316 16658
rect 5264 16594 5316 16600
rect 5184 14470 5304 14498
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 5184 12646 5212 14350
rect 5276 13938 5304 14470
rect 5368 14414 5396 20198
rect 5460 18970 5488 20590
rect 5448 18964 5500 18970
rect 5448 18906 5500 18912
rect 5448 18624 5500 18630
rect 5448 18566 5500 18572
rect 5460 18358 5488 18566
rect 5448 18352 5500 18358
rect 5448 18294 5500 18300
rect 5552 17882 5580 23802
rect 5644 21078 5672 26726
rect 5736 26586 5764 26794
rect 5724 26580 5776 26586
rect 5724 26522 5776 26528
rect 5828 26466 5856 31078
rect 5908 30728 5960 30734
rect 5908 30670 5960 30676
rect 5736 26438 5856 26466
rect 5736 23866 5764 26438
rect 5816 26376 5868 26382
rect 5816 26318 5868 26324
rect 5724 23860 5776 23866
rect 5724 23802 5776 23808
rect 5724 23724 5776 23730
rect 5724 23666 5776 23672
rect 5736 22234 5764 23666
rect 5828 23118 5856 26318
rect 5920 23168 5948 30670
rect 6092 30592 6144 30598
rect 6092 30534 6144 30540
rect 6000 29776 6052 29782
rect 6000 29718 6052 29724
rect 6012 25770 6040 29718
rect 6000 25764 6052 25770
rect 6000 25706 6052 25712
rect 6012 23236 6040 25706
rect 6104 24138 6132 30534
rect 6184 29708 6236 29714
rect 6184 29650 6236 29656
rect 6196 29510 6224 29650
rect 6184 29504 6236 29510
rect 6184 29446 6236 29452
rect 6196 28490 6224 29446
rect 6184 28484 6236 28490
rect 6184 28426 6236 28432
rect 6092 24132 6144 24138
rect 6092 24074 6144 24080
rect 6196 23730 6224 28426
rect 6288 25922 6316 31726
rect 6472 30938 6500 31758
rect 6656 31414 6684 32166
rect 6644 31408 6696 31414
rect 6644 31350 6696 31356
rect 6460 30932 6512 30938
rect 6460 30874 6512 30880
rect 6748 30682 6776 33458
rect 6840 32910 6868 34138
rect 6828 32904 6880 32910
rect 6828 32846 6880 32852
rect 6828 31952 6880 31958
rect 6828 31894 6880 31900
rect 6840 31822 6868 31894
rect 6828 31816 6880 31822
rect 6828 31758 6880 31764
rect 6748 30654 6868 30682
rect 6368 30592 6420 30598
rect 6368 30534 6420 30540
rect 6736 30592 6788 30598
rect 6736 30534 6788 30540
rect 6380 29782 6408 30534
rect 6644 30320 6696 30326
rect 6644 30262 6696 30268
rect 6656 29866 6684 30262
rect 6748 30258 6776 30534
rect 6736 30252 6788 30258
rect 6736 30194 6788 30200
rect 6564 29850 6684 29866
rect 6552 29844 6684 29850
rect 6604 29838 6684 29844
rect 6552 29786 6604 29792
rect 6368 29776 6420 29782
rect 6368 29718 6420 29724
rect 6380 29578 6408 29718
rect 6368 29572 6420 29578
rect 6368 29514 6420 29520
rect 6380 28558 6408 29514
rect 6656 28558 6684 29838
rect 6748 29714 6776 30194
rect 6736 29708 6788 29714
rect 6736 29650 6788 29656
rect 6840 29578 6868 30654
rect 6828 29572 6880 29578
rect 6828 29514 6880 29520
rect 6840 29102 6868 29514
rect 6828 29096 6880 29102
rect 6828 29038 6880 29044
rect 6368 28552 6420 28558
rect 6368 28494 6420 28500
rect 6644 28552 6696 28558
rect 6644 28494 6696 28500
rect 6368 28008 6420 28014
rect 6368 27950 6420 27956
rect 6380 26382 6408 27950
rect 6932 27606 6960 34886
rect 7024 34746 7052 35090
rect 7104 35080 7156 35086
rect 7104 35022 7156 35028
rect 7116 34746 7144 35022
rect 7286 34842 7342 35878
rect 7484 41386 7696 41414
rect 7484 34950 7512 41386
rect 7564 40520 7616 40526
rect 7564 40462 7616 40468
rect 7576 40186 7604 40462
rect 7564 40180 7616 40186
rect 7564 40122 7616 40128
rect 7932 40112 7984 40118
rect 7932 40054 7984 40060
rect 7944 39438 7972 40054
rect 7932 39432 7984 39438
rect 7932 39374 7984 39380
rect 7944 38962 7972 39374
rect 8128 39098 8156 42162
rect 8392 42152 8444 42158
rect 8392 42094 8444 42100
rect 8404 41818 8432 42094
rect 9036 42084 9088 42090
rect 9036 42026 9088 42032
rect 8576 42016 8628 42022
rect 8576 41958 8628 41964
rect 8944 42016 8996 42022
rect 8944 41958 8996 41964
rect 8392 41812 8444 41818
rect 8392 41754 8444 41760
rect 8404 41698 8432 41754
rect 8588 41750 8616 41958
rect 8576 41744 8628 41750
rect 8404 41670 8524 41698
rect 8576 41686 8628 41692
rect 8392 41608 8444 41614
rect 8392 41550 8444 41556
rect 8208 40928 8260 40934
rect 8208 40870 8260 40876
rect 8220 40050 8248 40870
rect 8208 40044 8260 40050
rect 8208 39986 8260 39992
rect 8220 39914 8248 39986
rect 8300 39976 8352 39982
rect 8300 39918 8352 39924
rect 8208 39908 8260 39914
rect 8208 39850 8260 39856
rect 8220 39098 8248 39850
rect 8312 39438 8340 39918
rect 8404 39642 8432 41550
rect 8392 39636 8444 39642
rect 8392 39578 8444 39584
rect 8496 39438 8524 41670
rect 8588 40526 8616 41686
rect 8760 41676 8812 41682
rect 8760 41618 8812 41624
rect 8576 40520 8628 40526
rect 8576 40462 8628 40468
rect 8300 39432 8352 39438
rect 8484 39432 8536 39438
rect 8352 39380 8432 39386
rect 8300 39374 8432 39380
rect 8484 39374 8536 39380
rect 8312 39358 8432 39374
rect 8116 39092 8168 39098
rect 8116 39034 8168 39040
rect 8208 39092 8260 39098
rect 8208 39034 8260 39040
rect 7656 38956 7708 38962
rect 7656 38898 7708 38904
rect 7932 38956 7984 38962
rect 7932 38898 7984 38904
rect 7668 38486 7696 38898
rect 7944 38826 7972 38898
rect 8128 38842 8156 39034
rect 8404 38894 8432 39358
rect 8772 38962 8800 41618
rect 8956 41206 8984 41958
rect 8944 41200 8996 41206
rect 8944 41142 8996 41148
rect 8944 40520 8996 40526
rect 8944 40462 8996 40468
rect 8760 38956 8812 38962
rect 8760 38898 8812 38904
rect 8392 38888 8444 38894
rect 8128 38826 8248 38842
rect 8392 38830 8444 38836
rect 7932 38820 7984 38826
rect 8128 38820 8260 38826
rect 8128 38814 8208 38820
rect 7932 38762 7984 38768
rect 8208 38762 8260 38768
rect 7748 38752 7800 38758
rect 7748 38694 7800 38700
rect 8300 38752 8352 38758
rect 8300 38694 8352 38700
rect 7656 38480 7708 38486
rect 7656 38422 7708 38428
rect 7564 37868 7616 37874
rect 7564 37810 7616 37816
rect 7576 37466 7604 37810
rect 7564 37460 7616 37466
rect 7564 37402 7616 37408
rect 7760 37262 7788 38694
rect 8024 38412 8076 38418
rect 8024 38354 8076 38360
rect 8036 37330 8064 38354
rect 8312 38350 8340 38694
rect 8772 38486 8800 38898
rect 8956 38826 8984 40462
rect 9048 40050 9076 42026
rect 9140 40186 9168 42162
rect 9680 40928 9732 40934
rect 9680 40870 9732 40876
rect 9128 40180 9180 40186
rect 9128 40122 9180 40128
rect 9692 40050 9720 40870
rect 9956 40452 10008 40458
rect 9956 40394 10008 40400
rect 9968 40186 9996 40394
rect 9956 40180 10008 40186
rect 9956 40122 10008 40128
rect 10244 40118 10272 42162
rect 10784 42016 10836 42022
rect 10784 41958 10836 41964
rect 12348 42016 12400 42022
rect 12348 41958 12400 41964
rect 10324 41540 10376 41546
rect 10324 41482 10376 41488
rect 10336 41274 10364 41482
rect 10324 41268 10376 41274
rect 10324 41210 10376 41216
rect 10796 40934 10824 41958
rect 12360 41614 12388 41958
rect 12438 41914 12494 42480
rect 17590 42458 17646 42480
rect 17590 42406 17592 42458
rect 17644 42406 17646 42458
rect 12716 42220 12768 42226
rect 12716 42162 12768 42168
rect 12438 41862 12440 41914
rect 12492 41862 12494 41914
rect 11888 41608 11940 41614
rect 11888 41550 11940 41556
rect 12348 41608 12400 41614
rect 12348 41550 12400 41556
rect 11900 41274 11928 41550
rect 12256 41472 12308 41478
rect 12256 41414 12308 41420
rect 11888 41268 11940 41274
rect 11888 41210 11940 41216
rect 11520 41132 11572 41138
rect 11520 41074 11572 41080
rect 11060 41064 11112 41070
rect 11060 41006 11112 41012
rect 10784 40928 10836 40934
rect 10784 40870 10836 40876
rect 10600 40384 10652 40390
rect 10600 40326 10652 40332
rect 10232 40112 10284 40118
rect 10232 40054 10284 40060
rect 10416 40112 10468 40118
rect 10416 40054 10468 40060
rect 9036 40044 9088 40050
rect 9036 39986 9088 39992
rect 9680 40044 9732 40050
rect 9680 39986 9732 39992
rect 9036 39840 9088 39846
rect 9036 39782 9088 39788
rect 9048 39438 9076 39782
rect 9036 39432 9088 39438
rect 9036 39374 9088 39380
rect 8944 38820 8996 38826
rect 8944 38762 8996 38768
rect 8760 38480 8812 38486
rect 8760 38422 8812 38428
rect 8300 38344 8352 38350
rect 8300 38286 8352 38292
rect 8208 38276 8260 38282
rect 8208 38218 8260 38224
rect 8392 38276 8444 38282
rect 8392 38218 8444 38224
rect 8116 38208 8168 38214
rect 8116 38150 8168 38156
rect 8128 37330 8156 38150
rect 8024 37324 8076 37330
rect 8024 37266 8076 37272
rect 8116 37324 8168 37330
rect 8116 37266 8168 37272
rect 7748 37256 7800 37262
rect 7748 37198 7800 37204
rect 8116 36576 8168 36582
rect 8116 36518 8168 36524
rect 8128 35222 8156 36518
rect 8116 35216 8168 35222
rect 8116 35158 8168 35164
rect 7932 35080 7984 35086
rect 7932 35022 7984 35028
rect 7472 34944 7524 34950
rect 7472 34886 7524 34892
rect 7748 34944 7800 34950
rect 7748 34886 7800 34892
rect 7286 34790 7288 34842
rect 7340 34790 7342 34842
rect 7012 34740 7064 34746
rect 7012 34682 7064 34688
rect 7104 34740 7156 34746
rect 7104 34682 7156 34688
rect 7116 33912 7144 34682
rect 7024 33884 7144 33912
rect 7024 32910 7052 33884
rect 7286 33754 7342 34790
rect 7564 33924 7616 33930
rect 7564 33866 7616 33872
rect 7286 33702 7288 33754
rect 7340 33702 7342 33754
rect 7012 32904 7064 32910
rect 7012 32846 7064 32852
rect 7104 32904 7156 32910
rect 7104 32846 7156 32852
rect 7012 31340 7064 31346
rect 7012 31282 7064 31288
rect 7024 31210 7052 31282
rect 7012 31204 7064 31210
rect 7012 31146 7064 31152
rect 7024 30666 7052 31146
rect 7012 30660 7064 30666
rect 7012 30602 7064 30608
rect 7024 29102 7052 30602
rect 7116 29850 7144 32846
rect 7286 32666 7342 33702
rect 7576 33658 7604 33866
rect 7564 33652 7616 33658
rect 7564 33594 7616 33600
rect 7760 33522 7788 34886
rect 7944 33998 7972 35022
rect 8024 34740 8076 34746
rect 8024 34682 8076 34688
rect 7932 33992 7984 33998
rect 7932 33934 7984 33940
rect 8036 33522 8064 34682
rect 8128 34066 8156 35158
rect 8220 34678 8248 38218
rect 8404 36922 8432 38218
rect 8772 38010 8800 38422
rect 8760 38004 8812 38010
rect 8760 37946 8812 37952
rect 8956 37262 8984 38762
rect 8944 37256 8996 37262
rect 8944 37198 8996 37204
rect 8668 37188 8720 37194
rect 8668 37130 8720 37136
rect 8392 36916 8444 36922
rect 8392 36858 8444 36864
rect 8680 36786 8708 37130
rect 8668 36780 8720 36786
rect 8668 36722 8720 36728
rect 8392 36576 8444 36582
rect 8392 36518 8444 36524
rect 8404 36378 8432 36518
rect 8392 36372 8444 36378
rect 8392 36314 8444 36320
rect 8944 35692 8996 35698
rect 8944 35634 8996 35640
rect 8956 35290 8984 35634
rect 9048 35630 9076 39374
rect 9692 39302 9720 39986
rect 10324 39432 10376 39438
rect 10324 39374 10376 39380
rect 9680 39296 9732 39302
rect 9680 39238 9732 39244
rect 9772 39296 9824 39302
rect 9772 39238 9824 39244
rect 9312 38344 9364 38350
rect 9312 38286 9364 38292
rect 9324 37942 9352 38286
rect 9312 37936 9364 37942
rect 9312 37878 9364 37884
rect 9784 37874 9812 39238
rect 10336 39098 10364 39374
rect 10324 39092 10376 39098
rect 10324 39034 10376 39040
rect 10232 38276 10284 38282
rect 10232 38218 10284 38224
rect 9956 38208 10008 38214
rect 9956 38150 10008 38156
rect 9772 37868 9824 37874
rect 9772 37810 9824 37816
rect 9220 37256 9272 37262
rect 9220 37198 9272 37204
rect 9404 37256 9456 37262
rect 9404 37198 9456 37204
rect 9232 36854 9260 37198
rect 9220 36848 9272 36854
rect 9220 36790 9272 36796
rect 9128 36712 9180 36718
rect 9128 36654 9180 36660
rect 9312 36712 9364 36718
rect 9312 36654 9364 36660
rect 9140 36378 9168 36654
rect 9128 36372 9180 36378
rect 9128 36314 9180 36320
rect 9324 36242 9352 36654
rect 9312 36236 9364 36242
rect 9312 36178 9364 36184
rect 9416 36174 9444 37198
rect 9588 36780 9640 36786
rect 9588 36722 9640 36728
rect 9600 36242 9628 36722
rect 9588 36236 9640 36242
rect 9588 36178 9640 36184
rect 9404 36168 9456 36174
rect 9404 36110 9456 36116
rect 9680 36168 9732 36174
rect 9680 36110 9732 36116
rect 9692 35698 9720 36110
rect 9968 35766 9996 38150
rect 10048 37188 10100 37194
rect 10048 37130 10100 37136
rect 9864 35760 9916 35766
rect 9864 35702 9916 35708
rect 9956 35760 10008 35766
rect 9956 35702 10008 35708
rect 9680 35692 9732 35698
rect 9680 35634 9732 35640
rect 9036 35624 9088 35630
rect 9036 35566 9088 35572
rect 9588 35624 9640 35630
rect 9588 35566 9640 35572
rect 8944 35284 8996 35290
rect 8944 35226 8996 35232
rect 8300 35080 8352 35086
rect 8300 35022 8352 35028
rect 8208 34672 8260 34678
rect 8208 34614 8260 34620
rect 8116 34060 8168 34066
rect 8116 34002 8168 34008
rect 7472 33516 7524 33522
rect 7472 33458 7524 33464
rect 7748 33516 7800 33522
rect 7748 33458 7800 33464
rect 8024 33516 8076 33522
rect 8024 33458 8076 33464
rect 7286 32614 7288 32666
rect 7340 32614 7342 32666
rect 7286 31578 7342 32614
rect 7484 31754 7512 33458
rect 8128 33454 8156 34002
rect 8312 33862 8340 35022
rect 8576 34672 8628 34678
rect 8576 34614 8628 34620
rect 8300 33856 8352 33862
rect 8300 33798 8352 33804
rect 7840 33448 7892 33454
rect 7840 33390 7892 33396
rect 8116 33448 8168 33454
rect 8116 33390 8168 33396
rect 7748 33312 7800 33318
rect 7748 33254 7800 33260
rect 7564 33040 7616 33046
rect 7564 32982 7616 32988
rect 7472 31748 7524 31754
rect 7472 31690 7524 31696
rect 7286 31526 7288 31578
rect 7340 31526 7342 31578
rect 7196 30592 7248 30598
rect 7196 30534 7248 30540
rect 7208 29850 7236 30534
rect 7286 30490 7342 31526
rect 7380 31272 7432 31278
rect 7380 31214 7432 31220
rect 7392 30598 7420 31214
rect 7380 30592 7432 30598
rect 7380 30534 7432 30540
rect 7286 30438 7288 30490
rect 7340 30438 7342 30490
rect 7104 29844 7156 29850
rect 7104 29786 7156 29792
rect 7196 29844 7248 29850
rect 7196 29786 7248 29792
rect 7286 29402 7342 30438
rect 7392 30258 7420 30534
rect 7380 30252 7432 30258
rect 7380 30194 7432 30200
rect 7392 29832 7420 30194
rect 7484 30190 7512 31690
rect 7576 31686 7604 32982
rect 7656 32768 7708 32774
rect 7656 32710 7708 32716
rect 7668 31890 7696 32710
rect 7656 31884 7708 31890
rect 7656 31826 7708 31832
rect 7760 31822 7788 33254
rect 7852 32502 7880 33390
rect 8128 32994 8156 33390
rect 8300 33040 8352 33046
rect 8128 32988 8300 32994
rect 8128 32982 8352 32988
rect 8128 32966 8340 32982
rect 8116 32904 8168 32910
rect 8116 32846 8168 32852
rect 8024 32768 8076 32774
rect 8024 32710 8076 32716
rect 7840 32496 7892 32502
rect 7840 32438 7892 32444
rect 8036 31890 8064 32710
rect 8024 31884 8076 31890
rect 8024 31826 8076 31832
rect 7748 31816 7800 31822
rect 7748 31758 7800 31764
rect 7932 31816 7984 31822
rect 7932 31758 7984 31764
rect 7564 31680 7616 31686
rect 7564 31622 7616 31628
rect 7944 31482 7972 31758
rect 8024 31748 8076 31754
rect 8024 31690 8076 31696
rect 8036 31482 8064 31690
rect 7932 31476 7984 31482
rect 7932 31418 7984 31424
rect 8024 31476 8076 31482
rect 8024 31418 8076 31424
rect 7656 31272 7708 31278
rect 7656 31214 7708 31220
rect 7564 30728 7616 30734
rect 7564 30670 7616 30676
rect 7472 30184 7524 30190
rect 7472 30126 7524 30132
rect 7392 29804 7512 29832
rect 7380 29708 7432 29714
rect 7380 29650 7432 29656
rect 7286 29350 7288 29402
rect 7340 29350 7342 29402
rect 7012 29096 7064 29102
rect 7012 29038 7064 29044
rect 7286 28314 7342 29350
rect 7392 29170 7420 29650
rect 7484 29306 7512 29804
rect 7472 29300 7524 29306
rect 7472 29242 7524 29248
rect 7380 29164 7432 29170
rect 7380 29106 7432 29112
rect 7472 29096 7524 29102
rect 7472 29038 7524 29044
rect 7380 28416 7432 28422
rect 7380 28358 7432 28364
rect 7286 28262 7288 28314
rect 7340 28262 7342 28314
rect 7196 28076 7248 28082
rect 7196 28018 7248 28024
rect 6920 27600 6972 27606
rect 6920 27542 6972 27548
rect 6460 26784 6512 26790
rect 6460 26726 6512 26732
rect 6368 26376 6420 26382
rect 6368 26318 6420 26324
rect 6288 25894 6408 25922
rect 6276 25832 6328 25838
rect 6276 25774 6328 25780
rect 6184 23724 6236 23730
rect 6184 23666 6236 23672
rect 6012 23208 6224 23236
rect 5920 23140 6040 23168
rect 5816 23112 5868 23118
rect 5816 23054 5868 23060
rect 5828 22438 5856 23054
rect 5908 22568 5960 22574
rect 5908 22510 5960 22516
rect 5816 22432 5868 22438
rect 5816 22374 5868 22380
rect 5724 22228 5776 22234
rect 5724 22170 5776 22176
rect 5724 22024 5776 22030
rect 5920 22012 5948 22510
rect 5776 21984 5948 22012
rect 5724 21966 5776 21972
rect 5632 21072 5684 21078
rect 5632 21014 5684 21020
rect 5632 20936 5684 20942
rect 5632 20878 5684 20884
rect 5644 19922 5672 20878
rect 5736 20806 5764 21966
rect 6012 21162 6040 23140
rect 5828 21134 6040 21162
rect 5724 20800 5776 20806
rect 5724 20742 5776 20748
rect 5632 19916 5684 19922
rect 5632 19858 5684 19864
rect 5644 19378 5672 19858
rect 5632 19372 5684 19378
rect 5632 19314 5684 19320
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 5644 17746 5672 19314
rect 5632 17740 5684 17746
rect 5632 17682 5684 17688
rect 5448 17332 5500 17338
rect 5448 17274 5500 17280
rect 5460 16590 5488 17274
rect 5448 16584 5500 16590
rect 5448 16526 5500 16532
rect 5540 16516 5592 16522
rect 5540 16458 5592 16464
rect 5552 16250 5580 16458
rect 5736 16454 5764 20742
rect 5724 16448 5776 16454
rect 5724 16390 5776 16396
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5460 15162 5488 15506
rect 5540 15428 5592 15434
rect 5540 15370 5592 15376
rect 5448 15156 5500 15162
rect 5448 15098 5500 15104
rect 5460 14618 5488 15098
rect 5448 14612 5500 14618
rect 5448 14554 5500 14560
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5448 14272 5500 14278
rect 5448 14214 5500 14220
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 5276 12434 5304 13874
rect 5460 13870 5488 14214
rect 5552 14006 5580 15370
rect 5724 14272 5776 14278
rect 5724 14214 5776 14220
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5356 12912 5408 12918
rect 5356 12854 5408 12860
rect 5184 12406 5304 12434
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 4896 9648 4948 9654
rect 4896 9590 4948 9596
rect 4896 8968 4948 8974
rect 4816 8928 4896 8956
rect 4816 7886 4844 8928
rect 4896 8910 4948 8916
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4816 7478 4844 7822
rect 4804 7472 4856 7478
rect 4804 7414 4856 7420
rect 4804 6928 4856 6934
rect 4804 6870 4856 6876
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4528 5024 4580 5030
rect 4528 4966 4580 4972
rect 4712 4548 4764 4554
rect 4712 4490 4764 4496
rect 4724 4282 4752 4490
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 4528 3596 4580 3602
rect 4528 3538 4580 3544
rect 4344 3528 4396 3534
rect 4344 3470 4396 3476
rect 4356 3126 4384 3470
rect 4344 3120 4396 3126
rect 4344 3062 4396 3068
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 4172 2650 4200 2994
rect 4436 2916 4488 2922
rect 4436 2858 4488 2864
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 4172 1970 4200 2586
rect 4448 2310 4476 2858
rect 4540 2650 4568 3538
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 4528 2644 4580 2650
rect 4528 2586 4580 2592
rect 4436 2304 4488 2310
rect 4436 2246 4488 2252
rect 4724 2038 4752 3334
rect 4816 2854 4844 6870
rect 4804 2848 4856 2854
rect 4804 2790 4856 2796
rect 4712 2032 4764 2038
rect 4712 1974 4764 1980
rect 4068 1964 4120 1970
rect 4068 1906 4120 1912
rect 4160 1964 4212 1970
rect 4160 1906 4212 1912
rect 4908 1358 4936 8230
rect 5000 7342 5028 10610
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 5092 9586 5120 10406
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 5092 7954 5120 8230
rect 5080 7948 5132 7954
rect 5080 7890 5132 7896
rect 4988 7336 5040 7342
rect 5184 7324 5212 12406
rect 5368 12170 5396 12854
rect 5356 12164 5408 12170
rect 5356 12106 5408 12112
rect 5264 11552 5316 11558
rect 5264 11494 5316 11500
rect 5276 11150 5304 11494
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5460 10266 5488 13330
rect 5736 13326 5764 14214
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 5540 13252 5592 13258
rect 5540 13194 5592 13200
rect 5552 11218 5580 13194
rect 5632 12776 5684 12782
rect 5632 12718 5684 12724
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5460 8974 5488 10202
rect 5264 8968 5316 8974
rect 5448 8968 5500 8974
rect 5264 8910 5316 8916
rect 5368 8928 5448 8956
rect 5276 7954 5304 8910
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 5368 7546 5396 8928
rect 5448 8910 5500 8916
rect 5552 8634 5580 11154
rect 5644 10674 5672 12718
rect 5724 12096 5776 12102
rect 5724 12038 5776 12044
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5644 9042 5672 10610
rect 5736 10470 5764 12038
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 4988 7278 5040 7284
rect 5092 7296 5212 7324
rect 5000 5302 5028 7278
rect 5092 5846 5120 7296
rect 5276 7206 5304 7482
rect 5460 7410 5488 7890
rect 5552 7886 5580 8570
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 5080 5840 5132 5846
rect 5080 5782 5132 5788
rect 4988 5296 5040 5302
rect 4988 5238 5040 5244
rect 5092 4570 5120 5782
rect 5000 4542 5120 4570
rect 5000 4282 5028 4542
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 4988 4276 5040 4282
rect 4988 4218 5040 4224
rect 5092 3738 5120 4422
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5184 3534 5212 7142
rect 5460 6798 5488 7346
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5276 5302 5304 6734
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 5368 5370 5396 5578
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5460 5302 5488 6734
rect 5552 5642 5580 6938
rect 5644 5710 5672 7482
rect 5736 7392 5764 9522
rect 5828 7562 5856 21134
rect 5908 21072 5960 21078
rect 5908 21014 5960 21020
rect 5920 18086 5948 21014
rect 6196 20602 6224 23208
rect 6288 22250 6316 25774
rect 6380 24954 6408 25894
rect 6368 24948 6420 24954
rect 6368 24890 6420 24896
rect 6368 24812 6420 24818
rect 6368 24754 6420 24760
rect 6380 24342 6408 24754
rect 6368 24336 6420 24342
rect 6368 24278 6420 24284
rect 6368 23724 6420 23730
rect 6368 23666 6420 23672
rect 6380 22386 6408 23666
rect 6472 22982 6500 26726
rect 6828 26376 6880 26382
rect 6828 26318 6880 26324
rect 6840 25956 6868 26318
rect 6932 26314 6960 27542
rect 7012 27328 7064 27334
rect 7012 27270 7064 27276
rect 7024 26382 7052 27270
rect 7208 27130 7236 28018
rect 7286 27226 7342 28262
rect 7286 27174 7288 27226
rect 7340 27174 7342 27226
rect 7196 27124 7248 27130
rect 7196 27066 7248 27072
rect 7104 26580 7156 26586
rect 7104 26522 7156 26528
rect 7116 26466 7144 26522
rect 7116 26438 7236 26466
rect 7012 26376 7064 26382
rect 7012 26318 7064 26324
rect 6920 26308 6972 26314
rect 6920 26250 6972 26256
rect 6920 25968 6972 25974
rect 6840 25928 6920 25956
rect 6552 25696 6604 25702
rect 6552 25638 6604 25644
rect 6736 25696 6788 25702
rect 6736 25638 6788 25644
rect 6564 25498 6592 25638
rect 6552 25492 6604 25498
rect 6552 25434 6604 25440
rect 6552 25356 6604 25362
rect 6552 25298 6604 25304
rect 6564 24614 6592 25298
rect 6644 24812 6696 24818
rect 6644 24754 6696 24760
rect 6552 24608 6604 24614
rect 6552 24550 6604 24556
rect 6656 23866 6684 24754
rect 6748 24274 6776 25638
rect 6840 24818 6868 25928
rect 6920 25910 6972 25916
rect 7208 25294 7236 26438
rect 7286 26138 7342 27174
rect 7392 26994 7420 28358
rect 7484 28014 7512 29038
rect 7472 28008 7524 28014
rect 7472 27950 7524 27956
rect 7472 27600 7524 27606
rect 7472 27542 7524 27548
rect 7484 26994 7512 27542
rect 7380 26988 7432 26994
rect 7380 26930 7432 26936
rect 7472 26988 7524 26994
rect 7472 26930 7524 26936
rect 7380 26784 7432 26790
rect 7380 26726 7432 26732
rect 7286 26086 7288 26138
rect 7340 26086 7342 26138
rect 7196 25288 7248 25294
rect 7196 25230 7248 25236
rect 7208 24954 7236 25230
rect 7286 25050 7342 26086
rect 7286 24998 7288 25050
rect 7340 24998 7342 25050
rect 7196 24948 7248 24954
rect 7196 24890 7248 24896
rect 6828 24812 6880 24818
rect 6828 24754 6880 24760
rect 6840 24682 6868 24754
rect 6828 24676 6880 24682
rect 6828 24618 6880 24624
rect 6736 24268 6788 24274
rect 6736 24210 6788 24216
rect 6644 23860 6696 23866
rect 6644 23802 6696 23808
rect 6552 23656 6604 23662
rect 6552 23598 6604 23604
rect 6460 22976 6512 22982
rect 6460 22918 6512 22924
rect 6380 22358 6500 22386
rect 6288 22222 6408 22250
rect 6276 21888 6328 21894
rect 6276 21830 6328 21836
rect 6184 20596 6236 20602
rect 6184 20538 6236 20544
rect 6000 20052 6052 20058
rect 6000 19994 6052 20000
rect 6012 18630 6040 19994
rect 6092 19508 6144 19514
rect 6092 19450 6144 19456
rect 6000 18624 6052 18630
rect 6000 18566 6052 18572
rect 6104 18426 6132 19450
rect 6092 18420 6144 18426
rect 6092 18362 6144 18368
rect 5908 18080 5960 18086
rect 5908 18022 5960 18028
rect 6000 16108 6052 16114
rect 6000 16050 6052 16056
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 5920 12442 5948 12786
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 6012 11014 6040 16050
rect 6092 15156 6144 15162
rect 6092 15098 6144 15104
rect 6104 14482 6132 15098
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 6196 14278 6224 20538
rect 6288 15366 6316 21830
rect 6380 20058 6408 22222
rect 6472 21690 6500 22358
rect 6460 21684 6512 21690
rect 6460 21626 6512 21632
rect 6460 21548 6512 21554
rect 6460 21490 6512 21496
rect 6368 20052 6420 20058
rect 6368 19994 6420 20000
rect 6368 19780 6420 19786
rect 6368 19722 6420 19728
rect 6380 18426 6408 19722
rect 6472 19242 6500 21490
rect 6460 19236 6512 19242
rect 6460 19178 6512 19184
rect 6460 18624 6512 18630
rect 6460 18566 6512 18572
rect 6368 18420 6420 18426
rect 6368 18362 6420 18368
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 6276 15360 6328 15366
rect 6276 15302 6328 15308
rect 6276 14476 6328 14482
rect 6276 14418 6328 14424
rect 6184 14272 6236 14278
rect 6184 14214 6236 14220
rect 6196 14006 6224 14214
rect 6184 14000 6236 14006
rect 6184 13942 6236 13948
rect 6184 13184 6236 13190
rect 6184 13126 6236 13132
rect 6196 12442 6224 13126
rect 6288 12850 6316 14418
rect 6276 12844 6328 12850
rect 6276 12786 6328 12792
rect 6184 12436 6236 12442
rect 6184 12378 6236 12384
rect 6276 12300 6328 12306
rect 6276 12242 6328 12248
rect 6092 11688 6144 11694
rect 6092 11630 6144 11636
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 6012 10062 6040 10610
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 6012 8906 6040 9862
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 6000 8424 6052 8430
rect 6000 8366 6052 8372
rect 5828 7534 5948 7562
rect 6012 7546 6040 8366
rect 5816 7404 5868 7410
rect 5736 7364 5816 7392
rect 5816 7346 5868 7352
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5540 5636 5592 5642
rect 5540 5578 5592 5584
rect 5264 5296 5316 5302
rect 5264 5238 5316 5244
rect 5448 5296 5500 5302
rect 5448 5238 5500 5244
rect 5276 4826 5304 5238
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5264 4480 5316 4486
rect 5264 4422 5316 4428
rect 5276 4214 5304 4422
rect 5264 4208 5316 4214
rect 5264 4150 5316 4156
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5460 3738 5488 4082
rect 5828 4010 5856 7346
rect 5816 4004 5868 4010
rect 5816 3946 5868 3952
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5736 3738 5764 3878
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 3884 1352 3936 1358
rect 3884 1294 3936 1300
rect 4896 1352 4948 1358
rect 4896 1294 4948 1300
rect 5736 1290 5764 3674
rect 5920 2774 5948 7534
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 6000 7268 6052 7274
rect 6000 7210 6052 7216
rect 6012 6322 6040 7210
rect 6104 7206 6132 11630
rect 6184 11552 6236 11558
rect 6184 11494 6236 11500
rect 6196 11082 6224 11494
rect 6184 11076 6236 11082
rect 6184 11018 6236 11024
rect 6288 10198 6316 12242
rect 6380 11336 6408 16186
rect 6472 12374 6500 18566
rect 6564 17678 6592 23598
rect 6644 23588 6696 23594
rect 6644 23530 6696 23536
rect 6656 23118 6684 23530
rect 6748 23186 6776 24210
rect 6840 23526 6868 24618
rect 6920 24200 6972 24206
rect 6920 24142 6972 24148
rect 6932 23866 6960 24142
rect 7196 24132 7248 24138
rect 7196 24074 7248 24080
rect 6920 23860 6972 23866
rect 6920 23802 6972 23808
rect 6828 23520 6880 23526
rect 6828 23462 6880 23468
rect 6736 23180 6788 23186
rect 6736 23122 6788 23128
rect 6644 23112 6696 23118
rect 6644 23054 6696 23060
rect 6656 22778 6684 23054
rect 6644 22772 6696 22778
rect 6644 22714 6696 22720
rect 6840 22710 6868 23462
rect 6828 22704 6880 22710
rect 6828 22646 6880 22652
rect 6736 22432 6788 22438
rect 6736 22374 6788 22380
rect 6748 21418 6776 22374
rect 6932 22094 6960 23802
rect 7104 22976 7156 22982
rect 7104 22918 7156 22924
rect 6932 22066 7052 22094
rect 6920 21956 6972 21962
rect 6920 21898 6972 21904
rect 6932 21486 6960 21898
rect 6920 21480 6972 21486
rect 6920 21422 6972 21428
rect 6736 21412 6788 21418
rect 6736 21354 6788 21360
rect 7024 21026 7052 22066
rect 6932 20998 7052 21026
rect 6736 20936 6788 20942
rect 6736 20878 6788 20884
rect 6828 20936 6880 20942
rect 6828 20878 6880 20884
rect 6644 20528 6696 20534
rect 6644 20470 6696 20476
rect 6656 19310 6684 20470
rect 6644 19304 6696 19310
rect 6644 19246 6696 19252
rect 6656 18970 6684 19246
rect 6644 18964 6696 18970
rect 6644 18906 6696 18912
rect 6656 18154 6684 18906
rect 6748 18630 6776 20878
rect 6840 20602 6868 20878
rect 6828 20596 6880 20602
rect 6828 20538 6880 20544
rect 6840 19514 6868 20538
rect 6932 20466 6960 20998
rect 7012 20868 7064 20874
rect 7012 20810 7064 20816
rect 6920 20460 6972 20466
rect 6920 20402 6972 20408
rect 6932 20262 6960 20402
rect 6920 20256 6972 20262
rect 6920 20198 6972 20204
rect 7024 20058 7052 20810
rect 7012 20052 7064 20058
rect 7012 19994 7064 20000
rect 7024 19514 7052 19994
rect 6828 19508 6880 19514
rect 6828 19450 6880 19456
rect 7012 19508 7064 19514
rect 7012 19450 7064 19456
rect 7024 18834 7052 19450
rect 7012 18828 7064 18834
rect 7012 18770 7064 18776
rect 7116 18714 7144 22918
rect 7208 21010 7236 24074
rect 7286 23962 7342 24998
rect 7286 23910 7288 23962
rect 7340 23910 7342 23962
rect 7286 22874 7342 23910
rect 7286 22822 7288 22874
rect 7340 22822 7342 22874
rect 7286 21786 7342 22822
rect 7286 21734 7288 21786
rect 7340 21734 7342 21786
rect 7196 21004 7248 21010
rect 7196 20946 7248 20952
rect 7286 20698 7342 21734
rect 7286 20646 7288 20698
rect 7340 20646 7342 20698
rect 7286 19610 7342 20646
rect 7392 20534 7420 26726
rect 7472 21888 7524 21894
rect 7472 21830 7524 21836
rect 7484 20942 7512 21830
rect 7472 20936 7524 20942
rect 7472 20878 7524 20884
rect 7380 20528 7432 20534
rect 7380 20470 7432 20476
rect 7380 20256 7432 20262
rect 7380 20198 7432 20204
rect 7286 19558 7288 19610
rect 7340 19558 7342 19610
rect 7196 18896 7248 18902
rect 7196 18838 7248 18844
rect 6840 18686 7144 18714
rect 6736 18624 6788 18630
rect 6736 18566 6788 18572
rect 6840 18442 6868 18686
rect 6748 18414 6868 18442
rect 7208 18426 7236 18838
rect 7286 18522 7342 19558
rect 7286 18470 7288 18522
rect 7340 18470 7342 18522
rect 7196 18420 7248 18426
rect 6644 18148 6696 18154
rect 6644 18090 6696 18096
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 6552 16584 6604 16590
rect 6552 16526 6604 16532
rect 6564 15570 6592 16526
rect 6748 16454 6776 18414
rect 7196 18362 7248 18368
rect 7104 18352 7156 18358
rect 7104 18294 7156 18300
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 6840 16640 6868 17818
rect 6920 17604 6972 17610
rect 6920 17546 6972 17552
rect 6932 16794 6960 17546
rect 7012 16992 7064 16998
rect 7012 16934 7064 16940
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 6840 16612 6960 16640
rect 6736 16448 6788 16454
rect 6736 16390 6788 16396
rect 6644 15904 6696 15910
rect 6644 15846 6696 15852
rect 6656 15638 6684 15846
rect 6644 15632 6696 15638
rect 6644 15574 6696 15580
rect 6552 15564 6604 15570
rect 6552 15506 6604 15512
rect 6828 15564 6880 15570
rect 6828 15506 6880 15512
rect 6736 15360 6788 15366
rect 6736 15302 6788 15308
rect 6552 14272 6604 14278
rect 6552 14214 6604 14220
rect 6564 13802 6592 14214
rect 6552 13796 6604 13802
rect 6552 13738 6604 13744
rect 6748 13274 6776 15302
rect 6840 15094 6868 15506
rect 6828 15088 6880 15094
rect 6828 15030 6880 15036
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 6840 13394 6868 14554
rect 6932 14498 6960 16612
rect 7024 14958 7052 16934
rect 7012 14952 7064 14958
rect 7012 14894 7064 14900
rect 6932 14470 7052 14498
rect 6920 14340 6972 14346
rect 6920 14282 6972 14288
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 6932 13326 6960 14282
rect 6920 13320 6972 13326
rect 6748 13246 6868 13274
rect 6920 13262 6972 13268
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6460 12368 6512 12374
rect 6460 12310 6512 12316
rect 6460 12232 6512 12238
rect 6564 12220 6592 12718
rect 6644 12368 6696 12374
rect 6644 12310 6696 12316
rect 6656 12238 6684 12310
rect 6512 12192 6592 12220
rect 6644 12232 6696 12238
rect 6460 12174 6512 12180
rect 6644 12174 6696 12180
rect 6656 11694 6684 12174
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 6380 11308 6684 11336
rect 6368 11212 6420 11218
rect 6368 11154 6420 11160
rect 6276 10192 6328 10198
rect 6276 10134 6328 10140
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6288 8974 6316 9318
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 6276 8492 6328 8498
rect 6276 8434 6328 8440
rect 6184 8016 6236 8022
rect 6184 7958 6236 7964
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 6092 5772 6144 5778
rect 6092 5714 6144 5720
rect 6104 5030 6132 5714
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 6104 3738 6132 4966
rect 6196 4758 6224 7958
rect 6288 7546 6316 8434
rect 6276 7540 6328 7546
rect 6276 7482 6328 7488
rect 6380 5846 6408 11154
rect 6460 11076 6512 11082
rect 6460 11018 6512 11024
rect 6552 11076 6604 11082
rect 6552 11018 6604 11024
rect 6472 10266 6500 11018
rect 6460 10260 6512 10266
rect 6460 10202 6512 10208
rect 6564 9586 6592 11018
rect 6656 9722 6684 11308
rect 6736 11076 6788 11082
rect 6736 11018 6788 11024
rect 6748 10810 6776 11018
rect 6736 10804 6788 10810
rect 6736 10746 6788 10752
rect 6736 10056 6788 10062
rect 6736 9998 6788 10004
rect 6644 9716 6696 9722
rect 6644 9658 6696 9664
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6644 8900 6696 8906
rect 6644 8842 6696 8848
rect 6460 8492 6512 8498
rect 6460 8434 6512 8440
rect 6472 8090 6500 8434
rect 6656 8294 6684 8842
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6564 7410 6592 7686
rect 6656 7410 6684 8230
rect 6748 7954 6776 9998
rect 6840 9654 6868 13246
rect 7024 12102 7052 14470
rect 7116 13530 7144 18294
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7208 17338 7236 17478
rect 7286 17434 7342 18470
rect 7392 18306 7420 20198
rect 7484 18426 7512 20878
rect 7576 20874 7604 30670
rect 7668 29646 7696 31214
rect 7748 30864 7800 30870
rect 7748 30806 7800 30812
rect 7656 29640 7708 29646
rect 7656 29582 7708 29588
rect 7668 26790 7696 29582
rect 7760 28150 7788 30806
rect 7932 30796 7984 30802
rect 7932 30738 7984 30744
rect 7944 29510 7972 30738
rect 7932 29504 7984 29510
rect 7932 29446 7984 29452
rect 8036 29322 8064 31418
rect 8128 31278 8156 32846
rect 8208 32496 8260 32502
rect 8208 32438 8260 32444
rect 8220 31804 8248 32438
rect 8300 31816 8352 31822
rect 8220 31776 8300 31804
rect 8116 31272 8168 31278
rect 8116 31214 8168 31220
rect 8220 30938 8248 31776
rect 8300 31758 8352 31764
rect 8208 30932 8260 30938
rect 8208 30874 8260 30880
rect 8116 30728 8168 30734
rect 8116 30670 8168 30676
rect 8300 30728 8352 30734
rect 8300 30670 8352 30676
rect 7944 29294 8064 29322
rect 7944 29170 7972 29294
rect 7932 29164 7984 29170
rect 7932 29106 7984 29112
rect 7944 28694 7972 29106
rect 8128 28966 8156 30670
rect 8312 30326 8340 30670
rect 8484 30388 8536 30394
rect 8484 30330 8536 30336
rect 8300 30320 8352 30326
rect 8300 30262 8352 30268
rect 8496 30258 8524 30330
rect 8208 30252 8260 30258
rect 8208 30194 8260 30200
rect 8484 30252 8536 30258
rect 8484 30194 8536 30200
rect 8220 29782 8248 30194
rect 8392 30048 8444 30054
rect 8392 29990 8444 29996
rect 8208 29776 8260 29782
rect 8208 29718 8260 29724
rect 8300 29776 8352 29782
rect 8300 29718 8352 29724
rect 8220 29510 8248 29718
rect 8208 29504 8260 29510
rect 8208 29446 8260 29452
rect 8208 29028 8260 29034
rect 8208 28970 8260 28976
rect 8116 28960 8168 28966
rect 8116 28902 8168 28908
rect 8220 28762 8248 28970
rect 8208 28756 8260 28762
rect 8208 28698 8260 28704
rect 7932 28688 7984 28694
rect 7932 28630 7984 28636
rect 8116 28620 8168 28626
rect 8116 28562 8168 28568
rect 7932 28552 7984 28558
rect 7932 28494 7984 28500
rect 7748 28144 7800 28150
rect 7748 28086 7800 28092
rect 7656 26784 7708 26790
rect 7656 26726 7708 26732
rect 7760 25906 7788 28086
rect 7944 28082 7972 28494
rect 7932 28076 7984 28082
rect 7932 28018 7984 28024
rect 7840 27872 7892 27878
rect 7840 27814 7892 27820
rect 7852 27538 7880 27814
rect 7840 27532 7892 27538
rect 7840 27474 7892 27480
rect 7944 27470 7972 28018
rect 8128 27946 8156 28562
rect 8208 28552 8260 28558
rect 8208 28494 8260 28500
rect 8220 28218 8248 28494
rect 8208 28212 8260 28218
rect 8208 28154 8260 28160
rect 8116 27940 8168 27946
rect 8116 27882 8168 27888
rect 8220 27470 8248 28154
rect 7932 27464 7984 27470
rect 7932 27406 7984 27412
rect 8208 27464 8260 27470
rect 8208 27406 8260 27412
rect 7840 26988 7892 26994
rect 7840 26930 7892 26936
rect 7852 26586 7880 26930
rect 8116 26920 8168 26926
rect 8116 26862 8168 26868
rect 7840 26580 7892 26586
rect 7840 26522 7892 26528
rect 8128 26382 8156 26862
rect 8116 26376 8168 26382
rect 8116 26318 8168 26324
rect 7748 25900 7800 25906
rect 7748 25842 7800 25848
rect 7656 24200 7708 24206
rect 7656 24142 7708 24148
rect 7668 22710 7696 24142
rect 8024 23316 8076 23322
rect 8024 23258 8076 23264
rect 7932 23112 7984 23118
rect 7932 23054 7984 23060
rect 7840 22976 7892 22982
rect 7840 22918 7892 22924
rect 7656 22704 7708 22710
rect 7656 22646 7708 22652
rect 7564 20868 7616 20874
rect 7564 20810 7616 20816
rect 7668 20754 7696 22646
rect 7748 22024 7800 22030
rect 7748 21966 7800 21972
rect 7760 20924 7788 21966
rect 7852 21554 7880 22918
rect 7944 22234 7972 23054
rect 7932 22228 7984 22234
rect 7932 22170 7984 22176
rect 8036 22094 8064 23258
rect 8128 22642 8156 26318
rect 8208 25764 8260 25770
rect 8208 25706 8260 25712
rect 8220 25294 8248 25706
rect 8312 25378 8340 29718
rect 8404 27878 8432 29990
rect 8496 29782 8524 30194
rect 8484 29776 8536 29782
rect 8484 29718 8536 29724
rect 8484 28008 8536 28014
rect 8484 27950 8536 27956
rect 8392 27872 8444 27878
rect 8392 27814 8444 27820
rect 8404 26586 8432 27814
rect 8496 27674 8524 27950
rect 8484 27668 8536 27674
rect 8484 27610 8536 27616
rect 8392 26580 8444 26586
rect 8392 26522 8444 26528
rect 8312 25350 8432 25378
rect 8208 25288 8260 25294
rect 8208 25230 8260 25236
rect 8208 24812 8260 24818
rect 8208 24754 8260 24760
rect 8220 23322 8248 24754
rect 8404 24052 8432 25350
rect 8484 24608 8536 24614
rect 8484 24550 8536 24556
rect 8496 24206 8524 24550
rect 8484 24200 8536 24206
rect 8484 24142 8536 24148
rect 8404 24024 8524 24052
rect 8300 23792 8352 23798
rect 8300 23734 8352 23740
rect 8208 23316 8260 23322
rect 8208 23258 8260 23264
rect 8312 23254 8340 23734
rect 8300 23248 8352 23254
rect 8300 23190 8352 23196
rect 8116 22636 8168 22642
rect 8116 22578 8168 22584
rect 8036 22066 8156 22094
rect 8024 22024 8076 22030
rect 8024 21966 8076 21972
rect 7932 21888 7984 21894
rect 7932 21830 7984 21836
rect 7840 21548 7892 21554
rect 7840 21490 7892 21496
rect 7840 20936 7892 20942
rect 7760 20896 7840 20924
rect 7840 20878 7892 20884
rect 7576 20726 7696 20754
rect 7576 19446 7604 20726
rect 7656 20324 7708 20330
rect 7656 20266 7708 20272
rect 7668 19718 7696 20266
rect 7656 19712 7708 19718
rect 7656 19654 7708 19660
rect 7564 19440 7616 19446
rect 7564 19382 7616 19388
rect 7564 18692 7616 18698
rect 7564 18634 7616 18640
rect 7576 18426 7604 18634
rect 7748 18624 7800 18630
rect 7748 18566 7800 18572
rect 7472 18420 7524 18426
rect 7472 18362 7524 18368
rect 7564 18420 7616 18426
rect 7564 18362 7616 18368
rect 7392 18278 7604 18306
rect 7760 18290 7788 18566
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7286 17382 7288 17434
rect 7340 17382 7342 17434
rect 7196 17332 7248 17338
rect 7196 17274 7248 17280
rect 7208 16590 7236 17274
rect 7196 16584 7248 16590
rect 7196 16526 7248 16532
rect 7208 15978 7236 16526
rect 7286 16346 7342 17382
rect 7392 16998 7420 17818
rect 7576 17762 7604 18278
rect 7656 18284 7708 18290
rect 7656 18226 7708 18232
rect 7748 18284 7800 18290
rect 7748 18226 7800 18232
rect 7668 17882 7696 18226
rect 7656 17876 7708 17882
rect 7656 17818 7708 17824
rect 7576 17734 7696 17762
rect 7472 17060 7524 17066
rect 7472 17002 7524 17008
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7380 16584 7432 16590
rect 7380 16526 7432 16532
rect 7286 16294 7288 16346
rect 7340 16294 7342 16346
rect 7196 15972 7248 15978
rect 7196 15914 7248 15920
rect 7208 15502 7236 15914
rect 7196 15496 7248 15502
rect 7196 15438 7248 15444
rect 7286 15258 7342 16294
rect 7392 16250 7420 16526
rect 7380 16244 7432 16250
rect 7380 16186 7432 16192
rect 7484 16130 7512 17002
rect 7564 16584 7616 16590
rect 7564 16526 7616 16532
rect 7392 16102 7512 16130
rect 7576 16114 7604 16526
rect 7564 16108 7616 16114
rect 7392 15910 7420 16102
rect 7564 16050 7616 16056
rect 7472 16040 7524 16046
rect 7472 15982 7524 15988
rect 7380 15904 7432 15910
rect 7380 15846 7432 15852
rect 7286 15206 7288 15258
rect 7340 15206 7342 15258
rect 7196 14816 7248 14822
rect 7196 14758 7248 14764
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 7116 12918 7144 13126
rect 7104 12912 7156 12918
rect 7104 12854 7156 12860
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 7208 11762 7236 14758
rect 7286 14170 7342 15206
rect 7392 14822 7420 15846
rect 7484 15706 7512 15982
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7576 15552 7604 16050
rect 7484 15524 7604 15552
rect 7484 14822 7512 15524
rect 7668 15484 7696 17734
rect 7760 17202 7788 18226
rect 7748 17196 7800 17202
rect 7748 17138 7800 17144
rect 7760 15638 7788 17138
rect 7852 16658 7880 20878
rect 7944 18578 7972 21830
rect 8036 21486 8064 21966
rect 8024 21480 8076 21486
rect 8024 21422 8076 21428
rect 8128 20618 8156 22066
rect 8300 22024 8352 22030
rect 8300 21966 8352 21972
rect 8312 20754 8340 21966
rect 8392 21888 8444 21894
rect 8392 21830 8444 21836
rect 8404 21554 8432 21830
rect 8392 21548 8444 21554
rect 8392 21490 8444 21496
rect 8312 20726 8432 20754
rect 8128 20590 8340 20618
rect 8116 20528 8168 20534
rect 8116 20470 8168 20476
rect 8024 20460 8076 20466
rect 8024 20402 8076 20408
rect 8036 19700 8064 20402
rect 8128 20330 8156 20470
rect 8208 20460 8260 20466
rect 8208 20402 8260 20408
rect 8116 20324 8168 20330
rect 8116 20266 8168 20272
rect 8116 19712 8168 19718
rect 8036 19672 8116 19700
rect 8036 18766 8064 19672
rect 8116 19654 8168 19660
rect 8220 19514 8248 20402
rect 8208 19508 8260 19514
rect 8208 19450 8260 19456
rect 8312 19394 8340 20590
rect 8404 20482 8432 20726
rect 8496 20602 8524 24024
rect 8588 20942 8616 34614
rect 8944 33856 8996 33862
rect 8944 33798 8996 33804
rect 8956 32842 8984 33798
rect 8944 32836 8996 32842
rect 8944 32778 8996 32784
rect 8944 32224 8996 32230
rect 8944 32166 8996 32172
rect 8956 32026 8984 32166
rect 8944 32020 8996 32026
rect 8944 31962 8996 31968
rect 9048 31686 9076 35566
rect 9220 35488 9272 35494
rect 9220 35430 9272 35436
rect 9128 35080 9180 35086
rect 9128 35022 9180 35028
rect 9140 34202 9168 35022
rect 9128 34196 9180 34202
rect 9128 34138 9180 34144
rect 9128 33992 9180 33998
rect 9128 33934 9180 33940
rect 9140 33522 9168 33934
rect 9232 33930 9260 35430
rect 9600 35018 9628 35566
rect 9876 35086 9904 35702
rect 10060 35562 10088 37130
rect 10244 36650 10272 38218
rect 10324 37120 10376 37126
rect 10324 37062 10376 37068
rect 10336 36922 10364 37062
rect 10324 36916 10376 36922
rect 10324 36858 10376 36864
rect 10232 36644 10284 36650
rect 10232 36586 10284 36592
rect 10324 36372 10376 36378
rect 10324 36314 10376 36320
rect 10336 36038 10364 36314
rect 10324 36032 10376 36038
rect 10324 35974 10376 35980
rect 10048 35556 10100 35562
rect 10048 35498 10100 35504
rect 9864 35080 9916 35086
rect 9864 35022 9916 35028
rect 9404 35012 9456 35018
rect 9404 34954 9456 34960
rect 9588 35012 9640 35018
rect 9588 34954 9640 34960
rect 9416 33998 9444 34954
rect 9876 34678 9904 35022
rect 9864 34672 9916 34678
rect 9864 34614 9916 34620
rect 10048 34604 10100 34610
rect 10048 34546 10100 34552
rect 10060 34202 10088 34546
rect 10048 34196 10100 34202
rect 10048 34138 10100 34144
rect 9404 33992 9456 33998
rect 9404 33934 9456 33940
rect 10232 33992 10284 33998
rect 10232 33934 10284 33940
rect 9220 33924 9272 33930
rect 9220 33866 9272 33872
rect 9128 33516 9180 33522
rect 9128 33458 9180 33464
rect 9232 32434 9260 33866
rect 9416 33538 9444 33934
rect 10244 33658 10272 33934
rect 10232 33652 10284 33658
rect 10232 33594 10284 33600
rect 9324 33522 9444 33538
rect 9312 33516 9444 33522
rect 9364 33510 9444 33516
rect 9312 33458 9364 33464
rect 9956 33448 10008 33454
rect 9956 33390 10008 33396
rect 9864 32836 9916 32842
rect 9864 32778 9916 32784
rect 9312 32768 9364 32774
rect 9312 32710 9364 32716
rect 9324 32570 9352 32710
rect 9312 32564 9364 32570
rect 9312 32506 9364 32512
rect 9220 32428 9272 32434
rect 9220 32370 9272 32376
rect 9324 31754 9352 32506
rect 9404 32360 9456 32366
rect 9404 32302 9456 32308
rect 9416 31754 9444 32302
rect 9312 31748 9364 31754
rect 9312 31690 9364 31696
rect 9404 31748 9456 31754
rect 9404 31690 9456 31696
rect 9036 31680 9088 31686
rect 9036 31622 9088 31628
rect 8668 31272 8720 31278
rect 8668 31214 8720 31220
rect 8680 31142 8708 31214
rect 8668 31136 8720 31142
rect 8668 31078 8720 31084
rect 8852 31136 8904 31142
rect 8852 31078 8904 31084
rect 8680 30394 8708 31078
rect 8864 30734 8892 31078
rect 8852 30728 8904 30734
rect 8852 30670 8904 30676
rect 8668 30388 8720 30394
rect 8668 30330 8720 30336
rect 8680 29782 8708 30330
rect 8760 30048 8812 30054
rect 8760 29990 8812 29996
rect 8668 29776 8720 29782
rect 8668 29718 8720 29724
rect 8668 29572 8720 29578
rect 8668 29514 8720 29520
rect 8680 28132 8708 29514
rect 8772 28626 8800 29990
rect 8760 28620 8812 28626
rect 8760 28562 8812 28568
rect 8760 28144 8812 28150
rect 8680 28104 8760 28132
rect 8760 28086 8812 28092
rect 8760 26988 8812 26994
rect 8760 26930 8812 26936
rect 8668 24812 8720 24818
rect 8668 24754 8720 24760
rect 8680 21146 8708 24754
rect 8772 24410 8800 26930
rect 8760 24404 8812 24410
rect 8760 24346 8812 24352
rect 8668 21140 8720 21146
rect 8668 21082 8720 21088
rect 8576 20936 8628 20942
rect 8576 20878 8628 20884
rect 8576 20800 8628 20806
rect 8576 20742 8628 20748
rect 8484 20596 8536 20602
rect 8484 20538 8536 20544
rect 8395 20454 8432 20482
rect 8395 20380 8423 20454
rect 8395 20352 8432 20380
rect 8404 19922 8432 20352
rect 8484 20256 8536 20262
rect 8484 20198 8536 20204
rect 8392 19916 8444 19922
rect 8392 19858 8444 19864
rect 8220 19366 8340 19394
rect 8024 18760 8076 18766
rect 8024 18702 8076 18708
rect 7944 18550 8156 18578
rect 7932 18284 7984 18290
rect 7932 18226 7984 18232
rect 8024 18284 8076 18290
rect 8024 18226 8076 18232
rect 7944 17338 7972 18226
rect 8036 17338 8064 18226
rect 7932 17332 7984 17338
rect 7932 17274 7984 17280
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 8024 17060 8076 17066
rect 8024 17002 8076 17008
rect 7840 16652 7892 16658
rect 7840 16594 7892 16600
rect 7840 16108 7892 16114
rect 7840 16050 7892 16056
rect 7748 15632 7800 15638
rect 7748 15574 7800 15580
rect 7576 15456 7696 15484
rect 7380 14816 7432 14822
rect 7380 14758 7432 14764
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 7286 14118 7288 14170
rect 7340 14118 7342 14170
rect 7286 13082 7342 14118
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7286 13030 7288 13082
rect 7340 13030 7342 13082
rect 7286 11994 7342 13030
rect 7380 12368 7432 12374
rect 7380 12310 7432 12316
rect 7286 11942 7288 11994
rect 7340 11942 7342 11994
rect 7196 11756 7248 11762
rect 7196 11698 7248 11704
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 7116 11014 7144 11630
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 6828 9648 6880 9654
rect 6828 9590 6880 9596
rect 6932 8974 6960 10474
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6932 8634 6960 8910
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 6736 7948 6788 7954
rect 6736 7890 6788 7896
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6932 7342 6960 7754
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6644 6724 6696 6730
rect 6644 6666 6696 6672
rect 6656 6390 6684 6666
rect 6644 6384 6696 6390
rect 6644 6326 6696 6332
rect 6932 6254 6960 7278
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 6368 5840 6420 5846
rect 6368 5782 6420 5788
rect 6380 5148 6408 5782
rect 6932 5658 6960 6190
rect 6840 5630 6960 5658
rect 6840 5386 6868 5630
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6564 5358 6868 5386
rect 6932 5370 6960 5510
rect 6920 5364 6972 5370
rect 6564 5234 6592 5358
rect 6920 5306 6972 5312
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6460 5160 6512 5166
rect 6288 5120 6460 5148
rect 6184 4752 6236 4758
rect 6184 4694 6236 4700
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 6092 3460 6144 3466
rect 6092 3402 6144 3408
rect 6104 3126 6132 3402
rect 6092 3120 6144 3126
rect 6092 3062 6144 3068
rect 6196 2922 6224 4694
rect 6288 3602 6316 5120
rect 6460 5102 6512 5108
rect 6368 4480 6420 4486
rect 6368 4422 6420 4428
rect 6276 3596 6328 3602
rect 6276 3538 6328 3544
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 6184 2916 6236 2922
rect 6184 2858 6236 2864
rect 5920 2746 6224 2774
rect 6196 1442 6224 2746
rect 6288 1562 6316 2994
rect 6276 1556 6328 1562
rect 6276 1498 6328 1504
rect 6196 1414 6316 1442
rect 5816 1352 5868 1358
rect 5816 1294 5868 1300
rect 5724 1284 5776 1290
rect 5724 1226 5776 1232
rect 3240 1216 3292 1222
rect 3240 1158 3292 1164
rect 5632 1216 5684 1222
rect 5632 1158 5684 1164
rect 5644 814 5672 1158
rect 5828 1018 5856 1294
rect 5816 1012 5868 1018
rect 5816 954 5868 960
rect 5632 808 5684 814
rect 2778 0 2834 800
rect 5632 750 5684 756
rect 6288 746 6316 1414
rect 6380 1358 6408 4422
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6472 2922 6500 3402
rect 6564 3058 6592 5170
rect 6644 4752 6696 4758
rect 6644 4694 6696 4700
rect 6656 4622 6684 4694
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6736 4548 6788 4554
rect 6736 4490 6788 4496
rect 6748 4010 6776 4490
rect 6736 4004 6788 4010
rect 6736 3946 6788 3952
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6656 3466 6684 3878
rect 6644 3460 6696 3466
rect 6644 3402 6696 3408
rect 6748 3058 6776 3946
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6840 3040 6868 3538
rect 6932 3534 6960 3878
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6920 3052 6972 3058
rect 6840 3012 6920 3040
rect 6460 2916 6512 2922
rect 6460 2858 6512 2864
rect 6564 2446 6592 2994
rect 6748 2446 6776 2994
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 6840 2106 6868 3012
rect 6920 2994 6972 3000
rect 6828 2100 6880 2106
rect 6828 2042 6880 2048
rect 6552 1760 6604 1766
rect 6552 1702 6604 1708
rect 6564 1494 6592 1702
rect 6552 1488 6604 1494
rect 6552 1430 6604 1436
rect 6840 1426 6868 2042
rect 7024 2038 7052 10610
rect 7116 9994 7144 10950
rect 7286 10906 7342 11942
rect 7286 10854 7288 10906
rect 7340 10854 7342 10906
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 7116 8974 7144 9930
rect 7208 9926 7236 10542
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7286 9818 7342 10854
rect 7392 10062 7420 12310
rect 7484 12238 7512 13466
rect 7576 13462 7604 15456
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7668 15026 7696 15302
rect 7656 15020 7708 15026
rect 7656 14962 7708 14968
rect 7748 14884 7800 14890
rect 7748 14826 7800 14832
rect 7760 14498 7788 14826
rect 7668 14470 7788 14498
rect 7668 14006 7696 14470
rect 7748 14340 7800 14346
rect 7748 14282 7800 14288
rect 7656 14000 7708 14006
rect 7656 13942 7708 13948
rect 7656 13796 7708 13802
rect 7656 13738 7708 13744
rect 7564 13456 7616 13462
rect 7564 13398 7616 13404
rect 7576 12986 7604 13398
rect 7668 13190 7696 13738
rect 7760 13530 7788 14282
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 7656 13184 7708 13190
rect 7708 13144 7788 13172
rect 7656 13126 7708 13132
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7656 12640 7708 12646
rect 7656 12582 7708 12588
rect 7668 12442 7696 12582
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7380 10056 7432 10062
rect 7380 9998 7432 10004
rect 7286 9766 7288 9818
rect 7340 9766 7342 9818
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 7116 7886 7144 8910
rect 7286 8730 7342 9766
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7286 8678 7288 8730
rect 7340 8678 7342 8730
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 7116 5030 7144 7822
rect 7286 7642 7342 8678
rect 7392 7954 7420 9454
rect 7484 8838 7512 12038
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 7576 9518 7604 11698
rect 7668 11218 7696 12038
rect 7656 11212 7708 11218
rect 7656 11154 7708 11160
rect 7656 10668 7708 10674
rect 7760 10656 7788 13144
rect 7852 12850 7880 16050
rect 7932 14272 7984 14278
rect 7932 14214 7984 14220
rect 7944 14074 7972 14214
rect 7932 14068 7984 14074
rect 7932 14010 7984 14016
rect 8036 13954 8064 17002
rect 8128 14600 8156 18550
rect 8220 17814 8248 19366
rect 8404 19334 8432 19858
rect 8496 19394 8524 20198
rect 8588 19718 8616 20742
rect 8864 20058 8892 30670
rect 8944 30660 8996 30666
rect 8944 30602 8996 30608
rect 8956 28762 8984 30602
rect 8944 28756 8996 28762
rect 8944 28698 8996 28704
rect 8944 27328 8996 27334
rect 8944 27270 8996 27276
rect 8956 27062 8984 27270
rect 8944 27056 8996 27062
rect 8944 26998 8996 27004
rect 8944 24200 8996 24206
rect 8944 24142 8996 24148
rect 8956 23866 8984 24142
rect 8944 23860 8996 23866
rect 8944 23802 8996 23808
rect 9048 22098 9076 31622
rect 9416 30938 9444 31690
rect 9876 31482 9904 32778
rect 9864 31476 9916 31482
rect 9864 31418 9916 31424
rect 9588 31408 9640 31414
rect 9588 31350 9640 31356
rect 9404 30932 9456 30938
rect 9404 30874 9456 30880
rect 9600 30258 9628 31350
rect 9772 30728 9824 30734
rect 9772 30670 9824 30676
rect 9864 30728 9916 30734
rect 9864 30670 9916 30676
rect 9680 30388 9732 30394
rect 9680 30330 9732 30336
rect 9496 30252 9548 30258
rect 9496 30194 9548 30200
rect 9588 30252 9640 30258
rect 9588 30194 9640 30200
rect 9508 30122 9536 30194
rect 9496 30116 9548 30122
rect 9496 30058 9548 30064
rect 9220 29606 9272 29612
rect 9272 29566 9444 29594
rect 9220 29548 9272 29554
rect 9220 29504 9272 29510
rect 9220 29446 9272 29452
rect 9232 29306 9260 29446
rect 9220 29300 9272 29306
rect 9220 29242 9272 29248
rect 9128 28960 9180 28966
rect 9128 28902 9180 28908
rect 9140 27674 9168 28902
rect 9416 28558 9444 29566
rect 9496 29504 9548 29510
rect 9496 29446 9548 29452
rect 9508 28966 9536 29446
rect 9496 28960 9548 28966
rect 9496 28902 9548 28908
rect 9588 28688 9640 28694
rect 9588 28630 9640 28636
rect 9220 28552 9272 28558
rect 9220 28494 9272 28500
rect 9404 28552 9456 28558
rect 9404 28494 9456 28500
rect 9128 27668 9180 27674
rect 9128 27610 9180 27616
rect 9140 25242 9168 27610
rect 9232 27538 9260 28494
rect 9496 28416 9548 28422
rect 9496 28358 9548 28364
rect 9220 27532 9272 27538
rect 9220 27474 9272 27480
rect 9232 26858 9260 27474
rect 9508 27470 9536 28358
rect 9496 27464 9548 27470
rect 9496 27406 9548 27412
rect 9496 27328 9548 27334
rect 9496 27270 9548 27276
rect 9508 27130 9536 27270
rect 9496 27124 9548 27130
rect 9496 27066 9548 27072
rect 9220 26852 9272 26858
rect 9220 26794 9272 26800
rect 9404 26036 9456 26042
rect 9404 25978 9456 25984
rect 9312 25900 9364 25906
rect 9312 25842 9364 25848
rect 9324 25702 9352 25842
rect 9220 25696 9272 25702
rect 9220 25638 9272 25644
rect 9312 25696 9364 25702
rect 9312 25638 9364 25644
rect 9232 25362 9260 25638
rect 9416 25430 9444 25978
rect 9600 25974 9628 28630
rect 9692 28558 9720 30330
rect 9784 29238 9812 30670
rect 9876 30190 9904 30670
rect 9864 30184 9916 30190
rect 9864 30126 9916 30132
rect 9876 29510 9904 30126
rect 9864 29504 9916 29510
rect 9864 29446 9916 29452
rect 9772 29232 9824 29238
rect 9772 29174 9824 29180
rect 9784 28694 9812 29174
rect 9772 28688 9824 28694
rect 9772 28630 9824 28636
rect 9680 28552 9732 28558
rect 9732 28512 9812 28540
rect 9680 28494 9732 28500
rect 9680 28416 9732 28422
rect 9680 28358 9732 28364
rect 9692 28218 9720 28358
rect 9680 28212 9732 28218
rect 9680 28154 9732 28160
rect 9784 28082 9812 28512
rect 9772 28076 9824 28082
rect 9772 28018 9824 28024
rect 9784 27946 9812 28018
rect 9772 27940 9824 27946
rect 9772 27882 9824 27888
rect 9772 26852 9824 26858
rect 9772 26794 9824 26800
rect 9784 26314 9812 26794
rect 9772 26308 9824 26314
rect 9772 26250 9824 26256
rect 9680 26240 9732 26246
rect 9680 26182 9732 26188
rect 9588 25968 9640 25974
rect 9588 25910 9640 25916
rect 9404 25424 9456 25430
rect 9404 25366 9456 25372
rect 9220 25356 9272 25362
rect 9220 25298 9272 25304
rect 9692 25294 9720 26182
rect 9772 25356 9824 25362
rect 9772 25298 9824 25304
rect 9312 25288 9364 25294
rect 9140 25214 9260 25242
rect 9312 25230 9364 25236
rect 9404 25288 9456 25294
rect 9404 25230 9456 25236
rect 9680 25288 9732 25294
rect 9680 25230 9732 25236
rect 9128 24812 9180 24818
rect 9128 24754 9180 24760
rect 9140 24614 9168 24754
rect 9128 24608 9180 24614
rect 9128 24550 9180 24556
rect 9140 24206 9168 24550
rect 9128 24200 9180 24206
rect 9128 24142 9180 24148
rect 9128 22976 9180 22982
rect 9128 22918 9180 22924
rect 9140 22710 9168 22918
rect 9128 22704 9180 22710
rect 9128 22646 9180 22652
rect 9036 22092 9088 22098
rect 9232 22094 9260 25214
rect 9324 24682 9352 25230
rect 9416 24954 9444 25230
rect 9404 24948 9456 24954
rect 9404 24890 9456 24896
rect 9588 24880 9640 24886
rect 9588 24822 9640 24828
rect 9404 24812 9456 24818
rect 9404 24754 9456 24760
rect 9312 24676 9364 24682
rect 9312 24618 9364 24624
rect 9416 24410 9444 24754
rect 9600 24410 9628 24822
rect 9404 24404 9456 24410
rect 9404 24346 9456 24352
rect 9588 24404 9640 24410
rect 9588 24346 9640 24352
rect 9680 24200 9732 24206
rect 9680 24142 9732 24148
rect 9588 23860 9640 23866
rect 9588 23802 9640 23808
rect 9600 23118 9628 23802
rect 9692 23798 9720 24142
rect 9784 24052 9812 25298
rect 9864 24064 9916 24070
rect 9784 24024 9864 24052
rect 9864 24006 9916 24012
rect 9680 23792 9732 23798
rect 9680 23734 9732 23740
rect 9876 23730 9904 24006
rect 9864 23724 9916 23730
rect 9784 23684 9864 23712
rect 9312 23112 9364 23118
rect 9312 23054 9364 23060
rect 9588 23112 9640 23118
rect 9588 23054 9640 23060
rect 9324 22778 9352 23054
rect 9312 22772 9364 22778
rect 9312 22714 9364 22720
rect 9784 22642 9812 23684
rect 9864 23666 9916 23672
rect 9968 22794 9996 33390
rect 10232 33380 10284 33386
rect 10232 33322 10284 33328
rect 10140 33312 10192 33318
rect 10140 33254 10192 33260
rect 10048 31340 10100 31346
rect 10048 31282 10100 31288
rect 10060 28762 10088 31282
rect 10048 28756 10100 28762
rect 10048 28698 10100 28704
rect 10152 22930 10180 33254
rect 10244 32910 10272 33322
rect 10232 32904 10284 32910
rect 10232 32846 10284 32852
rect 10232 29640 10284 29646
rect 10232 29582 10284 29588
rect 10244 29306 10272 29582
rect 10232 29300 10284 29306
rect 10232 29242 10284 29248
rect 10244 28082 10272 29242
rect 10232 28076 10284 28082
rect 10232 28018 10284 28024
rect 10244 27538 10272 28018
rect 10232 27532 10284 27538
rect 10232 27474 10284 27480
rect 10336 27130 10364 35974
rect 10428 34746 10456 40054
rect 10612 38282 10640 40326
rect 10796 39846 10824 40870
rect 11072 40458 11100 41006
rect 11428 40520 11480 40526
rect 11428 40462 11480 40468
rect 11060 40452 11112 40458
rect 11060 40394 11112 40400
rect 10876 40384 10928 40390
rect 10876 40326 10928 40332
rect 10888 40050 10916 40326
rect 11440 40050 11468 40462
rect 11532 40186 11560 41074
rect 11900 40730 11928 41210
rect 11888 40724 11940 40730
rect 11888 40666 11940 40672
rect 11796 40520 11848 40526
rect 11796 40462 11848 40468
rect 11612 40452 11664 40458
rect 11612 40394 11664 40400
rect 11520 40180 11572 40186
rect 11520 40122 11572 40128
rect 10876 40044 10928 40050
rect 10876 39986 10928 39992
rect 11428 40044 11480 40050
rect 11428 39986 11480 39992
rect 10784 39840 10836 39846
rect 10784 39782 10836 39788
rect 10796 39438 10824 39782
rect 10784 39432 10836 39438
rect 10784 39374 10836 39380
rect 10796 39098 10824 39374
rect 10784 39092 10836 39098
rect 10784 39034 10836 39040
rect 10600 38276 10652 38282
rect 10600 38218 10652 38224
rect 10508 36032 10560 36038
rect 10508 35974 10560 35980
rect 10520 35018 10548 35974
rect 10612 35834 10640 38218
rect 10692 37256 10744 37262
rect 10692 37198 10744 37204
rect 10704 36378 10732 37198
rect 10796 36378 10824 39034
rect 10968 38956 11020 38962
rect 10968 38898 11020 38904
rect 10980 38010 11008 38898
rect 11520 38752 11572 38758
rect 11520 38694 11572 38700
rect 10968 38004 11020 38010
rect 10968 37946 11020 37952
rect 10692 36372 10744 36378
rect 10692 36314 10744 36320
rect 10784 36372 10836 36378
rect 10784 36314 10836 36320
rect 10980 36242 11008 37946
rect 11532 37194 11560 38694
rect 11520 37188 11572 37194
rect 11520 37130 11572 37136
rect 11244 37120 11296 37126
rect 11244 37062 11296 37068
rect 11060 36780 11112 36786
rect 11060 36722 11112 36728
rect 11072 36378 11100 36722
rect 11060 36372 11112 36378
rect 11060 36314 11112 36320
rect 10968 36236 11020 36242
rect 10968 36178 11020 36184
rect 10692 36168 10744 36174
rect 10692 36110 10744 36116
rect 10600 35828 10652 35834
rect 10600 35770 10652 35776
rect 10508 35012 10560 35018
rect 10508 34954 10560 34960
rect 10416 34740 10468 34746
rect 10416 34682 10468 34688
rect 10416 34400 10468 34406
rect 10416 34342 10468 34348
rect 10428 33590 10456 34342
rect 10416 33584 10468 33590
rect 10416 33526 10468 33532
rect 10428 32978 10456 33526
rect 10416 32972 10468 32978
rect 10416 32914 10468 32920
rect 10428 32280 10456 32914
rect 10508 32292 10560 32298
rect 10428 32252 10508 32280
rect 10428 31804 10456 32252
rect 10508 32234 10560 32240
rect 10508 31816 10560 31822
rect 10428 31776 10508 31804
rect 10508 31758 10560 31764
rect 10612 31210 10640 35770
rect 10704 34202 10732 36110
rect 10876 35692 10928 35698
rect 10876 35634 10928 35640
rect 10784 35012 10836 35018
rect 10784 34954 10836 34960
rect 10796 34746 10824 34954
rect 10784 34740 10836 34746
rect 10784 34682 10836 34688
rect 10692 34196 10744 34202
rect 10692 34138 10744 34144
rect 10692 33516 10744 33522
rect 10692 33458 10744 33464
rect 10600 31204 10652 31210
rect 10600 31146 10652 31152
rect 10416 31136 10468 31142
rect 10416 31078 10468 31084
rect 10508 31136 10560 31142
rect 10508 31078 10560 31084
rect 10428 30734 10456 31078
rect 10416 30728 10468 30734
rect 10416 30670 10468 30676
rect 10520 30190 10548 31078
rect 10508 30184 10560 30190
rect 10508 30126 10560 30132
rect 10520 28966 10548 30126
rect 10600 29028 10652 29034
rect 10600 28970 10652 28976
rect 10508 28960 10560 28966
rect 10428 28920 10508 28948
rect 10428 27606 10456 28920
rect 10508 28902 10560 28908
rect 10508 28552 10560 28558
rect 10508 28494 10560 28500
rect 10520 28150 10548 28494
rect 10508 28144 10560 28150
rect 10508 28086 10560 28092
rect 10416 27600 10468 27606
rect 10416 27542 10468 27548
rect 10520 27470 10548 28086
rect 10508 27464 10560 27470
rect 10508 27406 10560 27412
rect 10324 27124 10376 27130
rect 10324 27066 10376 27072
rect 10612 26858 10640 28970
rect 10600 26852 10652 26858
rect 10600 26794 10652 26800
rect 10612 26024 10640 26794
rect 10520 25996 10640 26024
rect 10324 25832 10376 25838
rect 10324 25774 10376 25780
rect 10232 25696 10284 25702
rect 10232 25638 10284 25644
rect 10244 25158 10272 25638
rect 10232 25152 10284 25158
rect 10232 25094 10284 25100
rect 10336 24750 10364 25774
rect 10416 24880 10468 24886
rect 10416 24822 10468 24828
rect 10324 24744 10376 24750
rect 10324 24686 10376 24692
rect 10336 23730 10364 24686
rect 10324 23724 10376 23730
rect 10324 23666 10376 23672
rect 10232 23520 10284 23526
rect 10232 23462 10284 23468
rect 10244 23118 10272 23462
rect 10232 23112 10284 23118
rect 10232 23054 10284 23060
rect 10152 22902 10272 22930
rect 9876 22766 9996 22794
rect 10140 22772 10192 22778
rect 9772 22636 9824 22642
rect 9772 22578 9824 22584
rect 9680 22500 9732 22506
rect 9680 22442 9732 22448
rect 9692 22234 9720 22442
rect 9680 22228 9732 22234
rect 9680 22170 9732 22176
rect 9772 22228 9824 22234
rect 9772 22170 9824 22176
rect 9404 22160 9456 22166
rect 9784 22114 9812 22170
rect 9456 22108 9812 22114
rect 9404 22102 9812 22108
rect 9232 22066 9352 22094
rect 9416 22086 9812 22102
rect 9036 22034 9088 22040
rect 8944 22024 8996 22030
rect 8944 21966 8996 21972
rect 8760 20052 8812 20058
rect 8760 19994 8812 20000
rect 8852 20052 8904 20058
rect 8852 19994 8904 20000
rect 8668 19984 8720 19990
rect 8668 19926 8720 19932
rect 8576 19712 8628 19718
rect 8576 19654 8628 19660
rect 8496 19366 8616 19394
rect 8404 19306 8524 19334
rect 8208 17808 8260 17814
rect 8208 17750 8260 17756
rect 8392 17740 8444 17746
rect 8392 17682 8444 17688
rect 8208 17672 8260 17678
rect 8208 17614 8260 17620
rect 8220 17066 8248 17614
rect 8208 17060 8260 17066
rect 8208 17002 8260 17008
rect 8404 16998 8432 17682
rect 8496 17134 8524 19306
rect 8588 18986 8616 19366
rect 8680 19360 8708 19926
rect 8772 19514 8800 19994
rect 8760 19508 8812 19514
rect 8760 19450 8812 19456
rect 8956 19446 8984 21966
rect 9220 21548 9272 21554
rect 9220 21490 9272 21496
rect 9232 21146 9260 21490
rect 9220 21140 9272 21146
rect 9220 21082 9272 21088
rect 9220 20936 9272 20942
rect 9220 20878 9272 20884
rect 9036 20460 9088 20466
rect 9036 20402 9088 20408
rect 9128 20460 9180 20466
rect 9128 20402 9180 20408
rect 8944 19440 8996 19446
rect 8944 19382 8996 19388
rect 8760 19372 8812 19378
rect 8680 19332 8760 19360
rect 8760 19314 8812 19320
rect 8588 18958 8708 18986
rect 8576 18896 8628 18902
rect 8576 18838 8628 18844
rect 8484 17128 8536 17134
rect 8484 17070 8536 17076
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 8404 16658 8432 16934
rect 8392 16652 8444 16658
rect 8392 16594 8444 16600
rect 8208 16516 8260 16522
rect 8208 16458 8260 16464
rect 8220 16250 8248 16458
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 8496 15434 8524 17070
rect 8588 16590 8616 18838
rect 8680 18834 8708 18958
rect 8668 18828 8720 18834
rect 8668 18770 8720 18776
rect 8760 18760 8812 18766
rect 8760 18702 8812 18708
rect 8772 18358 8800 18702
rect 8760 18352 8812 18358
rect 8760 18294 8812 18300
rect 8956 17542 8984 19382
rect 9048 19174 9076 20402
rect 9140 19854 9168 20402
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 9036 19168 9088 19174
rect 9036 19110 9088 19116
rect 9036 18692 9088 18698
rect 9036 18634 9088 18640
rect 9048 18358 9076 18634
rect 9036 18352 9088 18358
rect 9036 18294 9088 18300
rect 9140 17954 9168 19790
rect 9232 19174 9260 20878
rect 9324 19990 9352 22066
rect 9588 21412 9640 21418
rect 9588 21354 9640 21360
rect 9404 21072 9456 21078
rect 9404 21014 9456 21020
rect 9416 20262 9444 21014
rect 9404 20256 9456 20262
rect 9404 20198 9456 20204
rect 9312 19984 9364 19990
rect 9312 19926 9364 19932
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 9232 18222 9260 19110
rect 9416 18834 9444 20198
rect 9404 18828 9456 18834
rect 9404 18770 9456 18776
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 9324 18290 9352 18702
rect 9312 18284 9364 18290
rect 9312 18226 9364 18232
rect 9600 18222 9628 21354
rect 9680 21072 9732 21078
rect 9680 21014 9732 21020
rect 9692 18766 9720 21014
rect 9772 20868 9824 20874
rect 9772 20810 9824 20816
rect 9784 20602 9812 20810
rect 9772 20596 9824 20602
rect 9772 20538 9824 20544
rect 9784 19786 9812 20538
rect 9772 19780 9824 19786
rect 9772 19722 9824 19728
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9220 18216 9272 18222
rect 9220 18158 9272 18164
rect 9588 18216 9640 18222
rect 9588 18158 9640 18164
rect 9220 18080 9272 18086
rect 9220 18022 9272 18028
rect 9048 17926 9168 17954
rect 8668 17536 8720 17542
rect 8668 17478 8720 17484
rect 8944 17536 8996 17542
rect 8944 17478 8996 17484
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 8680 16436 8708 17478
rect 8956 17202 8984 17478
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 8852 16788 8904 16794
rect 8852 16730 8904 16736
rect 8588 16408 8708 16436
rect 8588 15570 8616 16408
rect 8576 15564 8628 15570
rect 8576 15506 8628 15512
rect 8484 15428 8536 15434
rect 8484 15370 8536 15376
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8208 14612 8260 14618
rect 8128 14572 8208 14600
rect 8208 14554 8260 14560
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 8300 14272 8352 14278
rect 8300 14214 8352 14220
rect 7944 13926 8064 13954
rect 7840 12844 7892 12850
rect 7840 12786 7892 12792
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 7852 12102 7880 12174
rect 7840 12096 7892 12102
rect 7840 12038 7892 12044
rect 7944 11762 7972 13926
rect 8024 13796 8076 13802
rect 8024 13738 8076 13744
rect 8036 13462 8064 13738
rect 8024 13456 8076 13462
rect 8024 13398 8076 13404
rect 8220 12986 8248 14214
rect 8312 13870 8340 14214
rect 8404 13938 8432 14962
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 8208 12980 8260 12986
rect 8208 12922 8260 12928
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 7840 11688 7892 11694
rect 7840 11630 7892 11636
rect 7708 10628 7788 10656
rect 7656 10610 7708 10616
rect 7852 10554 7880 11630
rect 8220 11150 8248 12786
rect 8312 12782 8340 13806
rect 8496 13462 8524 15370
rect 8392 13456 8444 13462
rect 8392 13398 8444 13404
rect 8484 13456 8536 13462
rect 8484 13398 8536 13404
rect 8404 12850 8432 13398
rect 8588 13308 8616 15506
rect 8760 14476 8812 14482
rect 8760 14418 8812 14424
rect 8772 13870 8800 14418
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 8680 13530 8708 13670
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 8496 13280 8616 13308
rect 8392 12844 8444 12850
rect 8392 12786 8444 12792
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 7944 11014 7972 11086
rect 7932 11008 7984 11014
rect 7932 10950 7984 10956
rect 8024 11008 8076 11014
rect 8024 10950 8076 10956
rect 7923 10736 7975 10742
rect 8036 10724 8064 10950
rect 8312 10724 8340 11494
rect 7975 10696 8064 10724
rect 8266 10696 8340 10724
rect 7923 10678 7975 10684
rect 8116 10668 8168 10674
rect 8266 10656 8294 10696
rect 8168 10628 8294 10656
rect 8116 10610 8168 10616
rect 7668 10526 7880 10554
rect 7668 10198 7696 10526
rect 7748 10464 7800 10470
rect 7800 10424 8064 10452
rect 7748 10406 7800 10412
rect 8036 10248 8064 10424
rect 8208 10260 8260 10266
rect 8036 10220 8208 10248
rect 8208 10202 8260 10208
rect 7656 10192 7708 10198
rect 8496 10146 8524 13280
rect 8760 13252 8812 13258
rect 8760 13194 8812 13200
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8680 12442 8708 12922
rect 8772 12850 8800 13194
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 8588 10810 8616 12242
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 8576 10668 8628 10674
rect 8680 10656 8708 11698
rect 8628 10628 8708 10656
rect 8576 10610 8628 10616
rect 8680 10470 8708 10628
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 7656 10134 7708 10140
rect 7668 9722 7696 10134
rect 8036 10118 8524 10146
rect 8036 9874 8064 10118
rect 8392 9988 8444 9994
rect 8680 9976 8708 10406
rect 8772 9994 8800 12038
rect 8444 9948 8708 9976
rect 8760 9988 8812 9994
rect 8392 9930 8444 9936
rect 8760 9930 8812 9936
rect 8864 9926 8892 16730
rect 8956 16658 8984 17138
rect 8944 16652 8996 16658
rect 8944 16594 8996 16600
rect 8956 15570 8984 16594
rect 8944 15564 8996 15570
rect 8944 15506 8996 15512
rect 8956 15094 8984 15506
rect 8944 15088 8996 15094
rect 8944 15030 8996 15036
rect 8956 14482 8984 15030
rect 8944 14476 8996 14482
rect 8944 14418 8996 14424
rect 8956 12306 8984 14418
rect 8944 12300 8996 12306
rect 8944 12242 8996 12248
rect 9048 11642 9076 17926
rect 9232 17202 9260 18022
rect 9220 17196 9272 17202
rect 9496 17196 9548 17202
rect 9220 17138 9272 17144
rect 9416 17156 9496 17184
rect 9220 16516 9272 16522
rect 9220 16458 9272 16464
rect 9232 16250 9260 16458
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 9312 15428 9364 15434
rect 9312 15370 9364 15376
rect 9220 14952 9272 14958
rect 9220 14894 9272 14900
rect 9232 14770 9260 14894
rect 9140 14742 9260 14770
rect 9140 13938 9168 14742
rect 9128 13932 9180 13938
rect 9128 13874 9180 13880
rect 9140 12442 9168 13874
rect 9324 13802 9352 15370
rect 9416 14822 9444 17156
rect 9496 17138 9548 17144
rect 9692 16998 9720 18702
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9496 16448 9548 16454
rect 9496 16390 9548 16396
rect 9508 15910 9536 16390
rect 9692 16046 9720 16934
rect 9784 16454 9812 19722
rect 9772 16448 9824 16454
rect 9772 16390 9824 16396
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9496 15904 9548 15910
rect 9496 15846 9548 15852
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9496 14816 9548 14822
rect 9496 14758 9548 14764
rect 9404 14272 9456 14278
rect 9404 14214 9456 14220
rect 9312 13796 9364 13802
rect 9312 13738 9364 13744
rect 9416 13394 9444 14214
rect 9508 13938 9536 14758
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9588 14408 9640 14414
rect 9588 14350 9640 14356
rect 9600 14074 9628 14350
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 9784 12850 9812 14554
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 9128 12436 9180 12442
rect 9128 12378 9180 12384
rect 9232 12238 9260 12582
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9416 11762 9444 12038
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 9048 11614 9352 11642
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9036 11144 9088 11150
rect 9036 11086 9088 11092
rect 8944 11076 8996 11082
rect 8944 11018 8996 11024
rect 8956 10266 8984 11018
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 8944 9988 8996 9994
rect 8944 9930 8996 9936
rect 8300 9920 8352 9926
rect 8220 9880 8300 9908
rect 8220 9874 8248 9880
rect 7944 9846 8064 9874
rect 8216 9846 8248 9874
rect 8300 9862 8352 9868
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 7944 9738 7972 9846
rect 8216 9738 8244 9846
rect 8864 9738 8892 9862
rect 7656 9716 7708 9722
rect 7944 9710 8064 9738
rect 8216 9710 8432 9738
rect 7656 9658 7708 9664
rect 8036 9654 8064 9710
rect 8404 9654 8432 9710
rect 8496 9710 8892 9738
rect 8024 9648 8076 9654
rect 8024 9590 8076 9596
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7576 9178 7604 9454
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7564 9172 7616 9178
rect 7564 9114 7616 9120
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7668 8362 7696 9318
rect 8116 9036 8168 9042
rect 8116 8978 8168 8984
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 7656 8356 7708 8362
rect 7656 8298 7708 8304
rect 8036 8022 8064 8774
rect 8024 8016 8076 8022
rect 8024 7958 8076 7964
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 7286 7590 7288 7642
rect 7340 7590 7342 7642
rect 7196 7268 7248 7274
rect 7196 7210 7248 7216
rect 7104 5024 7156 5030
rect 7104 4966 7156 4972
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 7116 3398 7144 4014
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 7116 2854 7144 3334
rect 7104 2848 7156 2854
rect 7104 2790 7156 2796
rect 7012 2032 7064 2038
rect 7012 1974 7064 1980
rect 7208 1970 7236 7210
rect 7286 6554 7342 7590
rect 8128 7478 8156 8978
rect 8300 8900 8352 8906
rect 8300 8842 8352 8848
rect 8312 8634 8340 8842
rect 8496 8838 8524 9710
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8576 9376 8628 9382
rect 8576 9318 8628 9324
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8588 8634 8616 9318
rect 8680 8634 8708 9522
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 8220 8090 8248 8366
rect 8208 8084 8260 8090
rect 8208 8026 8260 8032
rect 8772 7546 8800 9454
rect 8956 8498 8984 9930
rect 9048 9722 9076 11086
rect 9140 11082 9168 11494
rect 9128 11076 9180 11082
rect 9128 11018 9180 11024
rect 9036 9716 9088 9722
rect 9036 9658 9088 9664
rect 9036 9444 9088 9450
rect 9036 9386 9088 9392
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8760 7540 8812 7546
rect 8760 7482 8812 7488
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 8128 7002 8156 7414
rect 8116 6996 8168 7002
rect 8116 6938 8168 6944
rect 8772 6866 8800 7482
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7286 6502 7288 6554
rect 7340 6502 7342 6554
rect 7286 5466 7342 6502
rect 7392 5642 7420 6598
rect 8956 6186 8984 8434
rect 9048 7818 9076 9386
rect 9140 9364 9168 11018
rect 9220 10124 9272 10130
rect 9220 10066 9272 10072
rect 9232 9722 9260 10066
rect 9220 9716 9272 9722
rect 9220 9658 9272 9664
rect 9324 9466 9352 11614
rect 9496 11280 9548 11286
rect 9496 11222 9548 11228
rect 9508 10674 9536 11222
rect 9692 11218 9720 12786
rect 9876 12434 9904 22766
rect 10060 22732 10140 22760
rect 9956 22636 10008 22642
rect 9956 22578 10008 22584
rect 9968 21554 9996 22578
rect 9956 21548 10008 21554
rect 9956 21490 10008 21496
rect 9956 20868 10008 20874
rect 9956 20810 10008 20816
rect 9968 20466 9996 20810
rect 10060 20806 10088 22732
rect 10140 22714 10192 22720
rect 10048 20800 10100 20806
rect 10048 20742 10100 20748
rect 9956 20460 10008 20466
rect 9956 20402 10008 20408
rect 9968 19854 9996 20402
rect 9956 19848 10008 19854
rect 9956 19790 10008 19796
rect 10140 19780 10192 19786
rect 10140 19722 10192 19728
rect 9956 19372 10008 19378
rect 9956 19314 10008 19320
rect 9968 18986 9996 19314
rect 9968 18958 10088 18986
rect 9956 18896 10008 18902
rect 9956 18838 10008 18844
rect 9968 14550 9996 18838
rect 10060 18222 10088 18958
rect 10152 18698 10180 19722
rect 10140 18692 10192 18698
rect 10140 18634 10192 18640
rect 10048 18216 10100 18222
rect 10048 18158 10100 18164
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 10060 17814 10088 18022
rect 10140 17876 10192 17882
rect 10140 17818 10192 17824
rect 10048 17808 10100 17814
rect 10048 17750 10100 17756
rect 10060 15978 10088 17750
rect 10048 15972 10100 15978
rect 10048 15914 10100 15920
rect 10048 15020 10100 15026
rect 10048 14962 10100 14968
rect 9956 14544 10008 14550
rect 9956 14486 10008 14492
rect 9968 13938 9996 14486
rect 10060 13938 10088 14962
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 9876 12406 10088 12434
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9588 10532 9640 10538
rect 9588 10474 9640 10480
rect 9600 9654 9628 10474
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 9692 9586 9720 10542
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9324 9438 9628 9466
rect 9496 9376 9548 9382
rect 9140 9336 9496 9364
rect 9496 9318 9548 9324
rect 9600 8974 9628 9438
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9692 9110 9720 9386
rect 9680 9104 9732 9110
rect 9680 9046 9732 9052
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9588 8968 9640 8974
rect 9588 8910 9640 8916
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 9140 7886 9168 8230
rect 9232 8090 9260 8910
rect 9680 8560 9732 8566
rect 9784 8548 9812 11698
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 9876 10674 9904 11086
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 9864 9988 9916 9994
rect 9968 9976 9996 11834
rect 9916 9948 9996 9976
rect 9864 9930 9916 9936
rect 9732 8520 9812 8548
rect 9864 8560 9916 8566
rect 9680 8502 9732 8508
rect 9864 8502 9916 8508
rect 9876 8412 9904 8502
rect 9416 8384 9904 8412
rect 9312 8356 9364 8362
rect 9416 8344 9444 8384
rect 9364 8316 9444 8344
rect 9312 8298 9364 8304
rect 9772 8288 9824 8294
rect 9772 8230 9824 8236
rect 9220 8084 9272 8090
rect 9220 8026 9272 8032
rect 9784 7954 9812 8230
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9036 7812 9088 7818
rect 9036 7754 9088 7760
rect 9404 7200 9456 7206
rect 9404 7142 9456 7148
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 8944 6180 8996 6186
rect 8944 6122 8996 6128
rect 7472 5772 7524 5778
rect 7472 5714 7524 5720
rect 7380 5636 7432 5642
rect 7380 5578 7432 5584
rect 7286 5414 7288 5466
rect 7340 5414 7342 5466
rect 7286 4378 7342 5414
rect 7286 4326 7288 4378
rect 7340 4326 7342 4378
rect 7286 3290 7342 4326
rect 7392 4146 7420 5578
rect 7484 4554 7512 5714
rect 8956 5710 8984 6122
rect 8944 5704 8996 5710
rect 8944 5646 8996 5652
rect 8668 5636 8720 5642
rect 8668 5578 8720 5584
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8496 5302 8524 5510
rect 7840 5296 7892 5302
rect 7840 5238 7892 5244
rect 8484 5296 8536 5302
rect 8484 5238 8536 5244
rect 7656 5092 7708 5098
rect 7656 5034 7708 5040
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7472 4548 7524 4554
rect 7472 4490 7524 4496
rect 7484 4282 7512 4490
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7380 4140 7432 4146
rect 7576 4128 7604 4762
rect 7668 4758 7696 5034
rect 7656 4752 7708 4758
rect 7656 4694 7708 4700
rect 7656 4140 7708 4146
rect 7576 4100 7656 4128
rect 7380 4082 7432 4088
rect 7656 4082 7708 4088
rect 7852 3466 7880 5238
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 7944 4826 7972 5170
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 8024 4752 8076 4758
rect 8024 4694 8076 4700
rect 7932 4004 7984 4010
rect 8036 3992 8064 4694
rect 8588 4146 8616 5170
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 7984 3964 8064 3992
rect 7932 3946 7984 3952
rect 7564 3460 7616 3466
rect 7564 3402 7616 3408
rect 7840 3460 7892 3466
rect 7840 3402 7892 3408
rect 7286 3238 7288 3290
rect 7340 3238 7342 3290
rect 7286 2202 7342 3238
rect 7576 2922 7604 3402
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7760 3126 7788 3334
rect 7748 3120 7800 3126
rect 7748 3062 7800 3068
rect 7564 2916 7616 2922
rect 7564 2858 7616 2864
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 7380 2304 7432 2310
rect 7380 2246 7432 2252
rect 7286 2150 7288 2202
rect 7340 2150 7342 2202
rect 7196 1964 7248 1970
rect 7196 1906 7248 1912
rect 6828 1420 6880 1426
rect 6828 1362 6880 1368
rect 6368 1352 6420 1358
rect 6368 1294 6420 1300
rect 7286 1114 7342 2150
rect 7392 1358 7420 2246
rect 7576 2106 7604 2382
rect 7564 2100 7616 2106
rect 7564 2042 7616 2048
rect 7472 1964 7524 1970
rect 7472 1906 7524 1912
rect 7484 1562 7512 1906
rect 7472 1556 7524 1562
rect 7472 1498 7524 1504
rect 7852 1358 7880 3402
rect 8680 3058 8708 5578
rect 9324 4690 9352 6258
rect 9416 5710 9444 7142
rect 9692 6322 9720 7822
rect 9784 6866 9812 7890
rect 10060 7546 10088 12406
rect 10152 11762 10180 17818
rect 10244 17066 10272 22902
rect 10336 22642 10364 23666
rect 10324 22636 10376 22642
rect 10324 22578 10376 22584
rect 10336 21554 10364 22578
rect 10324 21548 10376 21554
rect 10324 21490 10376 21496
rect 10428 20312 10456 24822
rect 10520 24750 10548 25996
rect 10600 25900 10652 25906
rect 10600 25842 10652 25848
rect 10612 25362 10640 25842
rect 10600 25356 10652 25362
rect 10600 25298 10652 25304
rect 10600 25152 10652 25158
rect 10600 25094 10652 25100
rect 10612 24954 10640 25094
rect 10600 24948 10652 24954
rect 10600 24890 10652 24896
rect 10508 24744 10560 24750
rect 10508 24686 10560 24692
rect 10508 24268 10560 24274
rect 10508 24210 10560 24216
rect 10520 23730 10548 24210
rect 10600 24200 10652 24206
rect 10600 24142 10652 24148
rect 10612 23866 10640 24142
rect 10600 23860 10652 23866
rect 10600 23802 10652 23808
rect 10508 23724 10560 23730
rect 10508 23666 10560 23672
rect 10508 22432 10560 22438
rect 10508 22374 10560 22380
rect 10520 21894 10548 22374
rect 10508 21888 10560 21894
rect 10508 21830 10560 21836
rect 10704 21536 10732 33458
rect 10784 33312 10836 33318
rect 10784 33254 10836 33260
rect 10796 24886 10824 33254
rect 10888 27010 10916 35634
rect 10980 35222 11008 36178
rect 11060 36100 11112 36106
rect 11060 36042 11112 36048
rect 11072 35698 11100 36042
rect 11060 35692 11112 35698
rect 11060 35634 11112 35640
rect 10968 35216 11020 35222
rect 10968 35158 11020 35164
rect 10980 34746 11008 35158
rect 11060 34944 11112 34950
rect 11060 34886 11112 34892
rect 10968 34740 11020 34746
rect 10968 34682 11020 34688
rect 11072 33998 11100 34886
rect 11060 33992 11112 33998
rect 11060 33934 11112 33940
rect 11072 31346 11100 33934
rect 11060 31340 11112 31346
rect 11060 31282 11112 31288
rect 11152 31272 11204 31278
rect 11152 31214 11204 31220
rect 10968 31136 11020 31142
rect 10968 31078 11020 31084
rect 10980 30938 11008 31078
rect 11164 30938 11192 31214
rect 10968 30932 11020 30938
rect 11152 30932 11204 30938
rect 10968 30874 11020 30880
rect 11072 30892 11152 30920
rect 10968 28688 11020 28694
rect 10968 28630 11020 28636
rect 11072 28642 11100 30892
rect 11152 30874 11204 30880
rect 11152 29164 11204 29170
rect 11152 29106 11204 29112
rect 11164 28762 11192 29106
rect 11152 28756 11204 28762
rect 11152 28698 11204 28704
rect 10980 28082 11008 28630
rect 11072 28626 11192 28642
rect 11072 28620 11204 28626
rect 11072 28614 11152 28620
rect 11152 28562 11204 28568
rect 11060 28416 11112 28422
rect 11060 28358 11112 28364
rect 11072 28218 11100 28358
rect 11060 28212 11112 28218
rect 11060 28154 11112 28160
rect 10968 28076 11020 28082
rect 10968 28018 11020 28024
rect 10888 26982 11008 27010
rect 10876 26920 10928 26926
rect 10876 26862 10928 26868
rect 10888 26246 10916 26862
rect 10876 26240 10928 26246
rect 10876 26182 10928 26188
rect 10888 25906 10916 26182
rect 10876 25900 10928 25906
rect 10876 25842 10928 25848
rect 10784 24880 10836 24886
rect 10784 24822 10836 24828
rect 10784 24064 10836 24070
rect 10784 24006 10836 24012
rect 10796 23254 10824 24006
rect 10784 23248 10836 23254
rect 10784 23190 10836 23196
rect 10888 23186 10916 25842
rect 10980 25242 11008 26982
rect 11072 26874 11100 28154
rect 11256 27130 11284 37062
rect 11624 36786 11652 40394
rect 11808 40050 11836 40462
rect 11796 40044 11848 40050
rect 11796 39986 11848 39992
rect 11808 38894 11836 39986
rect 11900 38962 11928 40666
rect 12268 40050 12296 41414
rect 12438 40826 12494 41862
rect 12728 41274 12756 42162
rect 12992 42152 13044 42158
rect 12992 42094 13044 42100
rect 16396 42152 16448 42158
rect 16396 42094 16448 42100
rect 17224 42152 17276 42158
rect 17224 42094 17276 42100
rect 12900 42016 12952 42022
rect 12900 41958 12952 41964
rect 12716 41268 12768 41274
rect 12716 41210 12768 41216
rect 12624 41132 12676 41138
rect 12624 41074 12676 41080
rect 12438 40774 12440 40826
rect 12492 40774 12494 40826
rect 12256 40044 12308 40050
rect 12256 39986 12308 39992
rect 12072 39568 12124 39574
rect 12072 39510 12124 39516
rect 11980 39296 12032 39302
rect 11980 39238 12032 39244
rect 11992 38962 12020 39238
rect 11888 38956 11940 38962
rect 11888 38898 11940 38904
rect 11980 38956 12032 38962
rect 11980 38898 12032 38904
rect 11796 38888 11848 38894
rect 11796 38830 11848 38836
rect 11900 38554 11928 38898
rect 12084 38554 12112 39510
rect 12268 39370 12296 39986
rect 12348 39976 12400 39982
rect 12348 39918 12400 39924
rect 12256 39364 12308 39370
rect 12256 39306 12308 39312
rect 12164 38752 12216 38758
rect 12164 38694 12216 38700
rect 11888 38548 11940 38554
rect 11888 38490 11940 38496
rect 12072 38548 12124 38554
rect 12072 38490 12124 38496
rect 11704 38480 11756 38486
rect 11704 38422 11756 38428
rect 11716 37398 11744 38422
rect 11796 38208 11848 38214
rect 11796 38150 11848 38156
rect 11808 37874 11836 38150
rect 11900 38010 11928 38490
rect 12072 38344 12124 38350
rect 12072 38286 12124 38292
rect 11888 38004 11940 38010
rect 11888 37946 11940 37952
rect 11796 37868 11848 37874
rect 11796 37810 11848 37816
rect 11704 37392 11756 37398
rect 11704 37334 11756 37340
rect 11900 37330 11928 37946
rect 12084 37942 12112 38286
rect 12072 37936 12124 37942
rect 12072 37878 12124 37884
rect 12072 37800 12124 37806
rect 12176 37788 12204 38694
rect 12124 37760 12204 37788
rect 12072 37742 12124 37748
rect 11980 37664 12032 37670
rect 11980 37606 12032 37612
rect 11888 37324 11940 37330
rect 11888 37266 11940 37272
rect 11612 36780 11664 36786
rect 11612 36722 11664 36728
rect 11796 36780 11848 36786
rect 11796 36722 11848 36728
rect 11704 36576 11756 36582
rect 11704 36518 11756 36524
rect 11612 36304 11664 36310
rect 11612 36246 11664 36252
rect 11428 36168 11480 36174
rect 11428 36110 11480 36116
rect 11440 31754 11468 36110
rect 11520 35828 11572 35834
rect 11520 35770 11572 35776
rect 11532 35630 11560 35770
rect 11624 35698 11652 36246
rect 11612 35692 11664 35698
rect 11612 35634 11664 35640
rect 11520 35624 11572 35630
rect 11520 35566 11572 35572
rect 11532 32502 11560 35566
rect 11716 34678 11744 36518
rect 11704 34672 11756 34678
rect 11704 34614 11756 34620
rect 11704 33924 11756 33930
rect 11704 33866 11756 33872
rect 11716 33658 11744 33866
rect 11704 33652 11756 33658
rect 11704 33594 11756 33600
rect 11704 33516 11756 33522
rect 11704 33458 11756 33464
rect 11612 33108 11664 33114
rect 11612 33050 11664 33056
rect 11624 32502 11652 33050
rect 11716 32842 11744 33458
rect 11704 32836 11756 32842
rect 11704 32778 11756 32784
rect 11520 32496 11572 32502
rect 11520 32438 11572 32444
rect 11612 32496 11664 32502
rect 11612 32438 11664 32444
rect 11716 32026 11744 32778
rect 11704 32020 11756 32026
rect 11704 31962 11756 31968
rect 11348 31726 11468 31754
rect 11244 27124 11296 27130
rect 11244 27066 11296 27072
rect 11072 26846 11192 26874
rect 11060 26784 11112 26790
rect 11060 26726 11112 26732
rect 11072 25974 11100 26726
rect 11060 25968 11112 25974
rect 11060 25910 11112 25916
rect 11072 25770 11100 25910
rect 11060 25764 11112 25770
rect 11060 25706 11112 25712
rect 10980 25214 11100 25242
rect 10968 25152 11020 25158
rect 10968 25094 11020 25100
rect 10980 24206 11008 25094
rect 10968 24200 11020 24206
rect 10968 24142 11020 24148
rect 11072 23866 11100 25214
rect 11060 23860 11112 23866
rect 11060 23802 11112 23808
rect 11164 23746 11192 26846
rect 11244 26852 11296 26858
rect 11244 26794 11296 26800
rect 11256 24188 11284 26794
rect 11348 25226 11376 31726
rect 11428 31680 11480 31686
rect 11428 31622 11480 31628
rect 11440 26994 11468 31622
rect 11704 31408 11756 31414
rect 11704 31350 11756 31356
rect 11716 30938 11744 31350
rect 11808 31278 11836 36722
rect 11900 35154 11928 37266
rect 11992 37194 12020 37606
rect 12072 37256 12124 37262
rect 12072 37198 12124 37204
rect 11980 37188 12032 37194
rect 11980 37130 12032 37136
rect 12084 36038 12112 37198
rect 12268 36922 12296 39306
rect 12360 37466 12388 39918
rect 12438 39738 12494 40774
rect 12636 40050 12664 41074
rect 12808 40384 12860 40390
rect 12808 40326 12860 40332
rect 12820 40050 12848 40326
rect 12624 40044 12676 40050
rect 12624 39986 12676 39992
rect 12808 40044 12860 40050
rect 12808 39986 12860 39992
rect 12532 39908 12584 39914
rect 12532 39850 12584 39856
rect 12438 39686 12440 39738
rect 12492 39686 12494 39738
rect 12438 38650 12494 39686
rect 12544 39030 12572 39850
rect 12912 39846 12940 41958
rect 13004 40934 13032 42094
rect 16028 42084 16080 42090
rect 16028 42026 16080 42032
rect 14004 41608 14056 41614
rect 14004 41550 14056 41556
rect 13084 41132 13136 41138
rect 13084 41074 13136 41080
rect 12992 40928 13044 40934
rect 12992 40870 13044 40876
rect 13096 40526 13124 41074
rect 13452 40928 13504 40934
rect 13452 40870 13504 40876
rect 13464 40526 13492 40870
rect 14016 40526 14044 41550
rect 15108 41540 15160 41546
rect 15108 41482 15160 41488
rect 14280 41472 14332 41478
rect 14280 41414 14332 41420
rect 14108 41386 14320 41414
rect 14108 41138 14136 41386
rect 15120 41274 15148 41482
rect 15752 41472 15804 41478
rect 15752 41414 15804 41420
rect 15108 41268 15160 41274
rect 15108 41210 15160 41216
rect 15764 41138 15792 41414
rect 14096 41132 14148 41138
rect 14096 41074 14148 41080
rect 14740 41132 14792 41138
rect 14740 41074 14792 41080
rect 15752 41132 15804 41138
rect 15752 41074 15804 41080
rect 14108 41002 14136 41074
rect 14648 41064 14700 41070
rect 14648 41006 14700 41012
rect 14096 40996 14148 41002
rect 14096 40938 14148 40944
rect 13084 40520 13136 40526
rect 13084 40462 13136 40468
rect 13452 40520 13504 40526
rect 13452 40462 13504 40468
rect 14004 40520 14056 40526
rect 14004 40462 14056 40468
rect 12624 39840 12676 39846
rect 12624 39782 12676 39788
rect 12900 39840 12952 39846
rect 12900 39782 12952 39788
rect 12636 39642 12664 39782
rect 12624 39636 12676 39642
rect 12624 39578 12676 39584
rect 12532 39024 12584 39030
rect 12532 38966 12584 38972
rect 12438 38598 12440 38650
rect 12492 38598 12494 38650
rect 12438 37562 12494 38598
rect 12544 38350 12572 38966
rect 12532 38344 12584 38350
rect 12532 38286 12584 38292
rect 12438 37510 12440 37562
rect 12492 37510 12494 37562
rect 12348 37460 12400 37466
rect 12348 37402 12400 37408
rect 12256 36916 12308 36922
rect 12256 36858 12308 36864
rect 12438 36474 12494 37510
rect 12544 36786 12572 38286
rect 12636 37738 12664 39578
rect 13096 39438 13124 40462
rect 13084 39432 13136 39438
rect 13084 39374 13136 39380
rect 13360 39296 13412 39302
rect 13360 39238 13412 39244
rect 13372 38350 13400 39238
rect 13084 38344 13136 38350
rect 13084 38286 13136 38292
rect 13360 38344 13412 38350
rect 13360 38286 13412 38292
rect 12624 37732 12676 37738
rect 12716 37732 12768 37738
rect 12676 37692 12716 37720
rect 12624 37674 12676 37680
rect 12716 37674 12768 37680
rect 13096 37466 13124 38286
rect 13268 37664 13320 37670
rect 13268 37606 13320 37612
rect 13084 37460 13136 37466
rect 13084 37402 13136 37408
rect 13096 36786 13124 37402
rect 13280 36786 13308 37606
rect 13372 37398 13400 38286
rect 13360 37392 13412 37398
rect 13360 37334 13412 37340
rect 13464 36786 13492 40462
rect 13820 39976 13872 39982
rect 13820 39918 13872 39924
rect 13832 39438 13860 39918
rect 13820 39432 13872 39438
rect 13820 39374 13872 39380
rect 13832 38758 13860 39374
rect 14016 38894 14044 40462
rect 14004 38888 14056 38894
rect 14004 38830 14056 38836
rect 13820 38752 13872 38758
rect 13820 38694 13872 38700
rect 14016 38486 14044 38830
rect 14004 38480 14056 38486
rect 14004 38422 14056 38428
rect 13820 38208 13872 38214
rect 13820 38150 13872 38156
rect 13636 37868 13688 37874
rect 13636 37810 13688 37816
rect 13648 37466 13676 37810
rect 13728 37800 13780 37806
rect 13728 37742 13780 37748
rect 13636 37460 13688 37466
rect 13636 37402 13688 37408
rect 12532 36780 12584 36786
rect 12532 36722 12584 36728
rect 13084 36780 13136 36786
rect 13084 36722 13136 36728
rect 13268 36780 13320 36786
rect 13268 36722 13320 36728
rect 13452 36780 13504 36786
rect 13452 36722 13504 36728
rect 12438 36422 12440 36474
rect 12492 36422 12494 36474
rect 12072 36032 12124 36038
rect 12072 35974 12124 35980
rect 12438 35386 12494 36422
rect 12900 35488 12952 35494
rect 12900 35430 12952 35436
rect 12438 35334 12440 35386
rect 12492 35334 12494 35386
rect 11888 35148 11940 35154
rect 11888 35090 11940 35096
rect 12256 34944 12308 34950
rect 12256 34886 12308 34892
rect 11888 34740 11940 34746
rect 11888 34682 11940 34688
rect 11900 33998 11928 34682
rect 12268 34678 12296 34886
rect 12256 34672 12308 34678
rect 12256 34614 12308 34620
rect 12348 34536 12400 34542
rect 12348 34478 12400 34484
rect 11888 33992 11940 33998
rect 11888 33934 11940 33940
rect 11980 33992 12032 33998
rect 11980 33934 12032 33940
rect 11992 33522 12020 33934
rect 12164 33856 12216 33862
rect 12164 33798 12216 33804
rect 11980 33516 12032 33522
rect 11980 33458 12032 33464
rect 11888 32972 11940 32978
rect 11888 32914 11940 32920
rect 11900 32842 11928 32914
rect 11888 32836 11940 32842
rect 11888 32778 11940 32784
rect 12072 32224 12124 32230
rect 12072 32166 12124 32172
rect 11980 32020 12032 32026
rect 11980 31962 12032 31968
rect 11888 31748 11940 31754
rect 11888 31690 11940 31696
rect 11900 31482 11928 31690
rect 11888 31476 11940 31482
rect 11888 31418 11940 31424
rect 11992 31414 12020 31962
rect 12084 31822 12112 32166
rect 12176 31890 12204 33798
rect 12256 32768 12308 32774
rect 12256 32710 12308 32716
rect 12268 32570 12296 32710
rect 12256 32564 12308 32570
rect 12256 32506 12308 32512
rect 12256 32428 12308 32434
rect 12256 32370 12308 32376
rect 12164 31884 12216 31890
rect 12164 31826 12216 31832
rect 12072 31816 12124 31822
rect 12072 31758 12124 31764
rect 12268 31754 12296 32370
rect 12176 31726 12296 31754
rect 11980 31408 12032 31414
rect 11980 31350 12032 31356
rect 11796 31272 11848 31278
rect 11796 31214 11848 31220
rect 11888 31204 11940 31210
rect 11888 31146 11940 31152
rect 11704 30932 11756 30938
rect 11624 30892 11704 30920
rect 11520 29572 11572 29578
rect 11520 29514 11572 29520
rect 11532 29306 11560 29514
rect 11520 29300 11572 29306
rect 11520 29242 11572 29248
rect 11520 28960 11572 28966
rect 11520 28902 11572 28908
rect 11532 28762 11560 28902
rect 11520 28756 11572 28762
rect 11520 28698 11572 28704
rect 11624 28218 11652 30892
rect 11704 30874 11756 30880
rect 11704 30048 11756 30054
rect 11704 29990 11756 29996
rect 11716 28422 11744 29990
rect 11900 29782 11928 31146
rect 12176 30734 12204 31726
rect 12256 31136 12308 31142
rect 12256 31078 12308 31084
rect 12164 30728 12216 30734
rect 12164 30670 12216 30676
rect 12072 30592 12124 30598
rect 12072 30534 12124 30540
rect 12084 30190 12112 30534
rect 11980 30184 12032 30190
rect 11980 30126 12032 30132
rect 12072 30184 12124 30190
rect 12072 30126 12124 30132
rect 11888 29776 11940 29782
rect 11888 29718 11940 29724
rect 11900 28490 11928 29718
rect 11992 28558 12020 30126
rect 12072 29164 12124 29170
rect 12072 29106 12124 29112
rect 12084 28762 12112 29106
rect 12072 28756 12124 28762
rect 12072 28698 12124 28704
rect 11980 28552 12032 28558
rect 11980 28494 12032 28500
rect 12072 28552 12124 28558
rect 12072 28494 12124 28500
rect 11888 28484 11940 28490
rect 11888 28426 11940 28432
rect 11704 28416 11756 28422
rect 11704 28358 11756 28364
rect 11612 28212 11664 28218
rect 11612 28154 11664 28160
rect 11612 28076 11664 28082
rect 11612 28018 11664 28024
rect 11520 28008 11572 28014
rect 11520 27950 11572 27956
rect 11428 26988 11480 26994
rect 11428 26930 11480 26936
rect 11532 26382 11560 27950
rect 11624 27674 11652 28018
rect 11612 27668 11664 27674
rect 11612 27610 11664 27616
rect 11796 27668 11848 27674
rect 11796 27610 11848 27616
rect 11808 27316 11836 27610
rect 11900 27470 11928 28426
rect 11980 28212 12032 28218
rect 11980 28154 12032 28160
rect 11888 27464 11940 27470
rect 11888 27406 11940 27412
rect 11808 27288 11928 27316
rect 11612 27124 11664 27130
rect 11612 27066 11664 27072
rect 11624 26586 11652 27066
rect 11704 26988 11756 26994
rect 11900 26978 11928 27288
rect 11704 26930 11756 26936
rect 11888 26972 11940 26978
rect 11612 26580 11664 26586
rect 11612 26522 11664 26528
rect 11520 26376 11572 26382
rect 11520 26318 11572 26324
rect 11532 25906 11560 26318
rect 11716 26246 11744 26930
rect 11888 26914 11940 26920
rect 11888 26852 11940 26858
rect 11888 26794 11940 26800
rect 11796 26512 11848 26518
rect 11796 26454 11848 26460
rect 11808 26382 11836 26454
rect 11900 26382 11928 26794
rect 11796 26376 11848 26382
rect 11796 26318 11848 26324
rect 11888 26376 11940 26382
rect 11888 26318 11940 26324
rect 11612 26240 11664 26246
rect 11612 26182 11664 26188
rect 11704 26240 11756 26246
rect 11704 26182 11756 26188
rect 11624 25906 11652 26182
rect 11520 25900 11572 25906
rect 11520 25842 11572 25848
rect 11612 25900 11664 25906
rect 11612 25842 11664 25848
rect 11428 25288 11480 25294
rect 11428 25230 11480 25236
rect 11336 25220 11388 25226
rect 11336 25162 11388 25168
rect 11440 24410 11468 25230
rect 11532 24886 11560 25842
rect 11716 25498 11744 26182
rect 11992 25650 12020 28154
rect 12084 27470 12112 28494
rect 12176 28422 12204 30670
rect 12268 30326 12296 31078
rect 12256 30320 12308 30326
rect 12256 30262 12308 30268
rect 12256 29504 12308 29510
rect 12256 29446 12308 29452
rect 12164 28416 12216 28422
rect 12164 28358 12216 28364
rect 12268 28234 12296 29446
rect 12360 28762 12388 34478
rect 12438 34298 12494 35334
rect 12912 35290 12940 35430
rect 12900 35284 12952 35290
rect 12900 35226 12952 35232
rect 13096 34950 13124 36722
rect 13280 36310 13308 36722
rect 13544 36576 13596 36582
rect 13544 36518 13596 36524
rect 13268 36304 13320 36310
rect 13268 36246 13320 36252
rect 13176 36168 13228 36174
rect 13176 36110 13228 36116
rect 13084 34944 13136 34950
rect 13084 34886 13136 34892
rect 12438 34246 12440 34298
rect 12492 34246 12494 34298
rect 12438 33210 12494 34246
rect 12992 33992 13044 33998
rect 12992 33934 13044 33940
rect 12532 33312 12584 33318
rect 12532 33254 12584 33260
rect 12438 33158 12440 33210
rect 12492 33158 12494 33210
rect 12438 32122 12494 33158
rect 12438 32070 12440 32122
rect 12492 32070 12494 32122
rect 12438 31034 12494 32070
rect 12544 31142 12572 33254
rect 12624 32904 12676 32910
rect 12624 32846 12676 32852
rect 12636 32366 12664 32846
rect 12716 32496 12768 32502
rect 12716 32438 12768 32444
rect 12624 32360 12676 32366
rect 12624 32302 12676 32308
rect 12728 31958 12756 32438
rect 12900 32224 12952 32230
rect 12900 32166 12952 32172
rect 12716 31952 12768 31958
rect 12716 31894 12768 31900
rect 12808 31952 12860 31958
rect 12808 31894 12860 31900
rect 12716 31816 12768 31822
rect 12716 31758 12768 31764
rect 12532 31136 12584 31142
rect 12532 31078 12584 31084
rect 12438 30982 12440 31034
rect 12492 30982 12494 31034
rect 12438 29946 12494 30982
rect 12728 30938 12756 31758
rect 12820 31278 12848 31894
rect 12808 31272 12860 31278
rect 12808 31214 12860 31220
rect 12716 30932 12768 30938
rect 12716 30874 12768 30880
rect 12532 30660 12584 30666
rect 12532 30602 12584 30608
rect 12624 30660 12676 30666
rect 12624 30602 12676 30608
rect 12544 30394 12572 30602
rect 12532 30388 12584 30394
rect 12532 30330 12584 30336
rect 12532 30252 12584 30258
rect 12636 30240 12664 30602
rect 12912 30394 12940 32166
rect 12808 30388 12860 30394
rect 12808 30330 12860 30336
rect 12900 30388 12952 30394
rect 12900 30330 12952 30336
rect 12584 30212 12664 30240
rect 12532 30194 12584 30200
rect 12438 29894 12440 29946
rect 12492 29894 12494 29946
rect 12438 28858 12494 29894
rect 12544 29102 12572 30194
rect 12820 29322 12848 30330
rect 12912 30002 12940 30330
rect 13004 30258 13032 33934
rect 13188 33454 13216 36110
rect 13360 36100 13412 36106
rect 13360 36042 13412 36048
rect 13372 35766 13400 36042
rect 13360 35760 13412 35766
rect 13360 35702 13412 35708
rect 13452 35760 13504 35766
rect 13452 35702 13504 35708
rect 13464 35578 13492 35702
rect 13556 35698 13584 36518
rect 13740 35698 13768 37742
rect 13832 37194 13860 38150
rect 13820 37188 13872 37194
rect 13820 37130 13872 37136
rect 14016 36174 14044 38422
rect 14108 37890 14136 40938
rect 14660 40458 14688 41006
rect 14648 40452 14700 40458
rect 14648 40394 14700 40400
rect 14660 40050 14688 40394
rect 14648 40044 14700 40050
rect 14648 39986 14700 39992
rect 14660 39506 14688 39986
rect 14752 39914 14780 41074
rect 15660 40928 15712 40934
rect 15660 40870 15712 40876
rect 15292 40452 15344 40458
rect 15292 40394 15344 40400
rect 15304 40050 15332 40394
rect 15476 40384 15528 40390
rect 15476 40326 15528 40332
rect 15384 40112 15436 40118
rect 15384 40054 15436 40060
rect 15292 40044 15344 40050
rect 15292 39986 15344 39992
rect 15200 39976 15252 39982
rect 15200 39918 15252 39924
rect 14740 39908 14792 39914
rect 14740 39850 14792 39856
rect 14648 39500 14700 39506
rect 14648 39442 14700 39448
rect 15212 38826 15240 39918
rect 15396 39438 15424 40054
rect 15384 39432 15436 39438
rect 15384 39374 15436 39380
rect 15384 39296 15436 39302
rect 15384 39238 15436 39244
rect 15396 39030 15424 39238
rect 15384 39024 15436 39030
rect 15384 38966 15436 38972
rect 15292 38956 15344 38962
rect 15292 38898 15344 38904
rect 15200 38820 15252 38826
rect 15200 38762 15252 38768
rect 14648 38752 14700 38758
rect 14648 38694 14700 38700
rect 14280 38548 14332 38554
rect 14280 38490 14332 38496
rect 14188 38344 14240 38350
rect 14188 38286 14240 38292
rect 14200 38010 14228 38286
rect 14188 38004 14240 38010
rect 14188 37946 14240 37952
rect 14108 37862 14228 37890
rect 14292 37874 14320 38490
rect 14200 37806 14228 37862
rect 14280 37868 14332 37874
rect 14280 37810 14332 37816
rect 14188 37800 14240 37806
rect 14188 37742 14240 37748
rect 14292 36786 14320 37810
rect 14464 37732 14516 37738
rect 14464 37674 14516 37680
rect 14372 36916 14424 36922
rect 14372 36858 14424 36864
rect 14280 36780 14332 36786
rect 14280 36722 14332 36728
rect 14292 36310 14320 36722
rect 14384 36666 14412 36858
rect 14476 36786 14504 37674
rect 14660 37262 14688 38694
rect 15212 37874 15240 38762
rect 15200 37868 15252 37874
rect 15200 37810 15252 37816
rect 15304 37856 15332 38898
rect 15384 37868 15436 37874
rect 15304 37828 15384 37856
rect 15200 37732 15252 37738
rect 15200 37674 15252 37680
rect 14924 37392 14976 37398
rect 14924 37334 14976 37340
rect 14556 37256 14608 37262
rect 14556 37198 14608 37204
rect 14648 37256 14700 37262
rect 14936 37210 14964 37334
rect 15212 37262 15240 37674
rect 15304 37398 15332 37828
rect 15384 37810 15436 37816
rect 15488 37670 15516 40326
rect 15672 39846 15700 40870
rect 15660 39840 15712 39846
rect 15660 39782 15712 39788
rect 15672 39574 15700 39782
rect 15660 39568 15712 39574
rect 15660 39510 15712 39516
rect 15764 39420 15792 41074
rect 16040 40934 16068 42026
rect 16212 42016 16264 42022
rect 16212 41958 16264 41964
rect 16028 40928 16080 40934
rect 16028 40870 16080 40876
rect 16224 39982 16252 41958
rect 16408 40730 16436 42094
rect 16672 42016 16724 42022
rect 16672 41958 16724 41964
rect 16684 41614 16712 41958
rect 16672 41608 16724 41614
rect 16672 41550 16724 41556
rect 16764 41132 16816 41138
rect 16764 41074 16816 41080
rect 16396 40724 16448 40730
rect 16396 40666 16448 40672
rect 16580 40520 16632 40526
rect 16580 40462 16632 40468
rect 16592 40050 16620 40462
rect 16580 40044 16632 40050
rect 16580 39986 16632 39992
rect 16212 39976 16264 39982
rect 16212 39918 16264 39924
rect 16776 39642 16804 41074
rect 17236 40662 17264 42094
rect 17316 41472 17368 41478
rect 17316 41414 17368 41420
rect 17224 40656 17276 40662
rect 17224 40598 17276 40604
rect 17132 40452 17184 40458
rect 17132 40394 17184 40400
rect 16948 40384 17000 40390
rect 16948 40326 17000 40332
rect 16764 39636 16816 39642
rect 16764 39578 16816 39584
rect 16960 39438 16988 40326
rect 17144 40050 17172 40394
rect 17236 40118 17264 40598
rect 17328 40526 17356 41414
rect 17590 41370 17646 42406
rect 20444 42356 20496 42362
rect 20444 42298 20496 42304
rect 20456 42226 20484 42298
rect 18144 42220 18196 42226
rect 18144 42162 18196 42168
rect 19892 42220 19944 42226
rect 19892 42162 19944 42168
rect 20444 42220 20496 42226
rect 20444 42162 20496 42168
rect 18052 42152 18104 42158
rect 18052 42094 18104 42100
rect 17590 41318 17592 41370
rect 17644 41318 17646 41370
rect 17316 40520 17368 40526
rect 17316 40462 17368 40468
rect 17224 40112 17276 40118
rect 17224 40054 17276 40060
rect 17132 40044 17184 40050
rect 17132 39986 17184 39992
rect 17328 39506 17356 40462
rect 17590 40282 17646 41318
rect 18064 40934 18092 42094
rect 18052 40928 18104 40934
rect 18052 40870 18104 40876
rect 18064 40526 18092 40870
rect 18052 40520 18104 40526
rect 18052 40462 18104 40468
rect 17590 40230 17592 40282
rect 17644 40230 17646 40282
rect 17316 39500 17368 39506
rect 17316 39442 17368 39448
rect 17500 39500 17552 39506
rect 17500 39442 17552 39448
rect 15844 39432 15896 39438
rect 15764 39392 15844 39420
rect 15844 39374 15896 39380
rect 16948 39432 17000 39438
rect 16948 39374 17000 39380
rect 15568 38888 15620 38894
rect 15568 38830 15620 38836
rect 15580 37874 15608 38830
rect 15856 37942 15884 39374
rect 17408 39364 17460 39370
rect 17408 39306 17460 39312
rect 17420 38962 17448 39306
rect 15936 38956 15988 38962
rect 15936 38898 15988 38904
rect 17224 38956 17276 38962
rect 17224 38898 17276 38904
rect 17408 38956 17460 38962
rect 17408 38898 17460 38904
rect 15844 37936 15896 37942
rect 15844 37878 15896 37884
rect 15568 37868 15620 37874
rect 15568 37810 15620 37816
rect 15476 37664 15528 37670
rect 15476 37606 15528 37612
rect 15752 37664 15804 37670
rect 15752 37606 15804 37612
rect 15292 37392 15344 37398
rect 15292 37334 15344 37340
rect 15660 37324 15712 37330
rect 15660 37266 15712 37272
rect 14648 37198 14700 37204
rect 14568 36922 14596 37198
rect 14844 37194 14964 37210
rect 15200 37256 15252 37262
rect 15200 37198 15252 37204
rect 15292 37256 15344 37262
rect 15292 37198 15344 37204
rect 14832 37188 14964 37194
rect 14884 37182 14964 37188
rect 14832 37130 14884 37136
rect 14556 36916 14608 36922
rect 14556 36858 14608 36864
rect 14464 36780 14516 36786
rect 14464 36722 14516 36728
rect 14924 36780 14976 36786
rect 14924 36722 14976 36728
rect 14556 36712 14608 36718
rect 14384 36660 14556 36666
rect 14384 36654 14608 36660
rect 14384 36638 14596 36654
rect 14280 36304 14332 36310
rect 14280 36246 14332 36252
rect 14004 36168 14056 36174
rect 14004 36110 14056 36116
rect 14556 36168 14608 36174
rect 14556 36110 14608 36116
rect 14648 36168 14700 36174
rect 14648 36110 14700 36116
rect 13544 35692 13596 35698
rect 13544 35634 13596 35640
rect 13728 35692 13780 35698
rect 13728 35634 13780 35640
rect 13372 35550 13492 35578
rect 13372 35018 13400 35550
rect 13544 35216 13596 35222
rect 13544 35158 13596 35164
rect 13360 35012 13412 35018
rect 13360 34954 13412 34960
rect 13268 34536 13320 34542
rect 13268 34478 13320 34484
rect 13176 33448 13228 33454
rect 13176 33390 13228 33396
rect 13188 32978 13216 33390
rect 13176 32972 13228 32978
rect 13176 32914 13228 32920
rect 13084 32904 13136 32910
rect 13084 32846 13136 32852
rect 13096 31142 13124 32846
rect 13176 32768 13228 32774
rect 13176 32710 13228 32716
rect 13188 31346 13216 32710
rect 13280 31482 13308 34478
rect 13372 33930 13400 34954
rect 13556 34610 13584 35158
rect 14568 35154 14596 36110
rect 14660 35766 14688 36110
rect 14648 35760 14700 35766
rect 14648 35702 14700 35708
rect 14556 35148 14608 35154
rect 14556 35090 14608 35096
rect 14568 34746 14596 35090
rect 14660 35018 14688 35702
rect 14936 35290 14964 36722
rect 15212 36310 15240 37198
rect 15304 36854 15332 37198
rect 15292 36848 15344 36854
rect 15292 36790 15344 36796
rect 15672 36718 15700 37266
rect 15764 36922 15792 37606
rect 15948 37466 15976 38898
rect 16580 38752 16632 38758
rect 16580 38694 16632 38700
rect 15936 37460 15988 37466
rect 15936 37402 15988 37408
rect 16488 37392 16540 37398
rect 16488 37334 16540 37340
rect 15844 37120 15896 37126
rect 15844 37062 15896 37068
rect 15856 36922 15884 37062
rect 15752 36916 15804 36922
rect 15752 36858 15804 36864
rect 15844 36916 15896 36922
rect 15844 36858 15896 36864
rect 15660 36712 15712 36718
rect 15660 36654 15712 36660
rect 15384 36576 15436 36582
rect 15384 36518 15436 36524
rect 15752 36576 15804 36582
rect 15752 36518 15804 36524
rect 15200 36304 15252 36310
rect 15200 36246 15252 36252
rect 15212 35986 15240 36246
rect 15120 35958 15240 35986
rect 15120 35766 15148 35958
rect 15108 35760 15160 35766
rect 15108 35702 15160 35708
rect 15200 35488 15252 35494
rect 15200 35430 15252 35436
rect 15292 35488 15344 35494
rect 15292 35430 15344 35436
rect 14924 35284 14976 35290
rect 14924 35226 14976 35232
rect 14648 35012 14700 35018
rect 14648 34954 14700 34960
rect 14556 34740 14608 34746
rect 14556 34682 14608 34688
rect 14660 34610 14688 34954
rect 15212 34610 15240 35430
rect 15304 34678 15332 35430
rect 15396 35086 15424 36518
rect 15764 36174 15792 36518
rect 15752 36168 15804 36174
rect 15752 36110 15804 36116
rect 15844 36032 15896 36038
rect 15844 35974 15896 35980
rect 16028 36032 16080 36038
rect 16028 35974 16080 35980
rect 15856 35766 15884 35974
rect 15844 35760 15896 35766
rect 15844 35702 15896 35708
rect 15568 35692 15620 35698
rect 15568 35634 15620 35640
rect 15580 35290 15608 35634
rect 15660 35624 15712 35630
rect 15660 35566 15712 35572
rect 15936 35624 15988 35630
rect 15936 35566 15988 35572
rect 15568 35284 15620 35290
rect 15568 35226 15620 35232
rect 15384 35080 15436 35086
rect 15384 35022 15436 35028
rect 15384 34944 15436 34950
rect 15384 34886 15436 34892
rect 15396 34746 15424 34886
rect 15384 34740 15436 34746
rect 15384 34682 15436 34688
rect 15568 34740 15620 34746
rect 15568 34682 15620 34688
rect 15292 34672 15344 34678
rect 15292 34614 15344 34620
rect 13544 34604 13596 34610
rect 13544 34546 13596 34552
rect 14188 34604 14240 34610
rect 14188 34546 14240 34552
rect 14648 34604 14700 34610
rect 14648 34546 14700 34552
rect 15200 34604 15252 34610
rect 15200 34546 15252 34552
rect 15476 34604 15528 34610
rect 15476 34546 15528 34552
rect 13452 34536 13504 34542
rect 13452 34478 13504 34484
rect 13360 33924 13412 33930
rect 13360 33866 13412 33872
rect 13372 32570 13400 33866
rect 13464 33862 13492 34478
rect 14200 33998 14228 34546
rect 14188 33992 14240 33998
rect 14188 33934 14240 33940
rect 14464 33992 14516 33998
rect 14464 33934 14516 33940
rect 13452 33856 13504 33862
rect 13452 33798 13504 33804
rect 14280 33856 14332 33862
rect 14280 33798 14332 33804
rect 14292 33590 14320 33798
rect 14280 33584 14332 33590
rect 14280 33526 14332 33532
rect 13728 33516 13780 33522
rect 13728 33458 13780 33464
rect 13360 32564 13412 32570
rect 13360 32506 13412 32512
rect 13360 31816 13412 31822
rect 13360 31758 13412 31764
rect 13268 31476 13320 31482
rect 13268 31418 13320 31424
rect 13176 31340 13228 31346
rect 13176 31282 13228 31288
rect 13268 31340 13320 31346
rect 13268 31282 13320 31288
rect 13084 31136 13136 31142
rect 13084 31078 13136 31084
rect 13096 30734 13124 31078
rect 13084 30728 13136 30734
rect 13084 30670 13136 30676
rect 12992 30252 13044 30258
rect 12992 30194 13044 30200
rect 12912 29974 13032 30002
rect 12900 29844 12952 29850
rect 12900 29786 12952 29792
rect 12728 29294 12848 29322
rect 12532 29096 12584 29102
rect 12532 29038 12584 29044
rect 12728 28966 12756 29294
rect 12912 29238 12940 29786
rect 13004 29646 13032 29974
rect 13096 29850 13124 30670
rect 13084 29844 13136 29850
rect 13084 29786 13136 29792
rect 12992 29640 13044 29646
rect 12992 29582 13044 29588
rect 13188 29510 13216 31282
rect 13176 29504 13228 29510
rect 13176 29446 13228 29452
rect 12900 29232 12952 29238
rect 12900 29174 12952 29180
rect 12992 29096 13044 29102
rect 12992 29038 13044 29044
rect 12716 28960 12768 28966
rect 12716 28902 12768 28908
rect 12438 28806 12440 28858
rect 12492 28806 12494 28858
rect 12348 28756 12400 28762
rect 12348 28698 12400 28704
rect 12176 28206 12296 28234
rect 12348 28212 12400 28218
rect 12072 27464 12124 27470
rect 12072 27406 12124 27412
rect 11900 25622 12020 25650
rect 11704 25492 11756 25498
rect 11704 25434 11756 25440
rect 11612 25152 11664 25158
rect 11612 25094 11664 25100
rect 11520 24880 11572 24886
rect 11520 24822 11572 24828
rect 11624 24818 11652 25094
rect 11796 24948 11848 24954
rect 11796 24890 11848 24896
rect 11612 24812 11664 24818
rect 11612 24754 11664 24760
rect 11428 24404 11480 24410
rect 11428 24346 11480 24352
rect 11336 24200 11388 24206
rect 11256 24160 11336 24188
rect 11336 24142 11388 24148
rect 11808 24138 11836 24890
rect 11428 24132 11480 24138
rect 11428 24074 11480 24080
rect 11796 24132 11848 24138
rect 11796 24074 11848 24080
rect 11440 23798 11468 24074
rect 11072 23718 11192 23746
rect 11428 23792 11480 23798
rect 11428 23734 11480 23740
rect 10876 23180 10928 23186
rect 10876 23122 10928 23128
rect 10784 23112 10836 23118
rect 10784 23054 10836 23060
rect 10796 22522 10824 23054
rect 10968 23044 11020 23050
rect 10968 22986 11020 22992
rect 10980 22642 11008 22986
rect 10968 22636 11020 22642
rect 10968 22578 11020 22584
rect 10796 22494 11008 22522
rect 10876 22024 10928 22030
rect 10876 21966 10928 21972
rect 10784 21888 10836 21894
rect 10784 21830 10836 21836
rect 10796 21554 10824 21830
rect 10888 21690 10916 21966
rect 10980 21894 11008 22494
rect 10968 21888 11020 21894
rect 10968 21830 11020 21836
rect 10876 21684 10928 21690
rect 10876 21626 10928 21632
rect 10612 21508 10732 21536
rect 10784 21548 10836 21554
rect 10508 20596 10560 20602
rect 10508 20538 10560 20544
rect 10336 20284 10456 20312
rect 10336 18154 10364 20284
rect 10416 19916 10468 19922
rect 10416 19858 10468 19864
rect 10428 18290 10456 19858
rect 10520 19854 10548 20538
rect 10508 19848 10560 19854
rect 10508 19790 10560 19796
rect 10520 18970 10548 19790
rect 10612 19428 10640 21508
rect 10784 21490 10836 21496
rect 10876 21412 10928 21418
rect 10796 21372 10876 21400
rect 10796 21332 10824 21372
rect 10876 21354 10928 21360
rect 10704 21304 10824 21332
rect 10704 20942 10732 21304
rect 10980 21298 11008 21830
rect 10888 21270 11008 21298
rect 10784 21140 10836 21146
rect 10784 21082 10836 21088
rect 10692 20936 10744 20942
rect 10692 20878 10744 20884
rect 10692 20596 10744 20602
rect 10692 20538 10744 20544
rect 10704 19990 10732 20538
rect 10796 20466 10824 21082
rect 10784 20460 10836 20466
rect 10784 20402 10836 20408
rect 10692 19984 10744 19990
rect 10692 19926 10744 19932
rect 10888 19768 10916 21270
rect 11072 21146 11100 23718
rect 11152 22568 11204 22574
rect 11152 22510 11204 22516
rect 11060 21140 11112 21146
rect 11060 21082 11112 21088
rect 11060 20800 11112 20806
rect 11060 20742 11112 20748
rect 11072 20534 11100 20742
rect 11060 20528 11112 20534
rect 11060 20470 11112 20476
rect 11060 20256 11112 20262
rect 11060 20198 11112 20204
rect 11072 19786 11100 20198
rect 11060 19780 11112 19786
rect 10888 19740 11008 19768
rect 10784 19440 10836 19446
rect 10612 19400 10732 19428
rect 10600 19236 10652 19242
rect 10600 19178 10652 19184
rect 10612 18970 10640 19178
rect 10508 18964 10560 18970
rect 10508 18906 10560 18912
rect 10600 18964 10652 18970
rect 10600 18906 10652 18912
rect 10600 18828 10652 18834
rect 10600 18770 10652 18776
rect 10416 18284 10468 18290
rect 10416 18226 10468 18232
rect 10324 18148 10376 18154
rect 10324 18090 10376 18096
rect 10428 17678 10456 18226
rect 10612 18222 10640 18770
rect 10600 18216 10652 18222
rect 10600 18158 10652 18164
rect 10416 17672 10468 17678
rect 10336 17632 10416 17660
rect 10232 17060 10284 17066
rect 10232 17002 10284 17008
rect 10336 16114 10364 17632
rect 10416 17614 10468 17620
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10508 16584 10560 16590
rect 10508 16526 10560 16532
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 10520 15638 10548 16526
rect 10612 16454 10640 17070
rect 10600 16448 10652 16454
rect 10600 16390 10652 16396
rect 10508 15632 10560 15638
rect 10508 15574 10560 15580
rect 10508 15360 10560 15366
rect 10508 15302 10560 15308
rect 10520 15026 10548 15302
rect 10508 15020 10560 15026
rect 10508 14962 10560 14968
rect 10520 14618 10548 14962
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10508 14068 10560 14074
rect 10508 14010 10560 14016
rect 10520 13938 10548 14010
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 10140 10736 10192 10742
rect 10244 10724 10272 13874
rect 10416 13456 10468 13462
rect 10416 13398 10468 13404
rect 10428 12646 10456 13398
rect 10416 12640 10468 12646
rect 10416 12582 10468 12588
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10336 11150 10364 11630
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 10192 10696 10272 10724
rect 10140 10678 10192 10684
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 9956 7472 10008 7478
rect 9956 7414 10008 7420
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9784 6322 9812 6802
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9968 5778 9996 7414
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9404 5296 9456 5302
rect 9404 5238 9456 5244
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 9324 4146 9352 4626
rect 9312 4140 9364 4146
rect 9232 4100 9312 4128
rect 9232 3670 9260 4100
rect 9312 4082 9364 4088
rect 9220 3664 9272 3670
rect 9220 3606 9272 3612
rect 9232 3534 9260 3606
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 8116 2848 8168 2854
rect 8116 2790 8168 2796
rect 8128 2514 8156 2790
rect 8116 2508 8168 2514
rect 8116 2450 8168 2456
rect 8220 2106 8248 2926
rect 8956 2650 8984 2994
rect 8944 2644 8996 2650
rect 8944 2586 8996 2592
rect 8208 2100 8260 2106
rect 8208 2042 8260 2048
rect 7380 1352 7432 1358
rect 7380 1294 7432 1300
rect 7840 1352 7892 1358
rect 7840 1294 7892 1300
rect 8392 1352 8444 1358
rect 8392 1294 8444 1300
rect 9220 1352 9272 1358
rect 9220 1294 9272 1300
rect 8300 1284 8352 1290
rect 8300 1226 8352 1232
rect 7286 1062 7288 1114
rect 7340 1062 7342 1114
rect 7286 1040 7342 1062
rect 8312 800 8340 1226
rect 8404 950 8432 1294
rect 8392 944 8444 950
rect 8392 886 8444 892
rect 9232 882 9260 1294
rect 9416 1290 9444 5238
rect 9508 5166 9536 5714
rect 10152 5234 10180 8230
rect 10244 8022 10272 10542
rect 10336 10538 10364 11086
rect 10324 10532 10376 10538
rect 10324 10474 10376 10480
rect 10324 9512 10376 9518
rect 10324 9454 10376 9460
rect 10232 8016 10284 8022
rect 10232 7958 10284 7964
rect 10336 7410 10364 9454
rect 10428 7886 10456 11154
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10612 8974 10640 9318
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10244 7002 10272 7346
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10244 6338 10272 6734
rect 10336 6458 10364 7142
rect 10428 6798 10456 7686
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10324 6452 10376 6458
rect 10324 6394 10376 6400
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10428 6338 10456 6394
rect 10244 6310 10456 6338
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 9496 5160 9548 5166
rect 9496 5102 9548 5108
rect 9956 5160 10008 5166
rect 9956 5102 10008 5108
rect 9508 4486 9536 5102
rect 9772 5092 9824 5098
rect 9772 5034 9824 5040
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9496 4480 9548 4486
rect 9496 4422 9548 4428
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9508 3534 9536 4014
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 9600 3058 9628 4558
rect 9692 3194 9720 4762
rect 9784 3534 9812 5034
rect 9968 4282 9996 5102
rect 10324 4548 10376 4554
rect 10324 4490 10376 4496
rect 10336 4282 10364 4490
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 10324 4276 10376 4282
rect 10324 4218 10376 4224
rect 9968 4146 9996 4218
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9600 2446 9628 2994
rect 9784 2774 9812 3470
rect 9784 2746 9904 2774
rect 9876 2650 9904 2746
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 9600 1970 9628 2382
rect 9588 1964 9640 1970
rect 9588 1906 9640 1912
rect 9680 1964 9732 1970
rect 9680 1906 9732 1912
rect 9404 1284 9456 1290
rect 9404 1226 9456 1232
rect 9692 1222 9720 1906
rect 9968 1426 9996 4082
rect 10428 3534 10456 6190
rect 10520 5642 10548 8298
rect 10612 8090 10640 8434
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10600 7200 10652 7206
rect 10600 7142 10652 7148
rect 10612 6934 10640 7142
rect 10600 6928 10652 6934
rect 10600 6870 10652 6876
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10612 6118 10640 6734
rect 10600 6112 10652 6118
rect 10600 6054 10652 6060
rect 10508 5636 10560 5642
rect 10508 5578 10560 5584
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 9956 1420 10008 1426
rect 9956 1362 10008 1368
rect 10060 1358 10088 3334
rect 10520 2446 10548 5170
rect 10612 3942 10640 6054
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10612 3126 10640 3878
rect 10704 3670 10732 19400
rect 10784 19382 10836 19388
rect 10796 18714 10824 19382
rect 10796 18686 10916 18714
rect 10784 18624 10836 18630
rect 10784 18566 10836 18572
rect 10796 17814 10824 18566
rect 10888 18290 10916 18686
rect 10980 18630 11008 19740
rect 11060 19722 11112 19728
rect 11060 19168 11112 19174
rect 11060 19110 11112 19116
rect 11072 18766 11100 19110
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 10968 18624 11020 18630
rect 10968 18566 11020 18572
rect 10876 18284 10928 18290
rect 10876 18226 10928 18232
rect 10784 17808 10836 17814
rect 10784 17750 10836 17756
rect 10888 16998 10916 18226
rect 10968 18148 11020 18154
rect 10968 18090 11020 18096
rect 11060 18148 11112 18154
rect 11060 18090 11112 18096
rect 10876 16992 10928 16998
rect 10876 16934 10928 16940
rect 10980 16522 11008 18090
rect 11072 16590 11100 18090
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 10968 16516 11020 16522
rect 10968 16458 11020 16464
rect 10784 16448 10836 16454
rect 10784 16390 10836 16396
rect 10796 16114 10824 16390
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 11072 13954 11100 14894
rect 10888 13938 11100 13954
rect 10876 13932 11100 13938
rect 10928 13926 11100 13932
rect 10876 13874 10928 13880
rect 11072 13734 11100 13926
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10796 12238 10824 12786
rect 11072 12238 11100 13670
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 10796 8566 10824 12174
rect 11072 10606 11100 12174
rect 11164 11898 11192 22510
rect 11244 22500 11296 22506
rect 11244 22442 11296 22448
rect 11256 22098 11284 22442
rect 11244 22092 11296 22098
rect 11244 22034 11296 22040
rect 11612 21888 11664 21894
rect 11612 21830 11664 21836
rect 11244 21548 11296 21554
rect 11244 21490 11296 21496
rect 11256 20942 11284 21490
rect 11624 21350 11652 21830
rect 11704 21548 11756 21554
rect 11704 21490 11756 21496
rect 11612 21344 11664 21350
rect 11612 21286 11664 21292
rect 11244 20936 11296 20942
rect 11716 20890 11744 21490
rect 11244 20878 11296 20884
rect 11624 20862 11744 20890
rect 11796 20936 11848 20942
rect 11796 20878 11848 20884
rect 11256 20726 11560 20754
rect 11256 20602 11284 20726
rect 11244 20596 11296 20602
rect 11244 20538 11296 20544
rect 11336 20596 11388 20602
rect 11336 20538 11388 20544
rect 11244 20392 11296 20398
rect 11244 20334 11296 20340
rect 11256 19854 11284 20334
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11256 19242 11284 19790
rect 11348 19378 11376 20538
rect 11532 19854 11560 20726
rect 11624 20466 11652 20862
rect 11808 20466 11836 20878
rect 11900 20534 11928 25622
rect 11980 25492 12032 25498
rect 11980 25434 12032 25440
rect 11992 25226 12020 25434
rect 12084 25294 12112 27406
rect 12072 25288 12124 25294
rect 12072 25230 12124 25236
rect 11980 25220 12032 25226
rect 11980 25162 12032 25168
rect 12176 24954 12204 28206
rect 12348 28154 12400 28160
rect 12256 26988 12308 26994
rect 12256 26930 12308 26936
rect 12268 26382 12296 26930
rect 12256 26376 12308 26382
rect 12256 26318 12308 26324
rect 12360 25974 12388 28154
rect 12438 27770 12494 28806
rect 12624 28756 12676 28762
rect 12624 28698 12676 28704
rect 12532 28552 12584 28558
rect 12532 28494 12584 28500
rect 12438 27718 12440 27770
rect 12492 27718 12494 27770
rect 12438 26682 12494 27718
rect 12544 27130 12572 28494
rect 12532 27124 12584 27130
rect 12532 27066 12584 27072
rect 12636 26874 12664 28698
rect 12728 28218 12756 28902
rect 12808 28552 12860 28558
rect 12808 28494 12860 28500
rect 12716 28212 12768 28218
rect 12716 28154 12768 28160
rect 12820 28064 12848 28494
rect 12728 28036 12848 28064
rect 12728 26994 12756 28036
rect 12808 27940 12860 27946
rect 12808 27882 12860 27888
rect 12820 27538 12848 27882
rect 12808 27532 12860 27538
rect 12808 27474 12860 27480
rect 12900 27464 12952 27470
rect 12900 27406 12952 27412
rect 12808 27396 12860 27402
rect 12808 27338 12860 27344
rect 12716 26988 12768 26994
rect 12716 26930 12768 26936
rect 12636 26846 12756 26874
rect 12438 26630 12440 26682
rect 12492 26630 12494 26682
rect 12348 25968 12400 25974
rect 12348 25910 12400 25916
rect 12438 25594 12494 26630
rect 12728 26450 12756 26846
rect 12532 26444 12584 26450
rect 12532 26386 12584 26392
rect 12716 26444 12768 26450
rect 12716 26386 12768 26392
rect 12438 25542 12440 25594
rect 12492 25542 12494 25594
rect 12256 25288 12308 25294
rect 12256 25230 12308 25236
rect 12164 24948 12216 24954
rect 12164 24890 12216 24896
rect 12164 24132 12216 24138
rect 12164 24074 12216 24080
rect 12176 23866 12204 24074
rect 12164 23860 12216 23866
rect 12164 23802 12216 23808
rect 12268 23050 12296 25230
rect 12348 25152 12400 25158
rect 12348 25094 12400 25100
rect 12164 23044 12216 23050
rect 12164 22986 12216 22992
rect 12256 23044 12308 23050
rect 12256 22986 12308 22992
rect 12072 22772 12124 22778
rect 12072 22714 12124 22720
rect 12084 20942 12112 22714
rect 12176 22234 12204 22986
rect 12268 22574 12296 22986
rect 12256 22568 12308 22574
rect 12256 22510 12308 22516
rect 12164 22228 12216 22234
rect 12164 22170 12216 22176
rect 12164 22092 12216 22098
rect 12164 22034 12216 22040
rect 12176 21554 12204 22034
rect 12360 22030 12388 25094
rect 12438 24506 12494 25542
rect 12544 25294 12572 26386
rect 12716 26308 12768 26314
rect 12636 26268 12716 26296
rect 12636 25702 12664 26268
rect 12716 26250 12768 26256
rect 12820 26042 12848 27338
rect 12912 27130 12940 27406
rect 12900 27124 12952 27130
rect 12900 27066 12952 27072
rect 12900 26988 12952 26994
rect 12900 26930 12952 26936
rect 12912 26450 12940 26930
rect 12900 26444 12952 26450
rect 12900 26386 12952 26392
rect 12912 26042 12940 26386
rect 12808 26036 12860 26042
rect 12808 25978 12860 25984
rect 12900 26036 12952 26042
rect 12900 25978 12952 25984
rect 12716 25968 12768 25974
rect 12716 25910 12768 25916
rect 12624 25696 12676 25702
rect 12624 25638 12676 25644
rect 12728 25362 12756 25910
rect 12820 25838 12848 25978
rect 12808 25832 12860 25838
rect 12808 25774 12860 25780
rect 12716 25356 12768 25362
rect 12716 25298 12768 25304
rect 12820 25294 12848 25774
rect 13004 25480 13032 29038
rect 13176 28484 13228 28490
rect 13176 28426 13228 28432
rect 13084 27872 13136 27878
rect 13084 27814 13136 27820
rect 13096 27470 13124 27814
rect 13188 27470 13216 28426
rect 13084 27464 13136 27470
rect 13084 27406 13136 27412
rect 13176 27464 13228 27470
rect 13176 27406 13228 27412
rect 13176 27124 13228 27130
rect 13176 27066 13228 27072
rect 13084 25696 13136 25702
rect 13084 25638 13136 25644
rect 12912 25452 13032 25480
rect 12532 25288 12584 25294
rect 12532 25230 12584 25236
rect 12808 25288 12860 25294
rect 12808 25230 12860 25236
rect 12438 24454 12440 24506
rect 12492 24454 12494 24506
rect 12438 23418 12494 24454
rect 12544 23662 12572 25230
rect 12912 24834 12940 25452
rect 12992 25356 13044 25362
rect 12992 25298 13044 25304
rect 12728 24806 12940 24834
rect 12624 24404 12676 24410
rect 12624 24346 12676 24352
rect 12532 23656 12584 23662
rect 12532 23598 12584 23604
rect 12438 23366 12440 23418
rect 12492 23366 12494 23418
rect 12438 22330 12494 23366
rect 12544 23322 12572 23598
rect 12532 23316 12584 23322
rect 12532 23258 12584 23264
rect 12636 22438 12664 24346
rect 12624 22432 12676 22438
rect 12624 22374 12676 22380
rect 12438 22278 12440 22330
rect 12492 22278 12494 22330
rect 12348 22024 12400 22030
rect 12348 21966 12400 21972
rect 12164 21548 12216 21554
rect 12348 21548 12400 21554
rect 12164 21490 12216 21496
rect 12268 21508 12348 21536
rect 12164 21004 12216 21010
rect 12164 20946 12216 20952
rect 12072 20936 12124 20942
rect 12072 20878 12124 20884
rect 11980 20868 12032 20874
rect 11980 20810 12032 20816
rect 11888 20528 11940 20534
rect 11888 20470 11940 20476
rect 11612 20460 11664 20466
rect 11612 20402 11664 20408
rect 11796 20460 11848 20466
rect 11796 20402 11848 20408
rect 11704 20324 11756 20330
rect 11704 20266 11756 20272
rect 11520 19848 11572 19854
rect 11520 19790 11572 19796
rect 11612 19440 11664 19446
rect 11612 19382 11664 19388
rect 11336 19372 11388 19378
rect 11336 19314 11388 19320
rect 11520 19372 11572 19378
rect 11520 19314 11572 19320
rect 11244 19236 11296 19242
rect 11244 19178 11296 19184
rect 11428 18828 11480 18834
rect 11428 18770 11480 18776
rect 11336 18760 11388 18766
rect 11336 18702 11388 18708
rect 11244 17740 11296 17746
rect 11244 17682 11296 17688
rect 11256 15026 11284 17682
rect 11348 15094 11376 18702
rect 11440 16794 11468 18770
rect 11532 17814 11560 19314
rect 11520 17808 11572 17814
rect 11520 17750 11572 17756
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 11428 16788 11480 16794
rect 11428 16730 11480 16736
rect 11428 16448 11480 16454
rect 11428 16390 11480 16396
rect 11440 15502 11468 16390
rect 11532 16114 11560 17614
rect 11624 17338 11652 19382
rect 11716 19174 11744 20266
rect 11704 19168 11756 19174
rect 11704 19110 11756 19116
rect 11704 18828 11756 18834
rect 11808 18816 11836 20402
rect 11992 19990 12020 20810
rect 12176 20466 12204 20946
rect 12268 20942 12296 21508
rect 12348 21490 12400 21496
rect 12348 21412 12400 21418
rect 12348 21354 12400 21360
rect 12360 21078 12388 21354
rect 12438 21242 12494 22278
rect 12728 22166 12756 24806
rect 12808 24744 12860 24750
rect 12808 24686 12860 24692
rect 12820 24070 12848 24686
rect 12808 24064 12860 24070
rect 12808 24006 12860 24012
rect 12820 23594 12848 24006
rect 12900 23656 12952 23662
rect 12900 23598 12952 23604
rect 12808 23588 12860 23594
rect 12808 23530 12860 23536
rect 12820 23118 12848 23530
rect 12808 23112 12860 23118
rect 12808 23054 12860 23060
rect 12820 22574 12848 23054
rect 12912 22982 12940 23598
rect 12900 22976 12952 22982
rect 12900 22918 12952 22924
rect 12808 22568 12860 22574
rect 12808 22510 12860 22516
rect 12716 22160 12768 22166
rect 12636 22120 12716 22148
rect 12532 22092 12584 22098
rect 12532 22034 12584 22040
rect 12544 21962 12572 22034
rect 12532 21956 12584 21962
rect 12532 21898 12584 21904
rect 12532 21344 12584 21350
rect 12532 21286 12584 21292
rect 12438 21190 12440 21242
rect 12492 21190 12494 21242
rect 12348 21072 12400 21078
rect 12348 21014 12400 21020
rect 12256 20936 12308 20942
rect 12256 20878 12308 20884
rect 12348 20936 12400 20942
rect 12348 20878 12400 20884
rect 12164 20460 12216 20466
rect 12164 20402 12216 20408
rect 12164 20324 12216 20330
rect 12268 20312 12296 20878
rect 12360 20398 12388 20878
rect 12348 20392 12400 20398
rect 12348 20334 12400 20340
rect 12216 20284 12296 20312
rect 12164 20266 12216 20272
rect 11980 19984 12032 19990
rect 11980 19926 12032 19932
rect 11980 19780 12032 19786
rect 11980 19722 12032 19728
rect 11992 19514 12020 19722
rect 12072 19712 12124 19718
rect 12072 19654 12124 19660
rect 11980 19508 12032 19514
rect 11980 19450 12032 19456
rect 12084 19446 12112 19654
rect 12072 19440 12124 19446
rect 12072 19382 12124 19388
rect 12268 18902 12296 20284
rect 12348 20256 12400 20262
rect 12348 20198 12400 20204
rect 12360 19854 12388 20198
rect 12438 20154 12494 21190
rect 12544 20806 12572 21286
rect 12532 20800 12584 20806
rect 12532 20742 12584 20748
rect 12532 20460 12584 20466
rect 12532 20402 12584 20408
rect 12438 20102 12440 20154
rect 12492 20102 12494 20154
rect 12348 19848 12400 19854
rect 12348 19790 12400 19796
rect 12256 18896 12308 18902
rect 12256 18838 12308 18844
rect 11756 18788 11836 18816
rect 11704 18770 11756 18776
rect 12164 18624 12216 18630
rect 12164 18566 12216 18572
rect 11716 18380 12020 18408
rect 11716 18290 11744 18380
rect 11704 18284 11756 18290
rect 11888 18284 11940 18290
rect 11704 18226 11756 18232
rect 11788 18244 11888 18272
rect 11788 18136 11816 18244
rect 11888 18226 11940 18232
rect 11788 18108 11836 18136
rect 11704 17536 11756 17542
rect 11704 17478 11756 17484
rect 11612 17332 11664 17338
rect 11612 17274 11664 17280
rect 11716 17202 11744 17478
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11808 16250 11836 18108
rect 11992 17678 12020 18380
rect 12176 18222 12204 18566
rect 12268 18290 12296 18838
rect 12256 18284 12308 18290
rect 12256 18226 12308 18232
rect 12164 18216 12216 18222
rect 12164 18158 12216 18164
rect 12360 18086 12388 19790
rect 12438 19066 12494 20102
rect 12438 19014 12440 19066
rect 12492 19014 12494 19066
rect 12164 18080 12216 18086
rect 12164 18022 12216 18028
rect 12348 18080 12400 18086
rect 12348 18022 12400 18028
rect 11980 17672 12032 17678
rect 11980 17614 12032 17620
rect 11992 17524 12020 17614
rect 11992 17496 12112 17524
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11796 16244 11848 16250
rect 11796 16186 11848 16192
rect 11520 16108 11572 16114
rect 11520 16050 11572 16056
rect 11428 15496 11480 15502
rect 11900 15450 11928 16934
rect 11980 16788 12032 16794
rect 11980 16730 12032 16736
rect 11992 16590 12020 16730
rect 11980 16584 12032 16590
rect 11980 16526 12032 16532
rect 12084 16046 12112 17496
rect 12176 16998 12204 18022
rect 12438 17978 12494 19014
rect 12544 18986 12572 20402
rect 12636 19378 12664 22120
rect 12716 22102 12768 22108
rect 12716 21344 12768 21350
rect 12716 21286 12768 21292
rect 12728 20942 12756 21286
rect 12820 21010 12848 22510
rect 12912 22098 12940 22918
rect 12900 22092 12952 22098
rect 12900 22034 12952 22040
rect 12900 21072 12952 21078
rect 12900 21014 12952 21020
rect 12808 21004 12860 21010
rect 12808 20946 12860 20952
rect 12716 20936 12768 20942
rect 12716 20878 12768 20884
rect 12820 20398 12848 20946
rect 12808 20392 12860 20398
rect 12808 20334 12860 20340
rect 12912 19514 12940 21014
rect 13004 19786 13032 25298
rect 13096 24886 13124 25638
rect 13188 25158 13216 27066
rect 13176 25152 13228 25158
rect 13176 25094 13228 25100
rect 13084 24880 13136 24886
rect 13084 24822 13136 24828
rect 13084 24268 13136 24274
rect 13084 24210 13136 24216
rect 13096 22030 13124 24210
rect 13188 23118 13216 25094
rect 13176 23112 13228 23118
rect 13176 23054 13228 23060
rect 13084 22024 13136 22030
rect 13136 21984 13216 22012
rect 13084 21966 13136 21972
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 12992 19780 13044 19786
rect 12992 19722 13044 19728
rect 12900 19508 12952 19514
rect 12900 19450 12952 19456
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12544 18958 12756 18986
rect 12624 18896 12676 18902
rect 12624 18838 12676 18844
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 12438 17926 12440 17978
rect 12492 17926 12494 17978
rect 12256 17060 12308 17066
rect 12256 17002 12308 17008
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 12164 16788 12216 16794
rect 12164 16730 12216 16736
rect 12176 16454 12204 16730
rect 12268 16726 12296 17002
rect 12438 16890 12494 17926
rect 12438 16838 12440 16890
rect 12492 16838 12494 16890
rect 12256 16720 12308 16726
rect 12256 16662 12308 16668
rect 12164 16448 12216 16454
rect 12164 16390 12216 16396
rect 12256 16448 12308 16454
rect 12256 16390 12308 16396
rect 12072 16040 12124 16046
rect 12072 15982 12124 15988
rect 12164 15972 12216 15978
rect 12268 15960 12296 16390
rect 12348 16244 12400 16250
rect 12348 16186 12400 16192
rect 12216 15932 12296 15960
rect 12164 15914 12216 15920
rect 12360 15892 12388 16186
rect 12268 15864 12388 15892
rect 11980 15496 12032 15502
rect 11428 15438 11480 15444
rect 11808 15444 11980 15450
rect 11808 15438 12032 15444
rect 11808 15434 12020 15438
rect 11796 15428 12020 15434
rect 11848 15422 12020 15428
rect 11796 15370 11848 15376
rect 12164 15360 12216 15366
rect 12164 15302 12216 15308
rect 12176 15094 12204 15302
rect 11336 15088 11388 15094
rect 11336 15030 11388 15036
rect 12164 15088 12216 15094
rect 12164 15030 12216 15036
rect 11244 15020 11296 15026
rect 11244 14962 11296 14968
rect 11888 14952 11940 14958
rect 11888 14894 11940 14900
rect 11900 14414 11928 14894
rect 11704 14408 11756 14414
rect 11704 14350 11756 14356
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 11624 13938 11652 14214
rect 11612 13932 11664 13938
rect 11612 13874 11664 13880
rect 11716 13734 11744 14350
rect 11980 14340 12032 14346
rect 11980 14282 12032 14288
rect 11992 13938 12020 14282
rect 11980 13932 12032 13938
rect 11980 13874 12032 13880
rect 11520 13728 11572 13734
rect 11520 13670 11572 13676
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11532 13462 11560 13670
rect 11520 13456 11572 13462
rect 11520 13398 11572 13404
rect 12176 13326 12204 14350
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 11336 13252 11388 13258
rect 11336 13194 11388 13200
rect 11348 12646 11376 13194
rect 11520 12912 11572 12918
rect 11520 12854 11572 12860
rect 11336 12640 11388 12646
rect 11336 12582 11388 12588
rect 11532 12374 11560 12854
rect 11888 12776 11940 12782
rect 11888 12718 11940 12724
rect 12268 12730 12296 15864
rect 12438 15802 12494 16838
rect 12438 15750 12440 15802
rect 12492 15750 12494 15802
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 12360 13870 12388 15438
rect 12438 14714 12494 15750
rect 12438 14662 12440 14714
rect 12492 14662 12494 14714
rect 12348 13864 12400 13870
rect 12348 13806 12400 13812
rect 12438 13626 12494 14662
rect 12438 13574 12440 13626
rect 12492 13574 12494 13626
rect 12348 13184 12400 13190
rect 12348 13126 12400 13132
rect 12360 12850 12388 13126
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 11900 12434 11928 12718
rect 12268 12702 12388 12730
rect 11900 12406 12020 12434
rect 11520 12368 11572 12374
rect 11520 12310 11572 12316
rect 11244 12164 11296 12170
rect 11244 12106 11296 12112
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 11164 10266 11192 10406
rect 11152 10260 11204 10266
rect 11152 10202 11204 10208
rect 11164 9674 11192 10202
rect 11256 10198 11284 12106
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11808 11150 11836 11630
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11244 10192 11296 10198
rect 11244 10134 11296 10140
rect 11532 9994 11560 10406
rect 11808 10062 11836 11086
rect 11888 10600 11940 10606
rect 11888 10542 11940 10548
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 11520 9988 11572 9994
rect 11520 9930 11572 9936
rect 10980 9646 11192 9674
rect 10980 9570 11008 9646
rect 11900 9586 11928 10542
rect 11992 10470 12020 12406
rect 12072 11756 12124 11762
rect 12124 11716 12296 11744
rect 12072 11698 12124 11704
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11152 9580 11204 9586
rect 10968 9564 11020 9570
rect 10876 9512 10928 9518
rect 10968 9506 11020 9512
rect 11072 9540 11152 9568
rect 11072 9466 11100 9540
rect 11152 9522 11204 9528
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 10928 9460 11100 9466
rect 10876 9454 11100 9460
rect 10888 9438 11100 9454
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 10784 8560 10836 8566
rect 10784 8502 10836 8508
rect 11256 8430 11284 9318
rect 11520 9104 11572 9110
rect 11520 9046 11572 9052
rect 10968 8424 11020 8430
rect 10968 8366 11020 8372
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 10980 7886 11008 8366
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10784 7812 10836 7818
rect 10784 7754 10836 7760
rect 10796 7546 10824 7754
rect 10980 7546 11008 7822
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 11336 7472 11388 7478
rect 11336 7414 11388 7420
rect 11348 6866 11376 7414
rect 11532 7410 11560 9046
rect 11624 8022 11652 9522
rect 11992 9382 12020 10406
rect 12072 9988 12124 9994
rect 12072 9930 12124 9936
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 11704 8900 11756 8906
rect 11704 8842 11756 8848
rect 11612 8016 11664 8022
rect 11612 7958 11664 7964
rect 11716 7886 11744 8842
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11348 4690 11376 6802
rect 11532 6322 11560 7346
rect 11520 6316 11572 6322
rect 11520 6258 11572 6264
rect 11716 5846 11744 7822
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11704 5840 11756 5846
rect 11704 5782 11756 5788
rect 11336 4684 11388 4690
rect 11336 4626 11388 4632
rect 10692 3664 10744 3670
rect 10692 3606 10744 3612
rect 11348 3602 11376 4626
rect 11716 4146 11744 5782
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10600 3120 10652 3126
rect 10600 3062 10652 3068
rect 10508 2440 10560 2446
rect 10508 2382 10560 2388
rect 10232 2372 10284 2378
rect 10232 2314 10284 2320
rect 10244 1562 10272 2314
rect 10232 1556 10284 1562
rect 10232 1498 10284 1504
rect 10612 1358 10640 3062
rect 10704 2650 10732 3470
rect 10968 3460 11020 3466
rect 10968 3402 11020 3408
rect 10980 2922 11008 3402
rect 11348 3126 11376 3538
rect 11808 3534 11836 4966
rect 11900 4214 11928 6598
rect 11992 5710 12020 6734
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11888 4208 11940 4214
rect 11888 4150 11940 4156
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 11336 3120 11388 3126
rect 11336 3062 11388 3068
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 11060 2916 11112 2922
rect 11060 2858 11112 2864
rect 11072 2666 11100 2858
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 10888 2638 11100 2666
rect 10888 2582 10916 2638
rect 10876 2576 10928 2582
rect 10876 2518 10928 2524
rect 11348 2514 11376 3062
rect 11624 3058 11652 3334
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 11336 2508 11388 2514
rect 11336 2450 11388 2456
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 11072 2106 11100 2246
rect 11060 2100 11112 2106
rect 11060 2042 11112 2048
rect 11348 1970 11376 2450
rect 11336 1964 11388 1970
rect 11336 1906 11388 1912
rect 11716 1358 11744 3130
rect 12084 2310 12112 9930
rect 12164 9580 12216 9586
rect 12164 9522 12216 9528
rect 12176 9110 12204 9522
rect 12164 9104 12216 9110
rect 12164 9046 12216 9052
rect 12268 7290 12296 11716
rect 12360 11354 12388 12702
rect 12438 12538 12494 13574
rect 12544 12850 12572 18226
rect 12636 17814 12664 18838
rect 12624 17808 12676 17814
rect 12624 17750 12676 17756
rect 12624 16788 12676 16794
rect 12728 16776 12756 18958
rect 12808 18896 12860 18902
rect 12808 18838 12860 18844
rect 12820 18154 12848 18838
rect 12912 18698 12940 19450
rect 12900 18692 12952 18698
rect 12900 18634 12952 18640
rect 12808 18148 12860 18154
rect 12808 18090 12860 18096
rect 12900 18080 12952 18086
rect 12900 18022 12952 18028
rect 12676 16748 12756 16776
rect 12624 16730 12676 16736
rect 12636 16114 12664 16730
rect 12808 16516 12860 16522
rect 12808 16458 12860 16464
rect 12624 16108 12676 16114
rect 12624 16050 12676 16056
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12636 13326 12664 14010
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12820 13190 12848 16458
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 12532 12844 12584 12850
rect 12532 12786 12584 12792
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 12438 12486 12440 12538
rect 12492 12486 12494 12538
rect 12438 11450 12494 12486
rect 12544 11778 12572 12786
rect 12636 12238 12664 12786
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12544 11762 12664 11778
rect 12820 11762 12848 12038
rect 12544 11756 12676 11762
rect 12544 11750 12624 11756
rect 12808 11756 12860 11762
rect 12624 11698 12676 11704
rect 12728 11716 12808 11744
rect 12438 11398 12440 11450
rect 12492 11398 12494 11450
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 12438 10362 12494 11398
rect 12636 11218 12664 11698
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 12636 10742 12664 11154
rect 12728 11082 12756 11716
rect 12808 11698 12860 11704
rect 12912 11626 12940 18022
rect 13004 17814 13032 19722
rect 13096 19514 13124 19790
rect 13084 19508 13136 19514
rect 13084 19450 13136 19456
rect 13084 19372 13136 19378
rect 13084 19314 13136 19320
rect 12992 17808 13044 17814
rect 12992 17750 13044 17756
rect 12992 14272 13044 14278
rect 12992 14214 13044 14220
rect 13004 14006 13032 14214
rect 12992 14000 13044 14006
rect 12992 13942 13044 13948
rect 12992 13728 13044 13734
rect 12992 13670 13044 13676
rect 13004 13326 13032 13670
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 12900 11620 12952 11626
rect 12900 11562 12952 11568
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 13004 11218 13032 11494
rect 12992 11212 13044 11218
rect 12992 11154 13044 11160
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 12624 10736 12676 10742
rect 12624 10678 12676 10684
rect 12438 10310 12440 10362
rect 12492 10310 12494 10362
rect 12438 9274 12494 10310
rect 12438 9222 12440 9274
rect 12492 9222 12494 9274
rect 12438 8186 12494 9222
rect 12728 9042 12756 11018
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 13004 9586 13032 10610
rect 13096 10266 13124 19314
rect 13188 18850 13216 21984
rect 13280 19394 13308 31282
rect 13372 23322 13400 31758
rect 13636 31204 13688 31210
rect 13636 31146 13688 31152
rect 13452 29844 13504 29850
rect 13452 29786 13504 29792
rect 13464 29170 13492 29786
rect 13648 29238 13676 31146
rect 13636 29232 13688 29238
rect 13636 29174 13688 29180
rect 13452 29164 13504 29170
rect 13452 29106 13504 29112
rect 13740 28506 13768 33458
rect 14188 32904 14240 32910
rect 14188 32846 14240 32852
rect 14096 32768 14148 32774
rect 14096 32710 14148 32716
rect 14108 32502 14136 32710
rect 14096 32496 14148 32502
rect 14096 32438 14148 32444
rect 14200 31958 14228 32846
rect 14476 32570 14504 33934
rect 14556 33312 14608 33318
rect 14556 33254 14608 33260
rect 14568 32910 14596 33254
rect 14556 32904 14608 32910
rect 14556 32846 14608 32852
rect 14464 32564 14516 32570
rect 14464 32506 14516 32512
rect 14372 32360 14424 32366
rect 14372 32302 14424 32308
rect 14188 31952 14240 31958
rect 14188 31894 14240 31900
rect 14384 31822 14412 32302
rect 14464 32224 14516 32230
rect 14464 32166 14516 32172
rect 14372 31816 14424 31822
rect 14372 31758 14424 31764
rect 14476 31668 14504 32166
rect 14384 31640 14504 31668
rect 14280 31340 14332 31346
rect 14280 31282 14332 31288
rect 14096 31272 14148 31278
rect 14096 31214 14148 31220
rect 14108 30938 14136 31214
rect 14096 30932 14148 30938
rect 14096 30874 14148 30880
rect 14292 30870 14320 31282
rect 14280 30864 14332 30870
rect 14280 30806 14332 30812
rect 14384 30734 14412 31640
rect 14660 31482 14688 34546
rect 14924 34536 14976 34542
rect 14924 34478 14976 34484
rect 14936 34202 14964 34478
rect 14924 34196 14976 34202
rect 14924 34138 14976 34144
rect 14936 33114 14964 34138
rect 15212 33658 15240 34546
rect 15384 34400 15436 34406
rect 15384 34342 15436 34348
rect 15200 33652 15252 33658
rect 15200 33594 15252 33600
rect 14924 33108 14976 33114
rect 14924 33050 14976 33056
rect 14936 32994 14964 33050
rect 14936 32966 15148 32994
rect 14924 32904 14976 32910
rect 14924 32846 14976 32852
rect 14936 32416 14964 32846
rect 15016 32428 15068 32434
rect 14936 32388 15016 32416
rect 14832 32292 14884 32298
rect 14832 32234 14884 32240
rect 14844 31822 14872 32234
rect 14832 31816 14884 31822
rect 14832 31758 14884 31764
rect 14648 31476 14700 31482
rect 14648 31418 14700 31424
rect 14464 31136 14516 31142
rect 14464 31078 14516 31084
rect 14372 30728 14424 30734
rect 14292 30688 14372 30716
rect 13912 30592 13964 30598
rect 13912 30534 13964 30540
rect 13924 29152 13952 30534
rect 14188 29776 14240 29782
rect 14188 29718 14240 29724
rect 14096 29640 14148 29646
rect 14096 29582 14148 29588
rect 13832 29124 13952 29152
rect 13832 28642 13860 29124
rect 14108 29102 14136 29582
rect 14096 29096 14148 29102
rect 14096 29038 14148 29044
rect 13912 29028 13964 29034
rect 13912 28970 13964 28976
rect 13924 28914 13952 28970
rect 14200 28914 14228 29718
rect 13924 28886 14228 28914
rect 13832 28614 13952 28642
rect 13740 28478 13860 28506
rect 13924 28490 13952 28614
rect 13728 28416 13780 28422
rect 13728 28358 13780 28364
rect 13636 28076 13688 28082
rect 13636 28018 13688 28024
rect 13452 27940 13504 27946
rect 13504 27900 13584 27928
rect 13452 27882 13504 27888
rect 13452 27056 13504 27062
rect 13452 26998 13504 27004
rect 13360 23316 13412 23322
rect 13360 23258 13412 23264
rect 13464 22778 13492 26998
rect 13556 26450 13584 27900
rect 13648 27130 13676 28018
rect 13636 27124 13688 27130
rect 13636 27066 13688 27072
rect 13740 26994 13768 28358
rect 13832 28234 13860 28478
rect 13912 28484 13964 28490
rect 13912 28426 13964 28432
rect 13832 28206 13952 28234
rect 13924 28098 13952 28206
rect 13924 28082 14136 28098
rect 13924 28076 14148 28082
rect 13924 28070 14096 28076
rect 14096 28018 14148 28024
rect 14200 27606 14228 28886
rect 13912 27600 13964 27606
rect 13912 27542 13964 27548
rect 14188 27600 14240 27606
rect 14188 27542 14240 27548
rect 13728 26988 13780 26994
rect 13728 26930 13780 26936
rect 13924 26790 13952 27542
rect 14004 27464 14056 27470
rect 14004 27406 14056 27412
rect 14016 26994 14044 27406
rect 14004 26988 14056 26994
rect 14004 26930 14056 26936
rect 14188 26920 14240 26926
rect 14188 26862 14240 26868
rect 13912 26784 13964 26790
rect 13912 26726 13964 26732
rect 14004 26784 14056 26790
rect 14004 26726 14056 26732
rect 13544 26444 13596 26450
rect 13544 26386 13596 26392
rect 13636 26376 13688 26382
rect 13636 26318 13688 26324
rect 13820 26376 13872 26382
rect 13820 26318 13872 26324
rect 13648 25974 13676 26318
rect 13636 25968 13688 25974
rect 13636 25910 13688 25916
rect 13544 25900 13596 25906
rect 13544 25842 13596 25848
rect 13556 23254 13584 25842
rect 13636 25832 13688 25838
rect 13636 25774 13688 25780
rect 13648 25498 13676 25774
rect 13636 25492 13688 25498
rect 13636 25434 13688 25440
rect 13636 25220 13688 25226
rect 13636 25162 13688 25168
rect 13648 24818 13676 25162
rect 13636 24812 13688 24818
rect 13636 24754 13688 24760
rect 13648 24410 13676 24754
rect 13636 24404 13688 24410
rect 13636 24346 13688 24352
rect 13832 24342 13860 26318
rect 13924 25702 13952 26726
rect 14016 26518 14044 26726
rect 14004 26512 14056 26518
rect 14004 26454 14056 26460
rect 14096 26512 14148 26518
rect 14096 26454 14148 26460
rect 13912 25696 13964 25702
rect 13912 25638 13964 25644
rect 14004 25220 14056 25226
rect 13924 25180 14004 25208
rect 13820 24336 13872 24342
rect 13820 24278 13872 24284
rect 13728 24200 13780 24206
rect 13728 24142 13780 24148
rect 13544 23248 13596 23254
rect 13544 23190 13596 23196
rect 13740 23118 13768 24142
rect 13728 23112 13780 23118
rect 13728 23054 13780 23060
rect 13832 23050 13860 24278
rect 13820 23044 13872 23050
rect 13820 22986 13872 22992
rect 13544 22976 13596 22982
rect 13544 22918 13596 22924
rect 13556 22778 13584 22918
rect 13452 22772 13504 22778
rect 13452 22714 13504 22720
rect 13544 22772 13596 22778
rect 13544 22714 13596 22720
rect 13636 22160 13688 22166
rect 13636 22102 13688 22108
rect 13452 22092 13504 22098
rect 13452 22034 13504 22040
rect 13464 21554 13492 22034
rect 13452 21548 13504 21554
rect 13452 21490 13504 21496
rect 13280 19366 13492 19394
rect 13360 19304 13412 19310
rect 13360 19246 13412 19252
rect 13188 18822 13308 18850
rect 13176 18760 13228 18766
rect 13176 18702 13228 18708
rect 13188 18290 13216 18702
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 13176 16516 13228 16522
rect 13176 16458 13228 16464
rect 13188 15434 13216 16458
rect 13176 15428 13228 15434
rect 13176 15370 13228 15376
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 13188 13938 13216 14418
rect 13176 13932 13228 13938
rect 13176 13874 13228 13880
rect 13280 12850 13308 18822
rect 13372 18630 13400 19246
rect 13464 18766 13492 19366
rect 13648 19174 13676 22102
rect 13832 21962 13860 22986
rect 13820 21956 13872 21962
rect 13820 21898 13872 21904
rect 13820 21684 13872 21690
rect 13820 21626 13872 21632
rect 13728 20800 13780 20806
rect 13728 20742 13780 20748
rect 13740 19378 13768 20742
rect 13728 19372 13780 19378
rect 13728 19314 13780 19320
rect 13636 19168 13688 19174
rect 13636 19110 13688 19116
rect 13452 18760 13504 18766
rect 13452 18702 13504 18708
rect 13360 18624 13412 18630
rect 13360 18566 13412 18572
rect 13372 17746 13400 18566
rect 13648 18358 13676 19110
rect 13832 18630 13860 21626
rect 13924 18970 13952 25180
rect 14004 25162 14056 25168
rect 14108 24698 14136 26454
rect 14200 26246 14228 26862
rect 14188 26240 14240 26246
rect 14188 26182 14240 26188
rect 14016 24670 14136 24698
rect 14016 24274 14044 24670
rect 14096 24608 14148 24614
rect 14096 24550 14148 24556
rect 14188 24608 14240 24614
rect 14188 24550 14240 24556
rect 14108 24410 14136 24550
rect 14096 24404 14148 24410
rect 14096 24346 14148 24352
rect 14200 24274 14228 24550
rect 14004 24268 14056 24274
rect 14004 24210 14056 24216
rect 14188 24268 14240 24274
rect 14188 24210 14240 24216
rect 14004 24064 14056 24070
rect 14004 24006 14056 24012
rect 14016 23798 14044 24006
rect 14004 23792 14056 23798
rect 14004 23734 14056 23740
rect 14292 23662 14320 30688
rect 14372 30670 14424 30676
rect 14372 30116 14424 30122
rect 14372 30058 14424 30064
rect 14384 29102 14412 30058
rect 14372 29096 14424 29102
rect 14372 29038 14424 29044
rect 14476 28762 14504 31078
rect 14936 30802 14964 32388
rect 15016 32370 15068 32376
rect 15120 31890 15148 32966
rect 15396 32910 15424 34342
rect 15488 34202 15516 34546
rect 15476 34196 15528 34202
rect 15476 34138 15528 34144
rect 15476 33992 15528 33998
rect 15580 33980 15608 34682
rect 15672 34678 15700 35566
rect 15660 34672 15712 34678
rect 15660 34614 15712 34620
rect 15948 34474 15976 35566
rect 16040 35222 16068 35974
rect 16028 35216 16080 35222
rect 16028 35158 16080 35164
rect 16500 35034 16528 37334
rect 16592 36174 16620 38694
rect 17236 38554 17264 38898
rect 17408 38820 17460 38826
rect 17408 38762 17460 38768
rect 17224 38548 17276 38554
rect 17224 38490 17276 38496
rect 17040 38412 17092 38418
rect 17092 38372 17172 38400
rect 17040 38354 17092 38360
rect 16856 37800 16908 37806
rect 16856 37742 16908 37748
rect 16672 36780 16724 36786
rect 16672 36722 16724 36728
rect 16684 36310 16712 36722
rect 16672 36304 16724 36310
rect 16672 36246 16724 36252
rect 16580 36168 16632 36174
rect 16580 36110 16632 36116
rect 16868 35698 16896 37742
rect 16948 37120 17000 37126
rect 16948 37062 17000 37068
rect 16960 36786 16988 37062
rect 16948 36780 17000 36786
rect 16948 36722 17000 36728
rect 17040 36712 17092 36718
rect 17040 36654 17092 36660
rect 17052 36174 17080 36654
rect 16948 36168 17000 36174
rect 16948 36110 17000 36116
rect 17040 36168 17092 36174
rect 17040 36110 17092 36116
rect 16856 35692 16908 35698
rect 16856 35634 16908 35640
rect 16672 35080 16724 35086
rect 16500 35028 16672 35034
rect 16500 35022 16724 35028
rect 16396 35012 16448 35018
rect 16396 34954 16448 34960
rect 16500 35006 16712 35022
rect 16408 34542 16436 34954
rect 16500 34950 16528 35006
rect 16488 34944 16540 34950
rect 16488 34886 16540 34892
rect 16304 34536 16356 34542
rect 16304 34478 16356 34484
rect 16396 34536 16448 34542
rect 16396 34478 16448 34484
rect 15936 34468 15988 34474
rect 15936 34410 15988 34416
rect 16316 34066 16344 34478
rect 16304 34060 16356 34066
rect 16304 34002 16356 34008
rect 15528 33952 15608 33980
rect 15660 33992 15712 33998
rect 15476 33934 15528 33940
rect 15660 33934 15712 33940
rect 15936 33992 15988 33998
rect 15936 33934 15988 33940
rect 15384 32904 15436 32910
rect 15384 32846 15436 32852
rect 15384 32564 15436 32570
rect 15384 32506 15436 32512
rect 15200 32496 15252 32502
rect 15200 32438 15252 32444
rect 15212 31958 15240 32438
rect 15292 32360 15344 32366
rect 15292 32302 15344 32308
rect 15200 31952 15252 31958
rect 15200 31894 15252 31900
rect 15108 31884 15160 31890
rect 15108 31826 15160 31832
rect 15120 31754 15148 31826
rect 15028 31726 15148 31754
rect 14924 30796 14976 30802
rect 14924 30738 14976 30744
rect 14556 30388 14608 30394
rect 14556 30330 14608 30336
rect 14464 28756 14516 28762
rect 14464 28698 14516 28704
rect 14372 28552 14424 28558
rect 14372 28494 14424 28500
rect 14384 27538 14412 28494
rect 14568 27878 14596 30330
rect 14924 30320 14976 30326
rect 14924 30262 14976 30268
rect 14832 29232 14884 29238
rect 14832 29174 14884 29180
rect 14648 29096 14700 29102
rect 14648 29038 14700 29044
rect 14660 28558 14688 29038
rect 14740 29028 14792 29034
rect 14740 28970 14792 28976
rect 14648 28552 14700 28558
rect 14648 28494 14700 28500
rect 14660 28218 14688 28494
rect 14648 28212 14700 28218
rect 14648 28154 14700 28160
rect 14556 27872 14608 27878
rect 14556 27814 14608 27820
rect 14372 27532 14424 27538
rect 14372 27474 14424 27480
rect 14568 27470 14596 27814
rect 14752 27470 14780 28970
rect 14844 28762 14872 29174
rect 14832 28756 14884 28762
rect 14832 28698 14884 28704
rect 14832 28416 14884 28422
rect 14832 28358 14884 28364
rect 14556 27464 14608 27470
rect 14556 27406 14608 27412
rect 14740 27464 14792 27470
rect 14740 27406 14792 27412
rect 14372 26988 14424 26994
rect 14372 26930 14424 26936
rect 14280 23656 14332 23662
rect 14280 23598 14332 23604
rect 14384 22982 14412 26930
rect 14464 26308 14516 26314
rect 14464 26250 14516 26256
rect 14476 24818 14504 26250
rect 14568 25906 14596 27406
rect 14844 26194 14872 28358
rect 14936 26314 14964 30262
rect 15028 30122 15056 31726
rect 15212 31414 15240 31894
rect 15200 31408 15252 31414
rect 15200 31350 15252 31356
rect 15304 31346 15332 32302
rect 15292 31340 15344 31346
rect 15292 31282 15344 31288
rect 15108 30864 15160 30870
rect 15108 30806 15160 30812
rect 15016 30116 15068 30122
rect 15016 30058 15068 30064
rect 15120 30002 15148 30806
rect 15200 30728 15252 30734
rect 15200 30670 15252 30676
rect 15212 30394 15240 30670
rect 15200 30388 15252 30394
rect 15200 30330 15252 30336
rect 15028 29974 15148 30002
rect 15028 27418 15056 29974
rect 15200 29640 15252 29646
rect 15200 29582 15252 29588
rect 15212 29102 15240 29582
rect 15304 29170 15332 31282
rect 15292 29164 15344 29170
rect 15292 29106 15344 29112
rect 15200 29096 15252 29102
rect 15200 29038 15252 29044
rect 15212 28694 15240 29038
rect 15200 28688 15252 28694
rect 15200 28630 15252 28636
rect 15396 28082 15424 32506
rect 15488 32366 15516 33934
rect 15672 32502 15700 33934
rect 15752 33856 15804 33862
rect 15752 33798 15804 33804
rect 15764 33658 15792 33798
rect 15752 33652 15804 33658
rect 15752 33594 15804 33600
rect 15948 33454 15976 33934
rect 15936 33448 15988 33454
rect 15936 33390 15988 33396
rect 15948 33130 15976 33390
rect 15948 33114 16068 33130
rect 15948 33108 16080 33114
rect 15948 33102 16028 33108
rect 16028 33050 16080 33056
rect 15752 32904 15804 32910
rect 15752 32846 15804 32852
rect 16212 32904 16264 32910
rect 16212 32846 16264 32852
rect 15660 32496 15712 32502
rect 15660 32438 15712 32444
rect 15568 32428 15620 32434
rect 15568 32370 15620 32376
rect 15476 32360 15528 32366
rect 15476 32302 15528 32308
rect 15476 31680 15528 31686
rect 15476 31622 15528 31628
rect 15488 30734 15516 31622
rect 15476 30728 15528 30734
rect 15476 30670 15528 30676
rect 15476 30252 15528 30258
rect 15476 30194 15528 30200
rect 15384 28076 15436 28082
rect 15384 28018 15436 28024
rect 15292 28008 15344 28014
rect 15292 27950 15344 27956
rect 15200 27464 15252 27470
rect 15028 27402 15148 27418
rect 15200 27406 15252 27412
rect 15028 27396 15160 27402
rect 15028 27390 15108 27396
rect 14924 26308 14976 26314
rect 14924 26250 14976 26256
rect 14660 26166 14872 26194
rect 14556 25900 14608 25906
rect 14556 25842 14608 25848
rect 14464 24812 14516 24818
rect 14464 24754 14516 24760
rect 14660 23474 14688 26166
rect 14832 26036 14884 26042
rect 14832 25978 14884 25984
rect 14740 25288 14792 25294
rect 14740 25230 14792 25236
rect 14752 24274 14780 25230
rect 14740 24268 14792 24274
rect 14740 24210 14792 24216
rect 14476 23446 14688 23474
rect 14096 22976 14148 22982
rect 14096 22918 14148 22924
rect 14372 22976 14424 22982
rect 14372 22918 14424 22924
rect 14108 22710 14136 22918
rect 14096 22704 14148 22710
rect 14096 22646 14148 22652
rect 14280 22704 14332 22710
rect 14280 22646 14332 22652
rect 14096 22500 14148 22506
rect 14096 22442 14148 22448
rect 14108 21418 14136 22442
rect 14292 21486 14320 22646
rect 14384 22166 14412 22918
rect 14372 22160 14424 22166
rect 14372 22102 14424 22108
rect 14372 21888 14424 21894
rect 14372 21830 14424 21836
rect 14384 21554 14412 21830
rect 14372 21548 14424 21554
rect 14372 21490 14424 21496
rect 14280 21480 14332 21486
rect 14280 21422 14332 21428
rect 14096 21412 14148 21418
rect 14096 21354 14148 21360
rect 14188 21344 14240 21350
rect 14188 21286 14240 21292
rect 14096 20936 14148 20942
rect 14096 20878 14148 20884
rect 14004 19848 14056 19854
rect 14004 19790 14056 19796
rect 13912 18964 13964 18970
rect 13912 18906 13964 18912
rect 13820 18624 13872 18630
rect 13820 18566 13872 18572
rect 13636 18352 13688 18358
rect 13636 18294 13688 18300
rect 13820 18352 13872 18358
rect 13820 18294 13872 18300
rect 13360 17740 13412 17746
rect 13360 17682 13412 17688
rect 13832 17270 13860 18294
rect 13912 17672 13964 17678
rect 14016 17660 14044 19790
rect 14108 19786 14136 20878
rect 14200 20534 14228 21286
rect 14372 20936 14424 20942
rect 14372 20878 14424 20884
rect 14188 20528 14240 20534
rect 14188 20470 14240 20476
rect 14280 19984 14332 19990
rect 14280 19926 14332 19932
rect 14188 19916 14240 19922
rect 14188 19858 14240 19864
rect 14096 19780 14148 19786
rect 14096 19722 14148 19728
rect 14200 19718 14228 19858
rect 14188 19712 14240 19718
rect 14188 19654 14240 19660
rect 14188 18760 14240 18766
rect 14188 18702 14240 18708
rect 14200 17882 14228 18702
rect 14188 17876 14240 17882
rect 14188 17818 14240 17824
rect 13964 17632 14044 17660
rect 13912 17614 13964 17620
rect 13820 17264 13872 17270
rect 13820 17206 13872 17212
rect 13544 17128 13596 17134
rect 13544 17070 13596 17076
rect 13556 14890 13584 17070
rect 13832 16658 13860 17206
rect 13924 16998 13952 17614
rect 14096 17604 14148 17610
rect 14148 17564 14228 17592
rect 14096 17546 14148 17552
rect 14004 17536 14056 17542
rect 14004 17478 14056 17484
rect 14016 17270 14044 17478
rect 14004 17264 14056 17270
rect 14004 17206 14056 17212
rect 13912 16992 13964 16998
rect 13912 16934 13964 16940
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 13544 14884 13596 14890
rect 13544 14826 13596 14832
rect 13544 14544 13596 14550
rect 13544 14486 13596 14492
rect 13452 14340 13504 14346
rect 13452 14282 13504 14288
rect 13464 13938 13492 14282
rect 13556 13938 13584 14486
rect 13452 13932 13504 13938
rect 13452 13874 13504 13880
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13268 12844 13320 12850
rect 13268 12786 13320 12792
rect 13176 12776 13228 12782
rect 13176 12718 13228 12724
rect 13188 11898 13216 12718
rect 13360 12640 13412 12646
rect 13360 12582 13412 12588
rect 13268 12436 13320 12442
rect 13268 12378 13320 12384
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 13280 11830 13308 12378
rect 13268 11824 13320 11830
rect 13268 11766 13320 11772
rect 13372 10742 13400 12582
rect 13360 10736 13412 10742
rect 13360 10678 13412 10684
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12438 8134 12440 8186
rect 12492 8134 12494 8186
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 12360 7478 12388 7686
rect 12348 7472 12400 7478
rect 12348 7414 12400 7420
rect 12268 7262 12388 7290
rect 12256 6724 12308 6730
rect 12256 6666 12308 6672
rect 12268 6458 12296 6666
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12164 5568 12216 5574
rect 12164 5510 12216 5516
rect 12176 4622 12204 5510
rect 12164 4616 12216 4622
rect 12164 4558 12216 4564
rect 12072 2304 12124 2310
rect 12072 2246 12124 2252
rect 10048 1352 10100 1358
rect 10048 1294 10100 1300
rect 10600 1352 10652 1358
rect 10600 1294 10652 1300
rect 11704 1352 11756 1358
rect 11704 1294 11756 1300
rect 11980 1284 12032 1290
rect 11980 1226 12032 1232
rect 9680 1216 9732 1222
rect 9680 1158 9732 1164
rect 9220 876 9272 882
rect 9220 818 9272 824
rect 6276 740 6328 746
rect 6276 682 6328 688
rect 8298 0 8354 800
rect 11992 746 12020 1226
rect 12360 1222 12388 7262
rect 12438 7098 12494 8134
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 12544 7546 12572 7822
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 12438 7046 12440 7098
rect 12492 7046 12494 7098
rect 12438 6010 12494 7046
rect 12636 6254 12664 7958
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12820 6934 12848 7822
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12912 7002 12940 7142
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 12808 6928 12860 6934
rect 12808 6870 12860 6876
rect 12624 6248 12676 6254
rect 12624 6190 12676 6196
rect 12438 5958 12440 6010
rect 12492 5958 12494 6010
rect 12438 4922 12494 5958
rect 12636 5846 12664 6190
rect 12624 5840 12676 5846
rect 12624 5782 12676 5788
rect 12900 5840 12952 5846
rect 12900 5782 12952 5788
rect 12636 5250 12664 5782
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 12544 5222 12664 5250
rect 12544 5098 12572 5222
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12532 5092 12584 5098
rect 12532 5034 12584 5040
rect 12438 4870 12440 4922
rect 12492 4870 12494 4922
rect 12438 3834 12494 4870
rect 12636 4758 12664 5102
rect 12624 4752 12676 4758
rect 12624 4694 12676 4700
rect 12820 4010 12848 5646
rect 12912 5166 12940 5782
rect 12900 5160 12952 5166
rect 12900 5102 12952 5108
rect 12808 4004 12860 4010
rect 12808 3946 12860 3952
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12438 3782 12440 3834
rect 12492 3782 12494 3834
rect 12438 2746 12494 3782
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 12728 3126 12756 3674
rect 12716 3120 12768 3126
rect 12716 3062 12768 3068
rect 12912 3058 12940 3878
rect 12900 3052 12952 3058
rect 12438 2694 12440 2746
rect 12492 2694 12494 2746
rect 12438 1658 12494 2694
rect 12820 3012 12900 3040
rect 12820 2514 12848 3012
rect 12900 2994 12952 3000
rect 13004 2774 13032 9522
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 13096 9110 13124 9318
rect 13084 9104 13136 9110
rect 13084 9046 13136 9052
rect 13360 8288 13412 8294
rect 13464 8242 13492 13874
rect 13544 13728 13596 13734
rect 13544 13670 13596 13676
rect 13556 12238 13584 13670
rect 13648 12306 13676 16050
rect 13832 15706 13860 16594
rect 13820 15700 13872 15706
rect 13820 15642 13872 15648
rect 13832 15026 13860 15642
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13832 14414 13860 14962
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13740 12442 13768 14214
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13636 12300 13688 12306
rect 13636 12242 13688 12248
rect 13832 12238 13860 14350
rect 13924 13870 13952 16934
rect 14004 15564 14056 15570
rect 14004 15506 14056 15512
rect 14016 14618 14044 15506
rect 14200 15502 14228 17564
rect 14188 15496 14240 15502
rect 14188 15438 14240 15444
rect 14188 15360 14240 15366
rect 14188 15302 14240 15308
rect 14096 15156 14148 15162
rect 14096 15098 14148 15104
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 13912 13864 13964 13870
rect 13912 13806 13964 13812
rect 13912 13252 13964 13258
rect 13912 13194 13964 13200
rect 13924 12850 13952 13194
rect 14108 12850 14136 15098
rect 14200 14618 14228 15302
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 14188 13320 14240 13326
rect 14188 13262 14240 13268
rect 14200 12986 14228 13262
rect 14188 12980 14240 12986
rect 14188 12922 14240 12928
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 13544 12232 13596 12238
rect 13544 12174 13596 12180
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 14292 11778 14320 19926
rect 14384 19854 14412 20878
rect 14476 19854 14504 23446
rect 14648 23248 14700 23254
rect 14648 23190 14700 23196
rect 14556 22024 14608 22030
rect 14556 21966 14608 21972
rect 14568 20534 14596 21966
rect 14660 21962 14688 23190
rect 14752 23118 14780 24210
rect 14740 23112 14792 23118
rect 14740 23054 14792 23060
rect 14648 21956 14700 21962
rect 14648 21898 14700 21904
rect 14844 21842 14872 25978
rect 14924 25696 14976 25702
rect 14924 25638 14976 25644
rect 14936 24886 14964 25638
rect 14924 24880 14976 24886
rect 14924 24822 14976 24828
rect 14924 24608 14976 24614
rect 14924 24550 14976 24556
rect 14936 24206 14964 24550
rect 14924 24200 14976 24206
rect 14924 24142 14976 24148
rect 14924 24064 14976 24070
rect 14924 24006 14976 24012
rect 14936 23798 14964 24006
rect 14924 23792 14976 23798
rect 14924 23734 14976 23740
rect 14924 23316 14976 23322
rect 14924 23258 14976 23264
rect 14936 22166 14964 23258
rect 14924 22160 14976 22166
rect 14924 22102 14976 22108
rect 14660 21814 14872 21842
rect 14660 21622 14688 21814
rect 15028 21672 15056 27390
rect 15108 27338 15160 27344
rect 15212 26364 15240 27406
rect 15304 27062 15332 27950
rect 15292 27056 15344 27062
rect 15292 26998 15344 27004
rect 15396 26994 15424 28018
rect 15384 26988 15436 26994
rect 15384 26930 15436 26936
rect 15488 26518 15516 30194
rect 15476 26512 15528 26518
rect 15476 26454 15528 26460
rect 15292 26376 15344 26382
rect 15212 26336 15292 26364
rect 15292 26318 15344 26324
rect 15200 25900 15252 25906
rect 15200 25842 15252 25848
rect 15212 25498 15240 25842
rect 15200 25492 15252 25498
rect 15200 25434 15252 25440
rect 15108 25424 15160 25430
rect 15108 25366 15160 25372
rect 15120 24342 15148 25366
rect 15304 25362 15332 26318
rect 15384 26308 15436 26314
rect 15384 26250 15436 26256
rect 15292 25356 15344 25362
rect 15292 25298 15344 25304
rect 15108 24336 15160 24342
rect 15108 24278 15160 24284
rect 15108 24200 15160 24206
rect 15108 24142 15160 24148
rect 15120 22778 15148 24142
rect 15200 23248 15252 23254
rect 15200 23190 15252 23196
rect 15108 22772 15160 22778
rect 15108 22714 15160 22720
rect 15108 22432 15160 22438
rect 15108 22374 15160 22380
rect 15120 22030 15148 22374
rect 15108 22024 15160 22030
rect 15108 21966 15160 21972
rect 14752 21644 15056 21672
rect 14648 21616 14700 21622
rect 14648 21558 14700 21564
rect 14556 20528 14608 20534
rect 14556 20470 14608 20476
rect 14648 20392 14700 20398
rect 14648 20334 14700 20340
rect 14372 19848 14424 19854
rect 14372 19790 14424 19796
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 14476 19700 14504 19790
rect 14384 19672 14504 19700
rect 14384 16250 14412 19672
rect 14464 19372 14516 19378
rect 14464 19314 14516 19320
rect 14476 18426 14504 19314
rect 14660 19310 14688 20334
rect 14752 20262 14780 21644
rect 14832 21548 14884 21554
rect 14832 21490 14884 21496
rect 14740 20256 14792 20262
rect 14740 20198 14792 20204
rect 14740 19712 14792 19718
rect 14740 19654 14792 19660
rect 14648 19304 14700 19310
rect 14648 19246 14700 19252
rect 14464 18420 14516 18426
rect 14464 18362 14516 18368
rect 14476 17678 14504 18362
rect 14464 17672 14516 17678
rect 14464 17614 14516 17620
rect 14752 17202 14780 19654
rect 14844 19514 14872 21490
rect 14924 21480 14976 21486
rect 14924 21422 14976 21428
rect 15108 21480 15160 21486
rect 15108 21422 15160 21428
rect 14936 20806 14964 21422
rect 15016 20936 15068 20942
rect 15120 20924 15148 21422
rect 15068 20896 15148 20924
rect 15016 20878 15068 20884
rect 14924 20800 14976 20806
rect 14924 20742 14976 20748
rect 14936 20466 14964 20742
rect 15108 20528 15160 20534
rect 15108 20470 15160 20476
rect 14924 20460 14976 20466
rect 14924 20402 14976 20408
rect 14924 19848 14976 19854
rect 14924 19790 14976 19796
rect 14832 19508 14884 19514
rect 14832 19450 14884 19456
rect 14832 18216 14884 18222
rect 14832 18158 14884 18164
rect 14844 17610 14872 18158
rect 14832 17604 14884 17610
rect 14832 17546 14884 17552
rect 14740 17196 14792 17202
rect 14740 17138 14792 17144
rect 14372 16244 14424 16250
rect 14372 16186 14424 16192
rect 14372 16040 14424 16046
rect 14372 15982 14424 15988
rect 14200 11750 14320 11778
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13648 11286 13676 11494
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13636 11280 13688 11286
rect 13636 11222 13688 11228
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13412 8236 13492 8242
rect 13360 8230 13492 8236
rect 13372 8214 13492 8230
rect 13464 8090 13492 8214
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13556 7750 13584 8978
rect 13636 8832 13688 8838
rect 13636 8774 13688 8780
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13452 7200 13504 7206
rect 13452 7142 13504 7148
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 13096 6458 13124 6734
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 13464 6322 13492 7142
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 13544 5772 13596 5778
rect 13544 5714 13596 5720
rect 13084 5704 13136 5710
rect 13084 5646 13136 5652
rect 13096 4214 13124 5646
rect 13176 5636 13228 5642
rect 13176 5578 13228 5584
rect 13084 4208 13136 4214
rect 13084 4150 13136 4156
rect 12912 2746 13032 2774
rect 12808 2508 12860 2514
rect 12808 2450 12860 2456
rect 12912 1834 12940 2746
rect 13096 2650 13124 4150
rect 13188 3602 13216 5578
rect 13556 4622 13584 5714
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 13544 4480 13596 4486
rect 13544 4422 13596 4428
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 13176 3596 13228 3602
rect 13176 3538 13228 3544
rect 13084 2644 13136 2650
rect 13084 2586 13136 2592
rect 13084 2372 13136 2378
rect 13084 2314 13136 2320
rect 12900 1828 12952 1834
rect 12900 1770 12952 1776
rect 12438 1606 12440 1658
rect 12492 1606 12494 1658
rect 12348 1216 12400 1222
rect 12348 1158 12400 1164
rect 12438 1040 12494 1606
rect 13096 1562 13124 2314
rect 13084 1556 13136 1562
rect 13084 1498 13136 1504
rect 13280 1358 13308 3878
rect 13556 3534 13584 4422
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13544 3392 13596 3398
rect 13544 3334 13596 3340
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 13372 2038 13400 2994
rect 13360 2032 13412 2038
rect 13360 1974 13412 1980
rect 13556 1970 13584 3334
rect 13544 1964 13596 1970
rect 13544 1906 13596 1912
rect 13544 1760 13596 1766
rect 13544 1702 13596 1708
rect 13556 1562 13584 1702
rect 13544 1556 13596 1562
rect 13544 1498 13596 1504
rect 13648 1358 13676 8774
rect 13268 1352 13320 1358
rect 13268 1294 13320 1300
rect 13636 1352 13688 1358
rect 13636 1294 13688 1300
rect 13740 1222 13768 11290
rect 14096 11144 14148 11150
rect 14096 11086 14148 11092
rect 14108 9926 14136 11086
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 13924 8838 13952 9590
rect 14108 9586 14136 9862
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14004 9444 14056 9450
rect 14004 9386 14056 9392
rect 14016 9178 14044 9386
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 14108 9042 14136 9522
rect 14096 9036 14148 9042
rect 14096 8978 14148 8984
rect 13912 8832 13964 8838
rect 13912 8774 13964 8780
rect 14108 8566 14136 8978
rect 14096 8560 14148 8566
rect 14096 8502 14148 8508
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 14004 7472 14056 7478
rect 14004 7414 14056 7420
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13832 7274 13860 7346
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 13832 6322 13860 7210
rect 14016 6322 14044 7414
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13832 5166 13860 6054
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 13832 3738 13860 5102
rect 14004 5092 14056 5098
rect 14004 5034 14056 5040
rect 14016 4282 14044 5034
rect 14108 4622 14136 7822
rect 14200 6458 14228 11750
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14292 10538 14320 11630
rect 14280 10532 14332 10538
rect 14280 10474 14332 10480
rect 14384 10418 14412 15982
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 14292 10390 14412 10418
rect 14292 10130 14320 10390
rect 14280 10124 14332 10130
rect 14280 10066 14332 10072
rect 14292 7886 14320 10066
rect 14476 9994 14504 15438
rect 14648 15020 14700 15026
rect 14648 14962 14700 14968
rect 14660 14074 14688 14962
rect 14752 14822 14780 17138
rect 14832 16448 14884 16454
rect 14832 16390 14884 16396
rect 14844 16182 14872 16390
rect 14832 16176 14884 16182
rect 14832 16118 14884 16124
rect 14832 15904 14884 15910
rect 14832 15846 14884 15852
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14752 14414 14780 14758
rect 14740 14408 14792 14414
rect 14740 14350 14792 14356
rect 14648 14068 14700 14074
rect 14648 14010 14700 14016
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 14648 13932 14700 13938
rect 14752 13920 14780 14010
rect 14844 13938 14872 15846
rect 14936 15162 14964 19790
rect 15120 19786 15148 20470
rect 15108 19780 15160 19786
rect 15108 19722 15160 19728
rect 15016 19236 15068 19242
rect 15016 19178 15068 19184
rect 15028 18426 15056 19178
rect 15120 18766 15148 19722
rect 15108 18760 15160 18766
rect 15108 18702 15160 18708
rect 15016 18420 15068 18426
rect 15016 18362 15068 18368
rect 15016 17672 15068 17678
rect 15016 17614 15068 17620
rect 15028 17202 15056 17614
rect 15120 17542 15148 18702
rect 15108 17536 15160 17542
rect 15108 17478 15160 17484
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 15028 16114 15056 17138
rect 15108 16652 15160 16658
rect 15108 16594 15160 16600
rect 15120 16522 15148 16594
rect 15108 16516 15160 16522
rect 15108 16458 15160 16464
rect 15016 16108 15068 16114
rect 15016 16050 15068 16056
rect 14924 15156 14976 15162
rect 14924 15098 14976 15104
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 14700 13892 14780 13920
rect 14832 13932 14884 13938
rect 14648 13874 14700 13880
rect 14832 13874 14884 13880
rect 14648 13320 14700 13326
rect 14648 13262 14700 13268
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14568 12102 14596 12786
rect 14556 12096 14608 12102
rect 14556 12038 14608 12044
rect 14660 10674 14688 13262
rect 14936 13258 14964 14758
rect 15028 14414 15056 16050
rect 15212 15178 15240 23190
rect 15304 22642 15332 25298
rect 15396 25294 15424 26250
rect 15384 25288 15436 25294
rect 15384 25230 15436 25236
rect 15476 24880 15528 24886
rect 15476 24822 15528 24828
rect 15384 23860 15436 23866
rect 15384 23802 15436 23808
rect 15292 22636 15344 22642
rect 15292 22578 15344 22584
rect 15304 22438 15332 22578
rect 15292 22432 15344 22438
rect 15292 22374 15344 22380
rect 15292 22160 15344 22166
rect 15292 22102 15344 22108
rect 15304 21962 15332 22102
rect 15292 21956 15344 21962
rect 15292 21898 15344 21904
rect 15304 19854 15332 21898
rect 15396 20874 15424 23802
rect 15488 22642 15516 24822
rect 15476 22636 15528 22642
rect 15476 22578 15528 22584
rect 15488 22030 15516 22578
rect 15580 22438 15608 32370
rect 15660 31816 15712 31822
rect 15660 31758 15712 31764
rect 15672 31482 15700 31758
rect 15660 31476 15712 31482
rect 15660 31418 15712 31424
rect 15660 31340 15712 31346
rect 15660 31282 15712 31288
rect 15672 29646 15700 31282
rect 15660 29640 15712 29646
rect 15660 29582 15712 29588
rect 15672 29238 15700 29582
rect 15660 29232 15712 29238
rect 15660 29174 15712 29180
rect 15764 28762 15792 32846
rect 16120 32836 16172 32842
rect 16120 32778 16172 32784
rect 16132 32570 16160 32778
rect 16120 32564 16172 32570
rect 16120 32506 16172 32512
rect 16028 31884 16080 31890
rect 16028 31826 16080 31832
rect 15936 31340 15988 31346
rect 15936 31282 15988 31288
rect 15948 30938 15976 31282
rect 15936 30932 15988 30938
rect 15936 30874 15988 30880
rect 15752 28756 15804 28762
rect 15752 28698 15804 28704
rect 15752 28552 15804 28558
rect 15752 28494 15804 28500
rect 15764 27674 15792 28494
rect 15752 27668 15804 27674
rect 15752 27610 15804 27616
rect 15660 26376 15712 26382
rect 15660 26318 15712 26324
rect 15844 26376 15896 26382
rect 15844 26318 15896 26324
rect 15672 24886 15700 26318
rect 15856 25702 15884 26318
rect 15844 25696 15896 25702
rect 15844 25638 15896 25644
rect 15752 25220 15804 25226
rect 15752 25162 15804 25168
rect 15660 24880 15712 24886
rect 15660 24822 15712 24828
rect 15660 24336 15712 24342
rect 15660 24278 15712 24284
rect 15568 22432 15620 22438
rect 15568 22374 15620 22380
rect 15580 22234 15608 22374
rect 15568 22228 15620 22234
rect 15568 22170 15620 22176
rect 15476 22024 15528 22030
rect 15476 21966 15528 21972
rect 15568 22024 15620 22030
rect 15568 21966 15620 21972
rect 15476 21888 15528 21894
rect 15476 21830 15528 21836
rect 15384 20868 15436 20874
rect 15384 20810 15436 20816
rect 15488 20534 15516 21830
rect 15476 20528 15528 20534
rect 15476 20470 15528 20476
rect 15384 20460 15436 20466
rect 15384 20402 15436 20408
rect 15292 19848 15344 19854
rect 15292 19790 15344 19796
rect 15396 19378 15424 20402
rect 15580 20330 15608 21966
rect 15672 21486 15700 24278
rect 15764 23798 15792 25162
rect 15856 24206 15884 25638
rect 16040 25430 16068 31826
rect 16120 31748 16172 31754
rect 16120 31690 16172 31696
rect 16132 31482 16160 31690
rect 16120 31476 16172 31482
rect 16120 31418 16172 31424
rect 16120 30184 16172 30190
rect 16120 30126 16172 30132
rect 16132 29578 16160 30126
rect 16120 29572 16172 29578
rect 16120 29514 16172 29520
rect 16224 28218 16252 32846
rect 16316 32298 16344 34002
rect 16488 33992 16540 33998
rect 16488 33934 16540 33940
rect 16396 32768 16448 32774
rect 16396 32710 16448 32716
rect 16304 32292 16356 32298
rect 16304 32234 16356 32240
rect 16316 31346 16344 32234
rect 16304 31340 16356 31346
rect 16304 31282 16356 31288
rect 16304 30048 16356 30054
rect 16304 29990 16356 29996
rect 16316 29578 16344 29990
rect 16304 29572 16356 29578
rect 16304 29514 16356 29520
rect 16304 28552 16356 28558
rect 16304 28494 16356 28500
rect 16212 28212 16264 28218
rect 16212 28154 16264 28160
rect 16120 28008 16172 28014
rect 16120 27950 16172 27956
rect 16132 25974 16160 27950
rect 16316 27878 16344 28494
rect 16304 27872 16356 27878
rect 16304 27814 16356 27820
rect 16212 26988 16264 26994
rect 16212 26930 16264 26936
rect 16120 25968 16172 25974
rect 16120 25910 16172 25916
rect 16028 25424 16080 25430
rect 16028 25366 16080 25372
rect 16028 24744 16080 24750
rect 16028 24686 16080 24692
rect 15936 24676 15988 24682
rect 15936 24618 15988 24624
rect 15948 24206 15976 24618
rect 15844 24200 15896 24206
rect 15844 24142 15896 24148
rect 15936 24200 15988 24206
rect 15936 24142 15988 24148
rect 15752 23792 15804 23798
rect 15752 23734 15804 23740
rect 15856 23730 15884 24142
rect 15844 23724 15896 23730
rect 15844 23666 15896 23672
rect 15752 23520 15804 23526
rect 15752 23462 15804 23468
rect 15844 23520 15896 23526
rect 15844 23462 15896 23468
rect 15764 23050 15792 23462
rect 15752 23044 15804 23050
rect 15752 22986 15804 22992
rect 15764 22642 15792 22986
rect 15856 22982 15884 23462
rect 15844 22976 15896 22982
rect 15844 22918 15896 22924
rect 15752 22636 15804 22642
rect 15752 22578 15804 22584
rect 15764 21554 15792 22578
rect 15936 22228 15988 22234
rect 15936 22170 15988 22176
rect 15844 21616 15896 21622
rect 15844 21558 15896 21564
rect 15752 21548 15804 21554
rect 15752 21490 15804 21496
rect 15660 21480 15712 21486
rect 15660 21422 15712 21428
rect 15660 21344 15712 21350
rect 15660 21286 15712 21292
rect 15672 20466 15700 21286
rect 15752 20868 15804 20874
rect 15752 20810 15804 20816
rect 15660 20460 15712 20466
rect 15660 20402 15712 20408
rect 15568 20324 15620 20330
rect 15568 20266 15620 20272
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 15488 19854 15516 20198
rect 15672 20058 15700 20402
rect 15660 20052 15712 20058
rect 15660 19994 15712 20000
rect 15476 19848 15528 19854
rect 15476 19790 15528 19796
rect 15568 19712 15620 19718
rect 15568 19654 15620 19660
rect 15580 19514 15608 19654
rect 15764 19514 15792 20810
rect 15568 19508 15620 19514
rect 15568 19450 15620 19456
rect 15752 19508 15804 19514
rect 15752 19450 15804 19456
rect 15384 19372 15436 19378
rect 15384 19314 15436 19320
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 15304 18748 15332 19246
rect 15568 19168 15620 19174
rect 15568 19110 15620 19116
rect 15384 18760 15436 18766
rect 15304 18720 15384 18748
rect 15384 18702 15436 18708
rect 15396 17610 15424 18702
rect 15476 18080 15528 18086
rect 15476 18022 15528 18028
rect 15488 17678 15516 18022
rect 15476 17672 15528 17678
rect 15476 17614 15528 17620
rect 15384 17604 15436 17610
rect 15384 17546 15436 17552
rect 15384 17264 15436 17270
rect 15384 17206 15436 17212
rect 15396 16658 15424 17206
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 15384 16652 15436 16658
rect 15384 16594 15436 16600
rect 15304 16182 15332 16594
rect 15396 16454 15424 16594
rect 15488 16590 15516 16934
rect 15476 16584 15528 16590
rect 15476 16526 15528 16532
rect 15580 16538 15608 19110
rect 15764 17066 15792 19450
rect 15856 18086 15884 21558
rect 15948 20942 15976 22170
rect 15936 20936 15988 20942
rect 15936 20878 15988 20884
rect 16040 20466 16068 24686
rect 16132 22098 16160 25910
rect 16224 24886 16252 26930
rect 16304 25900 16356 25906
rect 16304 25842 16356 25848
rect 16316 25226 16344 25842
rect 16408 25362 16436 32710
rect 16500 26926 16528 33934
rect 16580 33924 16632 33930
rect 16580 33866 16632 33872
rect 16592 31822 16620 33866
rect 16868 33522 16896 35634
rect 16960 35290 16988 36110
rect 16948 35284 17000 35290
rect 16948 35226 17000 35232
rect 16672 33516 16724 33522
rect 16672 33458 16724 33464
rect 16856 33516 16908 33522
rect 16856 33458 16908 33464
rect 16684 32570 16712 33458
rect 17052 33046 17080 36110
rect 17144 35086 17172 38372
rect 17420 38196 17448 38762
rect 17512 38350 17540 39442
rect 17590 39194 17646 40230
rect 17590 39142 17592 39194
rect 17644 39142 17646 39194
rect 17500 38344 17552 38350
rect 17500 38286 17552 38292
rect 17328 38168 17448 38196
rect 17328 37194 17356 38168
rect 17590 38106 17646 39142
rect 18064 39030 18092 40462
rect 18156 39642 18184 42162
rect 19340 42152 19392 42158
rect 19340 42094 19392 42100
rect 18604 42084 18656 42090
rect 18604 42026 18656 42032
rect 18236 41608 18288 41614
rect 18236 41550 18288 41556
rect 18512 41608 18564 41614
rect 18512 41550 18564 41556
rect 18248 40594 18276 41550
rect 18328 41200 18380 41206
rect 18328 41142 18380 41148
rect 18236 40588 18288 40594
rect 18236 40530 18288 40536
rect 18248 40186 18276 40530
rect 18236 40180 18288 40186
rect 18236 40122 18288 40128
rect 18144 39636 18196 39642
rect 18144 39578 18196 39584
rect 18248 39438 18276 40122
rect 18236 39432 18288 39438
rect 18236 39374 18288 39380
rect 18052 39024 18104 39030
rect 18052 38966 18104 38972
rect 18340 38962 18368 41142
rect 18524 40458 18552 41550
rect 18616 41206 18644 42026
rect 19064 42016 19116 42022
rect 19064 41958 19116 41964
rect 19076 41818 19104 41958
rect 19064 41812 19116 41818
rect 19064 41754 19116 41760
rect 18604 41200 18656 41206
rect 18604 41142 18656 41148
rect 18512 40452 18564 40458
rect 18512 40394 18564 40400
rect 18524 40050 18552 40394
rect 18512 40044 18564 40050
rect 18512 39986 18564 39992
rect 18420 39976 18472 39982
rect 18420 39918 18472 39924
rect 18432 39506 18460 39918
rect 18420 39500 18472 39506
rect 18420 39442 18472 39448
rect 18524 39438 18552 39986
rect 18512 39432 18564 39438
rect 18512 39374 18564 39380
rect 18328 38956 18380 38962
rect 18328 38898 18380 38904
rect 18880 38956 18932 38962
rect 18880 38898 18932 38904
rect 18512 38752 18564 38758
rect 18512 38694 18564 38700
rect 18524 38418 18552 38694
rect 18512 38412 18564 38418
rect 18512 38354 18564 38360
rect 17684 38344 17736 38350
rect 17684 38286 17736 38292
rect 17776 38344 17828 38350
rect 17776 38286 17828 38292
rect 17590 38054 17592 38106
rect 17644 38054 17646 38106
rect 17316 37188 17368 37194
rect 17316 37130 17368 37136
rect 17132 35080 17184 35086
rect 17132 35022 17184 35028
rect 17328 34474 17356 37130
rect 17590 37018 17646 38054
rect 17696 37126 17724 38286
rect 17788 37262 17816 38286
rect 18236 38208 18288 38214
rect 18236 38150 18288 38156
rect 18248 37942 18276 38150
rect 18236 37936 18288 37942
rect 18236 37878 18288 37884
rect 18052 37664 18104 37670
rect 18052 37606 18104 37612
rect 18420 37664 18472 37670
rect 18420 37606 18472 37612
rect 17776 37256 17828 37262
rect 17776 37198 17828 37204
rect 17868 37256 17920 37262
rect 17868 37198 17920 37204
rect 17684 37120 17736 37126
rect 17684 37062 17736 37068
rect 17590 36966 17592 37018
rect 17644 36966 17646 37018
rect 17500 36712 17552 36718
rect 17500 36654 17552 36660
rect 17408 36576 17460 36582
rect 17408 36518 17460 36524
rect 17420 35698 17448 36518
rect 17512 36242 17540 36654
rect 17500 36236 17552 36242
rect 17500 36178 17552 36184
rect 17590 35930 17646 36966
rect 17880 36904 17908 37198
rect 17696 36876 17908 36904
rect 17696 36650 17724 36876
rect 17776 36780 17828 36786
rect 17776 36722 17828 36728
rect 17684 36644 17736 36650
rect 17684 36586 17736 36592
rect 17788 36310 17816 36722
rect 17776 36304 17828 36310
rect 17776 36246 17828 36252
rect 17880 36174 17908 36876
rect 18064 36718 18092 37606
rect 18432 37262 18460 37606
rect 18236 37256 18288 37262
rect 18236 37198 18288 37204
rect 18420 37256 18472 37262
rect 18420 37198 18472 37204
rect 18248 36718 18276 37198
rect 18524 36922 18552 38354
rect 18892 38010 18920 38898
rect 19076 38554 19104 41754
rect 19352 41546 19380 42094
rect 19432 41744 19484 41750
rect 19432 41686 19484 41692
rect 19340 41540 19392 41546
rect 19340 41482 19392 41488
rect 19156 41472 19208 41478
rect 19352 41426 19380 41482
rect 19156 41414 19208 41420
rect 19168 40526 19196 41414
rect 19260 41398 19380 41426
rect 19260 41138 19288 41398
rect 19248 41132 19300 41138
rect 19248 41074 19300 41080
rect 19260 40594 19288 41074
rect 19248 40588 19300 40594
rect 19248 40530 19300 40536
rect 19156 40520 19208 40526
rect 19156 40462 19208 40468
rect 19444 40390 19472 41686
rect 19524 41676 19576 41682
rect 19524 41618 19576 41624
rect 19536 40934 19564 41618
rect 19800 40996 19852 41002
rect 19800 40938 19852 40944
rect 19524 40928 19576 40934
rect 19524 40870 19576 40876
rect 19432 40384 19484 40390
rect 19432 40326 19484 40332
rect 19444 39522 19472 40326
rect 19352 39494 19472 39522
rect 19064 38548 19116 38554
rect 19116 38508 19196 38536
rect 19064 38490 19116 38496
rect 18880 38004 18932 38010
rect 18880 37946 18932 37952
rect 19064 37868 19116 37874
rect 19064 37810 19116 37816
rect 19076 36922 19104 37810
rect 19168 37806 19196 38508
rect 19352 38486 19380 39494
rect 19432 39432 19484 39438
rect 19432 39374 19484 39380
rect 19444 39098 19472 39374
rect 19536 39370 19564 40870
rect 19708 39976 19760 39982
rect 19708 39918 19760 39924
rect 19524 39364 19576 39370
rect 19524 39306 19576 39312
rect 19432 39092 19484 39098
rect 19432 39034 19484 39040
rect 19340 38480 19392 38486
rect 19340 38422 19392 38428
rect 19352 37874 19380 38422
rect 19616 38344 19668 38350
rect 19616 38286 19668 38292
rect 19628 37874 19656 38286
rect 19340 37868 19392 37874
rect 19340 37810 19392 37816
rect 19616 37868 19668 37874
rect 19616 37810 19668 37816
rect 19156 37800 19208 37806
rect 19156 37742 19208 37748
rect 19168 37398 19196 37742
rect 19156 37392 19208 37398
rect 19156 37334 19208 37340
rect 18512 36916 18564 36922
rect 18512 36858 18564 36864
rect 19064 36916 19116 36922
rect 19064 36858 19116 36864
rect 18052 36712 18104 36718
rect 18052 36654 18104 36660
rect 18236 36712 18288 36718
rect 18236 36654 18288 36660
rect 18248 36174 18276 36654
rect 19168 36582 19196 37334
rect 19720 37330 19748 39918
rect 19708 37324 19760 37330
rect 19708 37266 19760 37272
rect 19248 36780 19300 36786
rect 19248 36722 19300 36728
rect 19524 36780 19576 36786
rect 19524 36722 19576 36728
rect 19260 36650 19288 36722
rect 19248 36644 19300 36650
rect 19248 36586 19300 36592
rect 19156 36576 19208 36582
rect 19156 36518 19208 36524
rect 19536 36242 19564 36722
rect 19720 36582 19748 37266
rect 19708 36576 19760 36582
rect 19708 36518 19760 36524
rect 19524 36236 19576 36242
rect 19524 36178 19576 36184
rect 17868 36168 17920 36174
rect 17868 36110 17920 36116
rect 18236 36168 18288 36174
rect 18236 36110 18288 36116
rect 18328 36168 18380 36174
rect 19720 36122 19748 36518
rect 18328 36110 18380 36116
rect 17590 35878 17592 35930
rect 17644 35878 17646 35930
rect 17408 35692 17460 35698
rect 17408 35634 17460 35640
rect 17500 35012 17552 35018
rect 17500 34954 17552 34960
rect 17512 34610 17540 34954
rect 17590 34842 17646 35878
rect 17880 35290 17908 36110
rect 18340 35986 18368 36110
rect 19444 36094 19748 36122
rect 18248 35958 18368 35986
rect 19156 36032 19208 36038
rect 19156 35974 19208 35980
rect 18248 35494 18276 35958
rect 18236 35488 18288 35494
rect 18236 35430 18288 35436
rect 18696 35488 18748 35494
rect 18696 35430 18748 35436
rect 17868 35284 17920 35290
rect 17868 35226 17920 35232
rect 17960 35080 18012 35086
rect 17960 35022 18012 35028
rect 17590 34790 17592 34842
rect 17644 34790 17646 34842
rect 17500 34604 17552 34610
rect 17500 34546 17552 34552
rect 17316 34468 17368 34474
rect 17316 34410 17368 34416
rect 17040 33040 17092 33046
rect 17040 32982 17092 32988
rect 17224 32768 17276 32774
rect 17224 32710 17276 32716
rect 16672 32564 16724 32570
rect 16672 32506 16724 32512
rect 17040 32428 17092 32434
rect 17040 32370 17092 32376
rect 16948 32360 17000 32366
rect 16948 32302 17000 32308
rect 16960 31890 16988 32302
rect 16948 31884 17000 31890
rect 16948 31826 17000 31832
rect 16580 31816 16632 31822
rect 16580 31758 16632 31764
rect 16592 30258 16620 31758
rect 17052 31754 17080 32370
rect 17132 32360 17184 32366
rect 17132 32302 17184 32308
rect 16776 31726 17080 31754
rect 16672 31136 16724 31142
rect 16672 31078 16724 31084
rect 16684 30666 16712 31078
rect 16672 30660 16724 30666
rect 16672 30602 16724 30608
rect 16580 30252 16632 30258
rect 16580 30194 16632 30200
rect 16580 29844 16632 29850
rect 16580 29786 16632 29792
rect 16488 26920 16540 26926
rect 16488 26862 16540 26868
rect 16592 26858 16620 29786
rect 16672 29164 16724 29170
rect 16672 29106 16724 29112
rect 16684 28472 16712 29106
rect 16776 28948 16804 31726
rect 17040 31680 17092 31686
rect 17040 31622 17092 31628
rect 16856 31340 16908 31346
rect 16856 31282 16908 31288
rect 16868 30394 16896 31282
rect 17052 31142 17080 31622
rect 17040 31136 17092 31142
rect 17040 31078 17092 31084
rect 16948 30592 17000 30598
rect 16948 30534 17000 30540
rect 16856 30388 16908 30394
rect 16856 30330 16908 30336
rect 16960 28994 16988 30534
rect 17052 29850 17080 31078
rect 17040 29844 17092 29850
rect 17040 29786 17092 29792
rect 17052 29102 17080 29786
rect 17144 29306 17172 32302
rect 17236 31958 17264 32710
rect 17224 31952 17276 31958
rect 17224 31894 17276 31900
rect 17328 31754 17356 34410
rect 17236 31726 17356 31754
rect 17590 33754 17646 34790
rect 17972 34610 18000 35022
rect 18248 34950 18276 35430
rect 18708 35222 18736 35430
rect 18696 35216 18748 35222
rect 18696 35158 18748 35164
rect 19168 35170 19196 35974
rect 19248 35692 19300 35698
rect 19248 35634 19300 35640
rect 19260 35290 19288 35634
rect 19248 35284 19300 35290
rect 19248 35226 19300 35232
rect 19340 35284 19392 35290
rect 19340 35226 19392 35232
rect 19352 35170 19380 35226
rect 19444 35222 19472 36094
rect 19524 36032 19576 36038
rect 19524 35974 19576 35980
rect 18236 34944 18288 34950
rect 18236 34886 18288 34892
rect 17960 34604 18012 34610
rect 17960 34546 18012 34552
rect 18328 34604 18380 34610
rect 18328 34546 18380 34552
rect 18512 34604 18564 34610
rect 18512 34546 18564 34552
rect 18340 33844 18368 34546
rect 18420 34400 18472 34406
rect 18420 34342 18472 34348
rect 18432 33998 18460 34342
rect 18524 34134 18552 34546
rect 18512 34128 18564 34134
rect 18512 34070 18564 34076
rect 18420 33992 18472 33998
rect 18420 33934 18472 33940
rect 18340 33816 18460 33844
rect 17590 33702 17592 33754
rect 17644 33702 17646 33754
rect 17590 32666 17646 33702
rect 18432 33658 18460 33816
rect 18524 33658 18552 34070
rect 18708 34066 18736 35158
rect 19168 35142 19380 35170
rect 19432 35216 19484 35222
rect 19432 35158 19484 35164
rect 19536 35086 19564 35974
rect 18880 35080 18932 35086
rect 18880 35022 18932 35028
rect 19524 35080 19576 35086
rect 19524 35022 19576 35028
rect 18696 34060 18748 34066
rect 18696 34002 18748 34008
rect 18788 33856 18840 33862
rect 18788 33798 18840 33804
rect 18420 33652 18472 33658
rect 18420 33594 18472 33600
rect 18512 33652 18564 33658
rect 18512 33594 18564 33600
rect 17868 33516 17920 33522
rect 17868 33458 17920 33464
rect 17590 32614 17592 32666
rect 17644 32614 17646 32666
rect 17132 29300 17184 29306
rect 17132 29242 17184 29248
rect 17040 29096 17092 29102
rect 17040 29038 17092 29044
rect 17132 29028 17184 29034
rect 16960 28966 17080 28994
rect 17132 28970 17184 28976
rect 16776 28920 16896 28948
rect 16868 28914 16896 28920
rect 16868 28886 16988 28914
rect 16764 28484 16816 28490
rect 16684 28444 16764 28472
rect 16764 28426 16816 28432
rect 16960 28200 16988 28886
rect 16776 28172 16988 28200
rect 16580 26852 16632 26858
rect 16580 26794 16632 26800
rect 16592 26314 16620 26794
rect 16672 26784 16724 26790
rect 16672 26726 16724 26732
rect 16684 26382 16712 26726
rect 16672 26376 16724 26382
rect 16672 26318 16724 26324
rect 16580 26308 16632 26314
rect 16580 26250 16632 26256
rect 16672 26240 16724 26246
rect 16672 26182 16724 26188
rect 16684 26042 16712 26182
rect 16672 26036 16724 26042
rect 16672 25978 16724 25984
rect 16396 25356 16448 25362
rect 16396 25298 16448 25304
rect 16304 25220 16356 25226
rect 16304 25162 16356 25168
rect 16672 25220 16724 25226
rect 16672 25162 16724 25168
rect 16212 24880 16264 24886
rect 16212 24822 16264 24828
rect 16212 24064 16264 24070
rect 16212 24006 16264 24012
rect 16224 23186 16252 24006
rect 16212 23180 16264 23186
rect 16212 23122 16264 23128
rect 16120 22092 16172 22098
rect 16316 22094 16344 25162
rect 16488 25152 16540 25158
rect 16488 25094 16540 25100
rect 16500 24954 16528 25094
rect 16488 24948 16540 24954
rect 16488 24890 16540 24896
rect 16120 22034 16172 22040
rect 16224 22066 16344 22094
rect 16120 21956 16172 21962
rect 16120 21898 16172 21904
rect 16132 21350 16160 21898
rect 16120 21344 16172 21350
rect 16120 21286 16172 21292
rect 16120 20528 16172 20534
rect 16120 20470 16172 20476
rect 16028 20460 16080 20466
rect 16028 20402 16080 20408
rect 16028 20324 16080 20330
rect 16028 20266 16080 20272
rect 16040 19922 16068 20266
rect 16028 19916 16080 19922
rect 16028 19858 16080 19864
rect 15936 18692 15988 18698
rect 15936 18634 15988 18640
rect 15948 18222 15976 18634
rect 16040 18290 16068 19858
rect 16028 18284 16080 18290
rect 16028 18226 16080 18232
rect 15936 18216 15988 18222
rect 15936 18158 15988 18164
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 15948 17610 15976 18158
rect 16028 18080 16080 18086
rect 16028 18022 16080 18028
rect 15844 17604 15896 17610
rect 15844 17546 15896 17552
rect 15936 17604 15988 17610
rect 15936 17546 15988 17552
rect 15856 17202 15884 17546
rect 15844 17196 15896 17202
rect 15844 17138 15896 17144
rect 15752 17060 15804 17066
rect 15752 17002 15804 17008
rect 15580 16510 15792 16538
rect 15384 16448 15436 16454
rect 15384 16390 15436 16396
rect 15568 16448 15620 16454
rect 15568 16390 15620 16396
rect 15292 16176 15344 16182
rect 15292 16118 15344 16124
rect 15212 15150 15332 15178
rect 15108 15020 15160 15026
rect 15108 14962 15160 14968
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 15120 14346 15148 14962
rect 15200 14612 15252 14618
rect 15200 14554 15252 14560
rect 15108 14340 15160 14346
rect 15108 14282 15160 14288
rect 15016 13728 15068 13734
rect 15016 13670 15068 13676
rect 15028 13308 15056 13670
rect 15120 13462 15148 14282
rect 15108 13456 15160 13462
rect 15108 13398 15160 13404
rect 15108 13320 15160 13326
rect 15028 13280 15108 13308
rect 14924 13252 14976 13258
rect 14924 13194 14976 13200
rect 14924 12980 14976 12986
rect 14924 12922 14976 12928
rect 14740 12844 14792 12850
rect 14740 12786 14792 12792
rect 14752 12238 14780 12786
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 14464 9988 14516 9994
rect 14464 9930 14516 9936
rect 14372 9648 14424 9654
rect 14372 9590 14424 9596
rect 14384 9110 14412 9590
rect 14372 9104 14424 9110
rect 14372 9046 14424 9052
rect 14372 8356 14424 8362
rect 14372 8298 14424 8304
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14292 6934 14320 7346
rect 14280 6928 14332 6934
rect 14280 6870 14332 6876
rect 14384 6798 14412 8298
rect 14476 6866 14504 9930
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 14660 8362 14688 9522
rect 14648 8356 14700 8362
rect 14648 8298 14700 8304
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14752 7410 14780 7822
rect 14740 7404 14792 7410
rect 14740 7346 14792 7352
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14752 6866 14780 7142
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14740 6860 14792 6866
rect 14740 6802 14792 6808
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 14004 4276 14056 4282
rect 14004 4218 14056 4224
rect 13820 3732 13872 3738
rect 13820 3674 13872 3680
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 13832 1426 13860 3130
rect 14200 2990 14228 6394
rect 14384 6322 14412 6734
rect 14936 6458 14964 12922
rect 15028 10810 15056 13280
rect 15108 13262 15160 13268
rect 15108 13184 15160 13190
rect 15108 13126 15160 13132
rect 15120 12306 15148 13126
rect 15108 12300 15160 12306
rect 15108 12242 15160 12248
rect 15212 11354 15240 14554
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 15200 11008 15252 11014
rect 15200 10950 15252 10956
rect 15016 10804 15068 10810
rect 15016 10746 15068 10752
rect 15212 10674 15240 10950
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 15108 9444 15160 9450
rect 15108 9386 15160 9392
rect 15120 7886 15148 9386
rect 15108 7880 15160 7886
rect 15108 7822 15160 7828
rect 15016 7812 15068 7818
rect 15016 7754 15068 7760
rect 15028 7410 15056 7754
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 15120 7274 15148 7822
rect 15108 7268 15160 7274
rect 15108 7210 15160 7216
rect 15016 6860 15068 6866
rect 15016 6802 15068 6808
rect 15028 6458 15056 6802
rect 14924 6452 14976 6458
rect 14924 6394 14976 6400
rect 15016 6452 15068 6458
rect 15016 6394 15068 6400
rect 14372 6316 14424 6322
rect 14372 6258 14424 6264
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 14280 5228 14332 5234
rect 14280 5170 14332 5176
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 14292 4282 14320 5170
rect 14384 4690 14412 5170
rect 14752 4826 14780 6258
rect 15016 6112 15068 6118
rect 15016 6054 15068 6060
rect 15028 5778 15056 6054
rect 15016 5772 15068 5778
rect 15016 5714 15068 5720
rect 14924 5704 14976 5710
rect 14924 5646 14976 5652
rect 14832 5228 14884 5234
rect 14832 5170 14884 5176
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14372 4684 14424 4690
rect 14372 4626 14424 4632
rect 14280 4276 14332 4282
rect 14280 4218 14332 4224
rect 14292 4146 14320 4218
rect 14384 4146 14412 4626
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14292 3534 14320 4082
rect 14384 3534 14412 4082
rect 14844 3534 14872 5170
rect 14936 5166 14964 5646
rect 15108 5568 15160 5574
rect 15304 5534 15332 15150
rect 15396 13938 15424 16390
rect 15476 16108 15528 16114
rect 15580 16096 15608 16390
rect 15528 16068 15608 16096
rect 15476 16050 15528 16056
rect 15580 15994 15608 16068
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 15488 15966 15608 15994
rect 15488 14482 15516 15966
rect 15672 15162 15700 16050
rect 15660 15156 15712 15162
rect 15580 15116 15660 15144
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 15384 13932 15436 13938
rect 15384 13874 15436 13880
rect 15580 13870 15608 15116
rect 15660 15098 15712 15104
rect 15764 14822 15792 16510
rect 15856 16454 15884 17138
rect 15844 16448 15896 16454
rect 15844 16390 15896 16396
rect 15844 16176 15896 16182
rect 15844 16118 15896 16124
rect 15856 15094 15884 16118
rect 15948 15502 15976 17546
rect 15936 15496 15988 15502
rect 15936 15438 15988 15444
rect 16040 15194 16068 18022
rect 15948 15166 16068 15194
rect 15844 15088 15896 15094
rect 15844 15030 15896 15036
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15568 13864 15620 13870
rect 15568 13806 15620 13812
rect 15672 13814 15700 14758
rect 15948 14482 15976 15166
rect 16132 15026 16160 20470
rect 16224 16998 16252 22066
rect 16304 21684 16356 21690
rect 16304 21626 16356 21632
rect 16316 20874 16344 21626
rect 16396 21344 16448 21350
rect 16396 21286 16448 21292
rect 16304 20868 16356 20874
rect 16304 20810 16356 20816
rect 16304 20324 16356 20330
rect 16304 20266 16356 20272
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 16224 15366 16252 16934
rect 16316 16590 16344 20266
rect 16304 16584 16356 16590
rect 16304 16526 16356 16532
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 16212 15360 16264 15366
rect 16212 15302 16264 15308
rect 16224 15162 16252 15302
rect 16212 15156 16264 15162
rect 16212 15098 16264 15104
rect 16120 15020 16172 15026
rect 16120 14962 16172 14968
rect 16028 14816 16080 14822
rect 16028 14758 16080 14764
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 15936 14476 15988 14482
rect 15936 14418 15988 14424
rect 15752 14272 15804 14278
rect 15752 14214 15804 14220
rect 15764 14056 15792 14214
rect 15764 14028 15884 14056
rect 15856 13938 15884 14028
rect 15844 13932 15896 13938
rect 15844 13874 15896 13880
rect 15936 13932 15988 13938
rect 15936 13874 15988 13880
rect 15672 13786 15792 13814
rect 15384 13728 15436 13734
rect 15384 13670 15436 13676
rect 15568 13728 15620 13734
rect 15568 13670 15620 13676
rect 15396 12442 15424 13670
rect 15580 12918 15608 13670
rect 15764 13394 15792 13786
rect 15948 13462 15976 13874
rect 15936 13456 15988 13462
rect 15936 13398 15988 13404
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 16040 13308 16068 14758
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 16132 13802 16160 14350
rect 16224 14074 16252 14758
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 16120 13796 16172 13802
rect 16120 13738 16172 13744
rect 15948 13280 16068 13308
rect 15844 13252 15896 13258
rect 15844 13194 15896 13200
rect 15568 12912 15620 12918
rect 15568 12854 15620 12860
rect 15384 12436 15436 12442
rect 15384 12378 15436 12384
rect 15856 11898 15884 13194
rect 15948 12186 15976 13280
rect 16028 12776 16080 12782
rect 16028 12718 16080 12724
rect 16040 12306 16068 12718
rect 16132 12714 16160 13738
rect 16224 13394 16252 13806
rect 16212 13388 16264 13394
rect 16212 13330 16264 13336
rect 16316 13326 16344 15846
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 16120 12708 16172 12714
rect 16120 12650 16172 12656
rect 16028 12300 16080 12306
rect 16028 12242 16080 12248
rect 15948 12158 16068 12186
rect 15936 12096 15988 12102
rect 15936 12038 15988 12044
rect 15844 11892 15896 11898
rect 15844 11834 15896 11840
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 15396 8430 15424 11290
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 15764 8838 15792 9318
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 15660 8492 15712 8498
rect 15660 8434 15712 8440
rect 15384 8424 15436 8430
rect 15436 8384 15608 8412
rect 15384 8366 15436 8372
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 15384 7336 15436 7342
rect 15384 7278 15436 7284
rect 15396 6866 15424 7278
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15396 5574 15424 6394
rect 15488 6254 15516 7346
rect 15476 6248 15528 6254
rect 15476 6190 15528 6196
rect 15108 5510 15160 5516
rect 15120 5166 15148 5510
rect 15212 5506 15332 5534
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 14924 5160 14976 5166
rect 14924 5102 14976 5108
rect 15108 5160 15160 5166
rect 15108 5102 15160 5108
rect 15016 5092 15068 5098
rect 15016 5034 15068 5040
rect 15028 4826 15056 5034
rect 15016 4820 15068 4826
rect 15016 4762 15068 4768
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 15016 4616 15068 4622
rect 15016 4558 15068 4564
rect 15028 4214 15056 4558
rect 15120 4264 15148 4626
rect 15212 4554 15240 5506
rect 15384 5160 15436 5166
rect 15304 5120 15384 5148
rect 15200 4548 15252 4554
rect 15200 4490 15252 4496
rect 15200 4276 15252 4282
rect 15120 4236 15200 4264
rect 15200 4218 15252 4224
rect 15016 4208 15068 4214
rect 15016 4150 15068 4156
rect 15304 3602 15332 5120
rect 15384 5102 15436 5108
rect 15580 5030 15608 8384
rect 15672 7546 15700 8434
rect 15660 7540 15712 7546
rect 15660 7482 15712 7488
rect 15752 6860 15804 6866
rect 15672 6820 15752 6848
rect 15672 5710 15700 6820
rect 15752 6802 15804 6808
rect 15856 6662 15884 11834
rect 15948 10742 15976 12038
rect 16040 11540 16068 12158
rect 16132 11694 16160 12650
rect 16316 12374 16344 13262
rect 16304 12368 16356 12374
rect 16304 12310 16356 12316
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 16040 11512 16160 11540
rect 15936 10736 15988 10742
rect 15936 10678 15988 10684
rect 16132 10674 16160 11512
rect 16028 10668 16080 10674
rect 16028 10610 16080 10616
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 16040 10266 16068 10610
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 16132 9586 16160 9862
rect 16120 9580 16172 9586
rect 16120 9522 16172 9528
rect 16212 9580 16264 9586
rect 16212 9522 16264 9528
rect 15936 9036 15988 9042
rect 15936 8978 15988 8984
rect 15948 8838 15976 8978
rect 15936 8832 15988 8838
rect 15936 8774 15988 8780
rect 15948 7886 15976 8774
rect 16028 8016 16080 8022
rect 16028 7958 16080 7964
rect 16132 7970 16160 9522
rect 16224 8090 16252 9522
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16316 8974 16344 9318
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16212 8084 16264 8090
rect 16212 8026 16264 8032
rect 15936 7880 15988 7886
rect 15936 7822 15988 7828
rect 15948 7206 15976 7822
rect 16040 7410 16068 7958
rect 16132 7942 16252 7970
rect 16028 7404 16080 7410
rect 16028 7346 16080 7352
rect 15936 7200 15988 7206
rect 15936 7142 15988 7148
rect 15844 6656 15896 6662
rect 15844 6598 15896 6604
rect 16028 6656 16080 6662
rect 16028 6598 16080 6604
rect 16040 6440 16068 6598
rect 15948 6412 16068 6440
rect 15948 6118 15976 6412
rect 16120 6384 16172 6390
rect 16120 6326 16172 6332
rect 16028 6248 16080 6254
rect 16028 6190 16080 6196
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15936 5772 15988 5778
rect 15936 5714 15988 5720
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 15672 5166 15700 5646
rect 15764 5574 15792 5646
rect 15752 5568 15804 5574
rect 15752 5510 15804 5516
rect 15660 5160 15712 5166
rect 15660 5102 15712 5108
rect 15764 5098 15792 5510
rect 15752 5092 15804 5098
rect 15752 5034 15804 5040
rect 15568 5024 15620 5030
rect 15568 4966 15620 4972
rect 15580 4706 15608 4966
rect 15488 4678 15608 4706
rect 15488 3602 15516 4678
rect 15568 4548 15620 4554
rect 15568 4490 15620 4496
rect 15580 3602 15608 4490
rect 15764 4486 15792 5034
rect 15948 4842 15976 5714
rect 16040 5574 16068 6190
rect 16028 5568 16080 5574
rect 16028 5510 16080 5516
rect 15948 4814 16068 4842
rect 16040 4758 16068 4814
rect 15844 4752 15896 4758
rect 15844 4694 15896 4700
rect 16028 4752 16080 4758
rect 16028 4694 16080 4700
rect 15752 4480 15804 4486
rect 15752 4422 15804 4428
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15568 3596 15620 3602
rect 15568 3538 15620 3544
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 14292 3058 14320 3470
rect 14384 3126 14412 3470
rect 14844 3194 14872 3470
rect 15580 3194 15608 3538
rect 14832 3188 14884 3194
rect 14832 3130 14884 3136
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 14372 3120 14424 3126
rect 14372 3062 14424 3068
rect 15660 3120 15712 3126
rect 15660 3062 15712 3068
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 14292 2650 14320 2994
rect 14924 2848 14976 2854
rect 14924 2790 14976 2796
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 14556 2508 14608 2514
rect 14556 2450 14608 2456
rect 14096 2304 14148 2310
rect 14096 2246 14148 2252
rect 13820 1420 13872 1426
rect 13820 1362 13872 1368
rect 14108 1222 14136 2246
rect 14568 1970 14596 2450
rect 14556 1964 14608 1970
rect 14556 1906 14608 1912
rect 14832 1964 14884 1970
rect 14832 1906 14884 1912
rect 14844 1562 14872 1906
rect 14832 1556 14884 1562
rect 14832 1498 14884 1504
rect 14936 1358 14964 2790
rect 15672 2774 15700 3062
rect 15764 3058 15792 4422
rect 15856 4146 15884 4694
rect 15936 4548 15988 4554
rect 15936 4490 15988 4496
rect 15948 4282 15976 4490
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 15844 4140 15896 4146
rect 15844 4082 15896 4088
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 15752 3052 15804 3058
rect 15752 2994 15804 3000
rect 15844 2848 15896 2854
rect 15844 2790 15896 2796
rect 15672 2746 15792 2774
rect 15660 2372 15712 2378
rect 15660 2314 15712 2320
rect 15672 1562 15700 2314
rect 15764 1766 15792 2746
rect 15752 1760 15804 1766
rect 15752 1702 15804 1708
rect 15660 1556 15712 1562
rect 15660 1498 15712 1504
rect 15856 1358 15884 2790
rect 15936 2304 15988 2310
rect 15936 2246 15988 2252
rect 15948 1426 15976 2246
rect 15936 1420 15988 1426
rect 15936 1362 15988 1368
rect 16040 1358 16068 3470
rect 16132 3126 16160 6326
rect 16120 3120 16172 3126
rect 16120 3062 16172 3068
rect 16224 2650 16252 7942
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16316 7206 16344 7890
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 16316 5642 16344 6258
rect 16304 5636 16356 5642
rect 16304 5578 16356 5584
rect 16316 4758 16344 5578
rect 16408 5370 16436 21286
rect 16500 19514 16528 24890
rect 16684 23118 16712 25162
rect 16776 23866 16804 28172
rect 16948 28076 17000 28082
rect 16948 28018 17000 28024
rect 16960 26994 16988 28018
rect 17052 27130 17080 28966
rect 17144 28218 17172 28970
rect 17132 28212 17184 28218
rect 17132 28154 17184 28160
rect 17040 27124 17092 27130
rect 17040 27066 17092 27072
rect 16948 26988 17000 26994
rect 16948 26930 17000 26936
rect 16960 26586 16988 26930
rect 16948 26580 17000 26586
rect 16948 26522 17000 26528
rect 16948 25968 17000 25974
rect 16948 25910 17000 25916
rect 16856 25832 16908 25838
rect 16856 25774 16908 25780
rect 16868 24274 16896 25774
rect 16960 24818 16988 25910
rect 16948 24812 17000 24818
rect 16948 24754 17000 24760
rect 16856 24268 16908 24274
rect 16856 24210 16908 24216
rect 16764 23860 16816 23866
rect 16764 23802 16816 23808
rect 16960 23526 16988 24754
rect 16948 23520 17000 23526
rect 16948 23462 17000 23468
rect 17052 23202 17080 27066
rect 17132 26784 17184 26790
rect 17132 26726 17184 26732
rect 17144 26586 17172 26726
rect 17132 26580 17184 26586
rect 17132 26522 17184 26528
rect 17132 26376 17184 26382
rect 17132 26318 17184 26324
rect 16868 23174 17080 23202
rect 16672 23112 16724 23118
rect 16672 23054 16724 23060
rect 16672 22976 16724 22982
rect 16672 22918 16724 22924
rect 16580 22772 16632 22778
rect 16580 22714 16632 22720
rect 16488 19508 16540 19514
rect 16488 19450 16540 19456
rect 16488 19372 16540 19378
rect 16488 19314 16540 19320
rect 16500 15706 16528 19314
rect 16592 16028 16620 22714
rect 16684 21622 16712 22918
rect 16764 22636 16816 22642
rect 16764 22578 16816 22584
rect 16776 21622 16804 22578
rect 16672 21616 16724 21622
rect 16672 21558 16724 21564
rect 16764 21616 16816 21622
rect 16764 21558 16816 21564
rect 16868 20618 16896 23174
rect 17040 23112 17092 23118
rect 17040 23054 17092 23060
rect 16948 22636 17000 22642
rect 16948 22578 17000 22584
rect 16960 20806 16988 22578
rect 17052 22574 17080 23054
rect 17144 22778 17172 26318
rect 17132 22772 17184 22778
rect 17132 22714 17184 22720
rect 17040 22568 17092 22574
rect 17040 22510 17092 22516
rect 17052 20924 17080 22510
rect 17132 22432 17184 22438
rect 17132 22374 17184 22380
rect 17144 22030 17172 22374
rect 17132 22024 17184 22030
rect 17132 21966 17184 21972
rect 17132 20936 17184 20942
rect 17052 20896 17132 20924
rect 17132 20878 17184 20884
rect 16948 20800 17000 20806
rect 16948 20742 17000 20748
rect 17040 20800 17092 20806
rect 17040 20742 17092 20748
rect 16684 20590 16896 20618
rect 16684 20534 16712 20590
rect 16672 20528 16724 20534
rect 16672 20470 16724 20476
rect 16764 20528 16816 20534
rect 16764 20470 16816 20476
rect 16672 20392 16724 20398
rect 16672 20334 16724 20340
rect 16684 19378 16712 20334
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16776 18850 16804 20470
rect 16948 20460 17000 20466
rect 16948 20402 17000 20408
rect 16856 20256 16908 20262
rect 16856 20198 16908 20204
rect 16868 19922 16896 20198
rect 16856 19916 16908 19922
rect 16856 19858 16908 19864
rect 16960 19514 16988 20402
rect 16948 19508 17000 19514
rect 16948 19450 17000 19456
rect 17052 19334 17080 20742
rect 17144 19378 17172 20878
rect 17236 20806 17264 31726
rect 17408 31680 17460 31686
rect 17408 31622 17460 31628
rect 17316 31340 17368 31346
rect 17316 31282 17368 31288
rect 17328 30938 17356 31282
rect 17316 30932 17368 30938
rect 17316 30874 17368 30880
rect 17420 30598 17448 31622
rect 17590 31578 17646 32614
rect 17880 32570 17908 33458
rect 18236 33312 18288 33318
rect 18236 33254 18288 33260
rect 18248 32842 18276 33254
rect 18236 32836 18288 32842
rect 18236 32778 18288 32784
rect 17868 32564 17920 32570
rect 17868 32506 17920 32512
rect 17684 32428 17736 32434
rect 17684 32370 17736 32376
rect 18144 32428 18196 32434
rect 18144 32370 18196 32376
rect 17590 31526 17592 31578
rect 17644 31526 17646 31578
rect 17408 30592 17460 30598
rect 17408 30534 17460 30540
rect 17590 30490 17646 31526
rect 17696 31464 17724 32370
rect 17776 32292 17828 32298
rect 17776 32234 17828 32240
rect 17788 31754 17816 32234
rect 17960 32224 18012 32230
rect 17960 32166 18012 32172
rect 17868 31952 17920 31958
rect 17868 31894 17920 31900
rect 17776 31748 17828 31754
rect 17776 31690 17828 31696
rect 17696 31436 17816 31464
rect 17788 30938 17816 31436
rect 17776 30932 17828 30938
rect 17776 30874 17828 30880
rect 17590 30438 17592 30490
rect 17644 30438 17646 30490
rect 17500 30252 17552 30258
rect 17500 30194 17552 30200
rect 17316 29504 17368 29510
rect 17316 29446 17368 29452
rect 17328 29170 17356 29446
rect 17316 29164 17368 29170
rect 17316 29106 17368 29112
rect 17408 29164 17460 29170
rect 17408 29106 17460 29112
rect 17316 28552 17368 28558
rect 17316 28494 17368 28500
rect 17328 27470 17356 28494
rect 17316 27464 17368 27470
rect 17316 27406 17368 27412
rect 17328 25838 17356 27406
rect 17420 26382 17448 29106
rect 17512 26382 17540 30194
rect 17590 29402 17646 30438
rect 17684 29504 17736 29510
rect 17684 29446 17736 29452
rect 17590 29350 17592 29402
rect 17644 29350 17646 29402
rect 17590 28314 17646 29350
rect 17696 29170 17724 29446
rect 17776 29300 17828 29306
rect 17776 29242 17828 29248
rect 17684 29164 17736 29170
rect 17684 29106 17736 29112
rect 17590 28262 17592 28314
rect 17644 28262 17646 28314
rect 17590 27226 17646 28262
rect 17684 27396 17736 27402
rect 17684 27338 17736 27344
rect 17590 27174 17592 27226
rect 17644 27174 17646 27226
rect 17408 26376 17460 26382
rect 17408 26318 17460 26324
rect 17500 26376 17552 26382
rect 17500 26318 17552 26324
rect 17316 25832 17368 25838
rect 17512 25786 17540 26318
rect 17316 25774 17368 25780
rect 17420 25758 17540 25786
rect 17590 26138 17646 27174
rect 17696 27130 17724 27338
rect 17684 27124 17736 27130
rect 17684 27066 17736 27072
rect 17590 26086 17592 26138
rect 17644 26086 17646 26138
rect 17420 25702 17448 25758
rect 17408 25696 17460 25702
rect 17408 25638 17460 25644
rect 17590 25050 17646 26086
rect 17590 24998 17592 25050
rect 17644 24998 17646 25050
rect 17316 24744 17368 24750
rect 17316 24686 17368 24692
rect 17328 23254 17356 24686
rect 17500 24132 17552 24138
rect 17500 24074 17552 24080
rect 17408 23520 17460 23526
rect 17408 23462 17460 23468
rect 17316 23248 17368 23254
rect 17316 23190 17368 23196
rect 17224 20800 17276 20806
rect 17224 20742 17276 20748
rect 17224 20596 17276 20602
rect 17224 20538 17276 20544
rect 17236 19922 17264 20538
rect 17224 19916 17276 19922
rect 17224 19858 17276 19864
rect 16684 18834 16804 18850
rect 16672 18828 16804 18834
rect 16724 18822 16804 18828
rect 16868 19306 17080 19334
rect 17132 19372 17184 19378
rect 17132 19314 17184 19320
rect 16672 18770 16724 18776
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 16776 18290 16804 18702
rect 16764 18284 16816 18290
rect 16764 18226 16816 18232
rect 16672 17672 16724 17678
rect 16672 17614 16724 17620
rect 16684 17202 16712 17614
rect 16868 17490 16896 19306
rect 17236 19258 17264 19858
rect 17144 19230 17264 19258
rect 17040 19168 17092 19174
rect 17040 19110 17092 19116
rect 17052 18698 17080 19110
rect 17040 18692 17092 18698
rect 17040 18634 17092 18640
rect 16948 17604 17000 17610
rect 16776 17462 16896 17490
rect 16940 17552 16948 17592
rect 16940 17546 17000 17552
rect 16776 17252 16804 17462
rect 16940 17354 16968 17546
rect 17144 17542 17172 19230
rect 17224 19168 17276 19174
rect 17224 19110 17276 19116
rect 17236 18766 17264 19110
rect 17224 18760 17276 18766
rect 17224 18702 17276 18708
rect 17224 18624 17276 18630
rect 17224 18566 17276 18572
rect 17236 17814 17264 18566
rect 17224 17808 17276 17814
rect 17224 17750 17276 17756
rect 17132 17536 17184 17542
rect 17132 17478 17184 17484
rect 16940 17326 17080 17354
rect 16776 17224 16896 17252
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16684 16640 16712 17138
rect 16764 16652 16816 16658
rect 16684 16612 16764 16640
rect 16764 16594 16816 16600
rect 16592 16000 16712 16028
rect 16684 15722 16712 16000
rect 16488 15700 16540 15706
rect 16488 15642 16540 15648
rect 16592 15694 16712 15722
rect 16592 15552 16620 15694
rect 16583 15524 16620 15552
rect 16488 15496 16540 15502
rect 16583 15484 16611 15524
rect 16583 15456 16620 15484
rect 16488 15438 16540 15444
rect 16500 13938 16528 15438
rect 16488 13932 16540 13938
rect 16488 13874 16540 13880
rect 16488 13320 16540 13326
rect 16488 13262 16540 13268
rect 16500 12782 16528 13262
rect 16592 12918 16620 15456
rect 16776 15026 16804 16594
rect 16868 15450 16896 17224
rect 17052 17202 17080 17326
rect 17132 17264 17184 17270
rect 17132 17206 17184 17212
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 16948 17060 17000 17066
rect 17144 17048 17172 17206
rect 16948 17002 17000 17008
rect 17052 17020 17172 17048
rect 16960 16130 16988 17002
rect 17052 16590 17080 17020
rect 17328 16810 17356 23190
rect 17420 22522 17448 23462
rect 17512 22778 17540 24074
rect 17590 23962 17646 24998
rect 17590 23910 17592 23962
rect 17644 23910 17646 23962
rect 17590 22874 17646 23910
rect 17684 23316 17736 23322
rect 17684 23258 17736 23264
rect 17590 22822 17592 22874
rect 17644 22822 17646 22874
rect 17500 22772 17552 22778
rect 17500 22714 17552 22720
rect 17420 22494 17540 22522
rect 17408 22432 17460 22438
rect 17408 22374 17460 22380
rect 17420 22234 17448 22374
rect 17408 22228 17460 22234
rect 17408 22170 17460 22176
rect 17408 22092 17460 22098
rect 17408 22034 17460 22040
rect 17420 18426 17448 22034
rect 17512 19922 17540 22494
rect 17590 21786 17646 22822
rect 17696 21894 17724 23258
rect 17788 22710 17816 29242
rect 17880 26994 17908 31894
rect 17972 31686 18000 32166
rect 18156 31890 18184 32370
rect 18144 31884 18196 31890
rect 18144 31826 18196 31832
rect 17960 31680 18012 31686
rect 17960 31622 18012 31628
rect 18248 31346 18276 32778
rect 18328 31816 18380 31822
rect 18328 31758 18380 31764
rect 17960 31340 18012 31346
rect 17960 31282 18012 31288
rect 18236 31340 18288 31346
rect 18236 31282 18288 31288
rect 17972 30258 18000 31282
rect 18052 30728 18104 30734
rect 18052 30670 18104 30676
rect 17960 30252 18012 30258
rect 17960 30194 18012 30200
rect 17972 29646 18000 30194
rect 17960 29640 18012 29646
rect 17960 29582 18012 29588
rect 17960 29096 18012 29102
rect 17960 29038 18012 29044
rect 17972 28218 18000 29038
rect 18064 28558 18092 30670
rect 18144 30592 18196 30598
rect 18144 30534 18196 30540
rect 18156 30258 18184 30534
rect 18236 30388 18288 30394
rect 18236 30330 18288 30336
rect 18144 30252 18196 30258
rect 18144 30194 18196 30200
rect 18156 29102 18184 30194
rect 18248 29714 18276 30330
rect 18236 29708 18288 29714
rect 18236 29650 18288 29656
rect 18340 29646 18368 31758
rect 18328 29640 18380 29646
rect 18328 29582 18380 29588
rect 18144 29096 18196 29102
rect 18144 29038 18196 29044
rect 18340 28762 18368 29582
rect 18328 28756 18380 28762
rect 18328 28698 18380 28704
rect 18052 28552 18104 28558
rect 18052 28494 18104 28500
rect 17960 28212 18012 28218
rect 17960 28154 18012 28160
rect 18340 28150 18368 28698
rect 18328 28144 18380 28150
rect 18328 28086 18380 28092
rect 18236 28076 18288 28082
rect 18236 28018 18288 28024
rect 17868 26988 17920 26994
rect 17868 26930 17920 26936
rect 18248 26518 18276 28018
rect 18432 27334 18460 33594
rect 18800 33522 18828 33798
rect 18788 33516 18840 33522
rect 18788 33458 18840 33464
rect 18788 32972 18840 32978
rect 18788 32914 18840 32920
rect 18512 31680 18564 31686
rect 18512 31622 18564 31628
rect 18524 30258 18552 31622
rect 18512 30252 18564 30258
rect 18512 30194 18564 30200
rect 18604 30184 18656 30190
rect 18604 30126 18656 30132
rect 18616 29782 18644 30126
rect 18696 30048 18748 30054
rect 18696 29990 18748 29996
rect 18604 29776 18656 29782
rect 18604 29718 18656 29724
rect 18708 29578 18736 29990
rect 18696 29572 18748 29578
rect 18696 29514 18748 29520
rect 18708 29102 18736 29514
rect 18696 29096 18748 29102
rect 18696 29038 18748 29044
rect 18708 28694 18736 29038
rect 18800 29034 18828 32914
rect 18788 29028 18840 29034
rect 18788 28970 18840 28976
rect 18696 28688 18748 28694
rect 18696 28630 18748 28636
rect 18512 28484 18564 28490
rect 18512 28426 18564 28432
rect 18420 27328 18472 27334
rect 18420 27270 18472 27276
rect 18420 26784 18472 26790
rect 18420 26726 18472 26732
rect 18236 26512 18288 26518
rect 18236 26454 18288 26460
rect 17960 26376 18012 26382
rect 17960 26318 18012 26324
rect 17868 24676 17920 24682
rect 17868 24618 17920 24624
rect 17880 23798 17908 24618
rect 17972 24070 18000 26318
rect 18236 26308 18288 26314
rect 18236 26250 18288 26256
rect 18052 25900 18104 25906
rect 18052 25842 18104 25848
rect 18064 25498 18092 25842
rect 18052 25492 18104 25498
rect 18052 25434 18104 25440
rect 18052 24948 18104 24954
rect 18052 24890 18104 24896
rect 17960 24064 18012 24070
rect 17960 24006 18012 24012
rect 17868 23792 17920 23798
rect 17868 23734 17920 23740
rect 17868 22976 17920 22982
rect 17868 22918 17920 22924
rect 17776 22704 17828 22710
rect 17776 22646 17828 22652
rect 17684 21888 17736 21894
rect 17684 21830 17736 21836
rect 17590 21734 17592 21786
rect 17644 21734 17646 21786
rect 17590 20698 17646 21734
rect 17788 21706 17816 22646
rect 17880 22642 17908 22918
rect 17868 22636 17920 22642
rect 17868 22578 17920 22584
rect 17788 21678 17908 21706
rect 17776 21412 17828 21418
rect 17776 21354 17828 21360
rect 17788 20942 17816 21354
rect 17684 20936 17736 20942
rect 17684 20878 17736 20884
rect 17776 20936 17828 20942
rect 17776 20878 17828 20884
rect 17590 20646 17592 20698
rect 17644 20646 17646 20698
rect 17500 19916 17552 19922
rect 17500 19858 17552 19864
rect 17590 19610 17646 20646
rect 17687 20618 17715 20878
rect 17880 20806 17908 21678
rect 17776 20800 17828 20806
rect 17776 20742 17828 20748
rect 17868 20800 17920 20806
rect 17868 20742 17920 20748
rect 17687 20590 17724 20618
rect 17590 19558 17592 19610
rect 17644 19558 17646 19610
rect 17590 18522 17646 19558
rect 17696 18698 17724 20590
rect 17788 19854 17816 20742
rect 17972 20618 18000 24006
rect 18064 22438 18092 24890
rect 18248 23186 18276 26250
rect 18432 25294 18460 26726
rect 18524 26042 18552 28426
rect 18696 28144 18748 28150
rect 18696 28086 18748 28092
rect 18604 27464 18656 27470
rect 18604 27406 18656 27412
rect 18616 26994 18644 27406
rect 18604 26988 18656 26994
rect 18604 26930 18656 26936
rect 18616 26234 18644 26930
rect 18708 26382 18736 28086
rect 18788 27396 18840 27402
rect 18788 27338 18840 27344
rect 18696 26376 18748 26382
rect 18696 26318 18748 26324
rect 18616 26206 18736 26234
rect 18512 26036 18564 26042
rect 18512 25978 18564 25984
rect 18708 25702 18736 26206
rect 18696 25696 18748 25702
rect 18696 25638 18748 25644
rect 18420 25288 18472 25294
rect 18420 25230 18472 25236
rect 18328 25220 18380 25226
rect 18328 25162 18380 25168
rect 18340 24818 18368 25162
rect 18432 24954 18460 25230
rect 18708 25226 18736 25638
rect 18696 25220 18748 25226
rect 18696 25162 18748 25168
rect 18420 24948 18472 24954
rect 18420 24890 18472 24896
rect 18328 24812 18380 24818
rect 18328 24754 18380 24760
rect 18340 24070 18368 24754
rect 18512 24608 18564 24614
rect 18512 24550 18564 24556
rect 18328 24064 18380 24070
rect 18328 24006 18380 24012
rect 18236 23180 18288 23186
rect 18236 23122 18288 23128
rect 18340 23118 18368 24006
rect 18144 23112 18196 23118
rect 18144 23054 18196 23060
rect 18328 23112 18380 23118
rect 18328 23054 18380 23060
rect 18052 22432 18104 22438
rect 18052 22374 18104 22380
rect 18052 22024 18104 22030
rect 18052 21966 18104 21972
rect 18064 20942 18092 21966
rect 18052 20936 18104 20942
rect 18052 20878 18104 20884
rect 18156 20874 18184 23054
rect 18236 22976 18288 22982
rect 18236 22918 18288 22924
rect 18248 22642 18276 22918
rect 18236 22636 18288 22642
rect 18236 22578 18288 22584
rect 18236 22160 18288 22166
rect 18236 22102 18288 22108
rect 18144 20868 18196 20874
rect 18144 20810 18196 20816
rect 17880 20590 18000 20618
rect 17880 20516 17908 20590
rect 17880 20488 18000 20516
rect 17776 19848 17828 19854
rect 17776 19790 17828 19796
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 17880 19496 17908 19790
rect 17880 19468 17917 19496
rect 17889 19394 17917 19468
rect 17849 19366 17917 19394
rect 17849 18816 17877 19366
rect 17972 19334 18000 20488
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 18064 19922 18092 19994
rect 18052 19916 18104 19922
rect 18052 19858 18104 19864
rect 18156 19446 18184 20810
rect 18248 20534 18276 22102
rect 18340 21962 18368 23054
rect 18420 22636 18472 22642
rect 18420 22578 18472 22584
rect 18328 21956 18380 21962
rect 18328 21898 18380 21904
rect 18328 21344 18380 21350
rect 18328 21286 18380 21292
rect 18236 20528 18288 20534
rect 18236 20470 18288 20476
rect 18236 20052 18288 20058
rect 18236 19994 18288 20000
rect 18144 19440 18196 19446
rect 18144 19382 18196 19388
rect 17972 19306 18092 19334
rect 17960 19168 18012 19174
rect 17960 19110 18012 19116
rect 17849 18788 17908 18816
rect 17684 18692 17736 18698
rect 17684 18634 17736 18640
rect 17590 18470 17592 18522
rect 17644 18470 17646 18522
rect 17408 18420 17460 18426
rect 17408 18362 17460 18368
rect 17408 18284 17460 18290
rect 17408 18226 17460 18232
rect 17420 17270 17448 18226
rect 17500 17808 17552 17814
rect 17500 17750 17552 17756
rect 17408 17264 17460 17270
rect 17408 17206 17460 17212
rect 17408 17060 17460 17066
rect 17408 17002 17460 17008
rect 17144 16782 17356 16810
rect 17040 16584 17092 16590
rect 17040 16526 17092 16532
rect 16960 16102 17080 16130
rect 17052 16046 17080 16102
rect 17040 16040 17092 16046
rect 17040 15982 17092 15988
rect 16948 15972 17000 15978
rect 16948 15914 17000 15920
rect 16960 15552 16988 15914
rect 17040 15564 17092 15570
rect 16960 15524 17040 15552
rect 17040 15506 17092 15512
rect 16868 15422 17080 15450
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16764 15020 16816 15026
rect 16764 14962 16816 14968
rect 16672 14068 16724 14074
rect 16672 14010 16724 14016
rect 16580 12912 16632 12918
rect 16580 12854 16632 12860
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 16684 10996 16712 14010
rect 16868 13870 16896 15302
rect 16948 15156 17000 15162
rect 16948 15098 17000 15104
rect 16960 15026 16988 15098
rect 16948 15020 17000 15026
rect 16948 14962 17000 14968
rect 16960 14056 16988 14962
rect 17052 14414 17080 15422
rect 17040 14408 17092 14414
rect 17040 14350 17092 14356
rect 16960 14028 17080 14056
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 16764 13864 16816 13870
rect 16764 13806 16816 13812
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16776 13530 16804 13806
rect 16764 13524 16816 13530
rect 16764 13466 16816 13472
rect 16856 13524 16908 13530
rect 16856 13466 16908 13472
rect 16764 12844 16816 12850
rect 16764 12786 16816 12792
rect 16776 12102 16804 12786
rect 16868 12288 16896 13466
rect 16960 12646 16988 13874
rect 17052 13410 17080 14028
rect 17144 13530 17172 16782
rect 17316 16720 17368 16726
rect 17316 16662 17368 16668
rect 17328 14600 17356 16662
rect 17420 16658 17448 17002
rect 17408 16652 17460 16658
rect 17408 16594 17460 16600
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 17236 14572 17356 14600
rect 17132 13524 17184 13530
rect 17132 13466 17184 13472
rect 17052 13382 17172 13410
rect 16948 12640 17000 12646
rect 16948 12582 17000 12588
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 16868 12260 16988 12288
rect 16960 12170 16988 12260
rect 16856 12164 16908 12170
rect 16856 12106 16908 12112
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16764 12096 16816 12102
rect 16764 12038 16816 12044
rect 16868 11830 16896 12106
rect 16856 11824 16908 11830
rect 16856 11766 16908 11772
rect 17052 11762 17080 12582
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 16684 10968 16896 10996
rect 16672 10600 16724 10606
rect 16672 10542 16724 10548
rect 16684 10198 16712 10542
rect 16672 10192 16724 10198
rect 16672 10134 16724 10140
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16500 8566 16528 8774
rect 16488 8560 16540 8566
rect 16488 8502 16540 8508
rect 16592 7546 16620 8910
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16684 7886 16712 8366
rect 16868 8090 16896 10968
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 17052 8974 17080 9318
rect 17040 8968 17092 8974
rect 17040 8910 17092 8916
rect 17052 8566 17080 8910
rect 17040 8560 17092 8566
rect 17040 8502 17092 8508
rect 16856 8084 16908 8090
rect 16856 8026 16908 8032
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16948 7812 17000 7818
rect 16948 7754 17000 7760
rect 16856 7744 16908 7750
rect 16856 7686 16908 7692
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 16488 6792 16540 6798
rect 16488 6734 16540 6740
rect 16500 6390 16528 6734
rect 16580 6724 16632 6730
rect 16580 6666 16632 6672
rect 16488 6384 16540 6390
rect 16488 6326 16540 6332
rect 16592 6202 16620 6666
rect 16764 6316 16816 6322
rect 16764 6258 16816 6264
rect 16500 6174 16620 6202
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 16500 5234 16528 6174
rect 16580 6112 16632 6118
rect 16580 6054 16632 6060
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 16396 5160 16448 5166
rect 16396 5102 16448 5108
rect 16304 4752 16356 4758
rect 16304 4694 16356 4700
rect 16408 4690 16436 5102
rect 16396 4684 16448 4690
rect 16396 4626 16448 4632
rect 16488 4276 16540 4282
rect 16488 4218 16540 4224
rect 16500 3602 16528 4218
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 16592 3534 16620 6054
rect 16776 3942 16804 6258
rect 16868 6118 16896 7686
rect 16960 7410 16988 7754
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 17144 7002 17172 13382
rect 17236 11234 17264 14572
rect 17316 14476 17368 14482
rect 17316 14418 17368 14424
rect 17328 13682 17356 14418
rect 17420 13802 17448 14758
rect 17408 13796 17460 13802
rect 17408 13738 17460 13744
rect 17328 13654 17448 13682
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 17328 11354 17356 11494
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17236 11206 17356 11234
rect 17224 8084 17276 8090
rect 17224 8026 17276 8032
rect 17132 6996 17184 7002
rect 17132 6938 17184 6944
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 17132 6792 17184 6798
rect 17132 6734 17184 6740
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 16960 5846 16988 6734
rect 16948 5840 17000 5846
rect 16948 5782 17000 5788
rect 17040 5704 17092 5710
rect 17040 5646 17092 5652
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 16868 4622 16896 5170
rect 16948 5024 17000 5030
rect 16948 4966 17000 4972
rect 16856 4616 16908 4622
rect 16856 4558 16908 4564
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16868 3670 16896 4558
rect 16960 4146 16988 4966
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 16948 4004 17000 4010
rect 16948 3946 17000 3952
rect 16856 3664 16908 3670
rect 16856 3606 16908 3612
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 16488 3460 16540 3466
rect 16488 3402 16540 3408
rect 16500 3126 16528 3402
rect 16488 3120 16540 3126
rect 16488 3062 16540 3068
rect 16212 2644 16264 2650
rect 16212 2586 16264 2592
rect 16224 2446 16252 2586
rect 16212 2440 16264 2446
rect 16212 2382 16264 2388
rect 16672 2372 16724 2378
rect 16672 2314 16724 2320
rect 16580 1896 16632 1902
rect 16580 1838 16632 1844
rect 16592 1358 16620 1838
rect 16684 1562 16712 2314
rect 16776 1902 16804 3470
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 16868 2922 16896 2994
rect 16960 2990 16988 3946
rect 17052 3738 17080 5646
rect 17144 4554 17172 6734
rect 17236 6390 17264 8026
rect 17328 6798 17356 11206
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 17224 6384 17276 6390
rect 17224 6326 17276 6332
rect 17236 5658 17264 6326
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17328 5778 17356 6258
rect 17316 5772 17368 5778
rect 17316 5714 17368 5720
rect 17236 5642 17356 5658
rect 17236 5636 17368 5642
rect 17236 5630 17316 5636
rect 17316 5578 17368 5584
rect 17224 5568 17276 5574
rect 17224 5510 17276 5516
rect 17132 4548 17184 4554
rect 17132 4490 17184 4496
rect 17236 4214 17264 5510
rect 17316 5228 17368 5234
rect 17316 5170 17368 5176
rect 17328 4758 17356 5170
rect 17316 4752 17368 4758
rect 17316 4694 17368 4700
rect 17316 4616 17368 4622
rect 17316 4558 17368 4564
rect 17224 4208 17276 4214
rect 17224 4150 17276 4156
rect 17040 3732 17092 3738
rect 17040 3674 17092 3680
rect 17328 3584 17356 4558
rect 17144 3556 17356 3584
rect 17040 3460 17092 3466
rect 17040 3402 17092 3408
rect 16948 2984 17000 2990
rect 16948 2926 17000 2932
rect 16856 2916 16908 2922
rect 16856 2858 16908 2864
rect 16868 1970 16896 2858
rect 17052 2310 17080 3402
rect 17144 3058 17172 3556
rect 17236 3466 17264 3556
rect 17224 3460 17276 3466
rect 17224 3402 17276 3408
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 17040 2304 17092 2310
rect 17040 2246 17092 2252
rect 17144 1970 17172 2994
rect 17328 2310 17356 2994
rect 17316 2304 17368 2310
rect 17316 2246 17368 2252
rect 16856 1964 16908 1970
rect 16856 1906 16908 1912
rect 17132 1964 17184 1970
rect 17132 1906 17184 1912
rect 16764 1896 16816 1902
rect 16764 1838 16816 1844
rect 16856 1760 16908 1766
rect 16856 1702 16908 1708
rect 16672 1556 16724 1562
rect 16672 1498 16724 1504
rect 16868 1358 16896 1702
rect 14924 1352 14976 1358
rect 14924 1294 14976 1300
rect 15844 1352 15896 1358
rect 15844 1294 15896 1300
rect 16028 1352 16080 1358
rect 16028 1294 16080 1300
rect 16580 1352 16632 1358
rect 16580 1294 16632 1300
rect 16856 1352 16908 1358
rect 16856 1294 16908 1300
rect 16040 1222 16068 1294
rect 13728 1216 13780 1222
rect 13728 1158 13780 1164
rect 14096 1216 14148 1222
rect 14096 1158 14148 1164
rect 16028 1216 16080 1222
rect 16028 1158 16080 1164
rect 17420 1018 17448 13654
rect 17512 13258 17540 17750
rect 17590 17434 17646 18470
rect 17776 18420 17828 18426
rect 17776 18362 17828 18368
rect 17684 17536 17736 17542
rect 17684 17478 17736 17484
rect 17590 17382 17592 17434
rect 17644 17382 17646 17434
rect 17590 16346 17646 17382
rect 17696 17338 17724 17478
rect 17684 17332 17736 17338
rect 17684 17274 17736 17280
rect 17788 17184 17816 18362
rect 17880 18154 17908 18788
rect 17972 18630 18000 19110
rect 18064 18986 18092 19306
rect 18064 18958 18184 18986
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 18156 18578 18184 18958
rect 18248 18834 18276 19994
rect 18340 19990 18368 21286
rect 18432 21146 18460 22578
rect 18420 21140 18472 21146
rect 18420 21082 18472 21088
rect 18420 20936 18472 20942
rect 18420 20878 18472 20884
rect 18328 19984 18380 19990
rect 18328 19926 18380 19932
rect 18328 19508 18380 19514
rect 18328 19450 18380 19456
rect 18236 18828 18288 18834
rect 18236 18770 18288 18776
rect 18340 18766 18368 19450
rect 18432 19378 18460 20878
rect 18524 19802 18552 24550
rect 18604 23724 18656 23730
rect 18604 23666 18656 23672
rect 18616 23526 18644 23666
rect 18604 23520 18656 23526
rect 18604 23462 18656 23468
rect 18708 22624 18736 25162
rect 18800 22778 18828 27338
rect 18788 22772 18840 22778
rect 18788 22714 18840 22720
rect 18788 22636 18840 22642
rect 18708 22596 18788 22624
rect 18788 22578 18840 22584
rect 18892 22438 18920 35022
rect 19156 34944 19208 34950
rect 19156 34886 19208 34892
rect 18972 32428 19024 32434
rect 18972 32370 19024 32376
rect 18984 31482 19012 32370
rect 19064 31680 19116 31686
rect 19064 31622 19116 31628
rect 19076 31482 19104 31622
rect 18972 31476 19024 31482
rect 18972 31418 19024 31424
rect 19064 31476 19116 31482
rect 19064 31418 19116 31424
rect 19168 31346 19196 34886
rect 19340 34400 19392 34406
rect 19340 34342 19392 34348
rect 19352 33998 19380 34342
rect 19340 33992 19392 33998
rect 19340 33934 19392 33940
rect 19352 33590 19380 33934
rect 19340 33584 19392 33590
rect 19340 33526 19392 33532
rect 19616 32904 19668 32910
rect 19616 32846 19668 32852
rect 19340 32564 19392 32570
rect 19340 32506 19392 32512
rect 19248 31816 19300 31822
rect 19248 31758 19300 31764
rect 19156 31340 19208 31346
rect 19156 31282 19208 31288
rect 19168 30734 19196 31282
rect 19260 30802 19288 31758
rect 19352 31754 19380 32506
rect 19524 32496 19576 32502
rect 19524 32438 19576 32444
rect 19432 32224 19484 32230
rect 19432 32166 19484 32172
rect 19444 31804 19472 32166
rect 19536 31906 19564 32438
rect 19628 32434 19656 32846
rect 19708 32768 19760 32774
rect 19708 32710 19760 32716
rect 19616 32428 19668 32434
rect 19616 32370 19668 32376
rect 19720 32230 19748 32710
rect 19708 32224 19760 32230
rect 19708 32166 19760 32172
rect 19536 31878 19656 31906
rect 19524 31816 19576 31822
rect 19444 31776 19524 31804
rect 19524 31758 19576 31764
rect 19340 31748 19392 31754
rect 19340 31690 19392 31696
rect 19352 31634 19380 31690
rect 19352 31606 19472 31634
rect 19340 31476 19392 31482
rect 19340 31418 19392 31424
rect 19248 30796 19300 30802
rect 19248 30738 19300 30744
rect 19156 30728 19208 30734
rect 19156 30670 19208 30676
rect 19168 30394 19196 30670
rect 19248 30660 19300 30666
rect 19248 30602 19300 30608
rect 19156 30388 19208 30394
rect 19156 30330 19208 30336
rect 19260 30326 19288 30602
rect 19352 30326 19380 31418
rect 19444 30954 19472 31606
rect 19628 31346 19656 31878
rect 19616 31340 19668 31346
rect 19616 31282 19668 31288
rect 19812 31278 19840 40938
rect 19800 31272 19852 31278
rect 19800 31214 19852 31220
rect 19444 30926 19564 30954
rect 19432 30864 19484 30870
rect 19432 30806 19484 30812
rect 19248 30320 19300 30326
rect 19248 30262 19300 30268
rect 19340 30320 19392 30326
rect 19340 30262 19392 30268
rect 19248 29708 19300 29714
rect 19248 29650 19300 29656
rect 19260 29034 19288 29650
rect 19248 29028 19300 29034
rect 19248 28970 19300 28976
rect 19260 28558 19288 28970
rect 19248 28552 19300 28558
rect 19248 28494 19300 28500
rect 19352 28218 19380 30262
rect 19444 29170 19472 30806
rect 19536 30394 19564 30926
rect 19524 30388 19576 30394
rect 19524 30330 19576 30336
rect 19800 30116 19852 30122
rect 19800 30058 19852 30064
rect 19524 29776 19576 29782
rect 19524 29718 19576 29724
rect 19432 29164 19484 29170
rect 19432 29106 19484 29112
rect 19340 28212 19392 28218
rect 19340 28154 19392 28160
rect 18972 28076 19024 28082
rect 18972 28018 19024 28024
rect 18984 27878 19012 28018
rect 18972 27872 19024 27878
rect 18972 27814 19024 27820
rect 19064 27872 19116 27878
rect 19064 27814 19116 27820
rect 18696 22432 18748 22438
rect 18696 22374 18748 22380
rect 18880 22432 18932 22438
rect 18880 22374 18932 22380
rect 18708 21554 18736 22374
rect 18880 22092 18932 22098
rect 18880 22034 18932 22040
rect 18788 21888 18840 21894
rect 18788 21830 18840 21836
rect 18696 21548 18748 21554
rect 18696 21490 18748 21496
rect 18708 20942 18736 21490
rect 18800 21350 18828 21830
rect 18892 21554 18920 22034
rect 18880 21548 18932 21554
rect 18880 21490 18932 21496
rect 18788 21344 18840 21350
rect 18788 21286 18840 21292
rect 18984 20992 19012 27814
rect 19076 27538 19104 27814
rect 19064 27532 19116 27538
rect 19064 27474 19116 27480
rect 19064 27328 19116 27334
rect 19064 27270 19116 27276
rect 19076 26994 19104 27270
rect 19064 26988 19116 26994
rect 19064 26930 19116 26936
rect 19352 26926 19380 28154
rect 19340 26920 19392 26926
rect 19340 26862 19392 26868
rect 19064 26852 19116 26858
rect 19064 26794 19116 26800
rect 18800 20964 19012 20992
rect 18696 20936 18748 20942
rect 18696 20878 18748 20884
rect 18604 20596 18656 20602
rect 18604 20538 18656 20544
rect 18616 19990 18644 20538
rect 18708 20466 18736 20878
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 18604 19984 18656 19990
rect 18604 19926 18656 19932
rect 18524 19774 18736 19802
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 18512 19440 18564 19446
rect 18512 19382 18564 19388
rect 18420 19372 18472 19378
rect 18420 19314 18472 19320
rect 18524 19242 18552 19382
rect 18420 19236 18472 19242
rect 18420 19178 18472 19184
rect 18512 19236 18564 19242
rect 18512 19178 18564 19184
rect 18328 18760 18380 18766
rect 18328 18702 18380 18708
rect 17972 18426 18000 18566
rect 18156 18550 18368 18578
rect 18340 18426 18368 18550
rect 17960 18420 18012 18426
rect 17960 18362 18012 18368
rect 18236 18420 18288 18426
rect 18236 18362 18288 18368
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 17960 18284 18012 18290
rect 17960 18226 18012 18232
rect 18144 18284 18196 18290
rect 18144 18226 18196 18232
rect 17868 18148 17920 18154
rect 17868 18090 17920 18096
rect 17972 17814 18000 18226
rect 17960 17808 18012 17814
rect 17960 17750 18012 17756
rect 17868 17740 17920 17746
rect 17868 17682 17920 17688
rect 17880 17270 17908 17682
rect 17972 17270 18000 17750
rect 18052 17672 18104 17678
rect 18156 17660 18184 18226
rect 18248 17678 18276 18362
rect 18432 18290 18460 19178
rect 18512 18828 18564 18834
rect 18512 18770 18564 18776
rect 18420 18284 18472 18290
rect 18420 18226 18472 18232
rect 18328 18148 18380 18154
rect 18328 18090 18380 18096
rect 18104 17632 18184 17660
rect 18236 17672 18288 17678
rect 18052 17614 18104 17620
rect 18236 17614 18288 17620
rect 18052 17332 18104 17338
rect 18052 17274 18104 17280
rect 18144 17332 18196 17338
rect 18144 17274 18196 17280
rect 17868 17264 17920 17270
rect 17868 17206 17920 17212
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 17687 17156 17816 17184
rect 17687 16980 17715 17156
rect 17687 16952 17724 16980
rect 17590 16294 17592 16346
rect 17644 16294 17646 16346
rect 17590 15258 17646 16294
rect 17696 15502 17724 16952
rect 17776 16584 17828 16590
rect 17776 16526 17828 16532
rect 17684 15496 17736 15502
rect 17684 15438 17736 15444
rect 17590 15206 17592 15258
rect 17644 15206 17646 15258
rect 17590 14170 17646 15206
rect 17788 15162 17816 16526
rect 18064 16402 18092 17274
rect 17880 16374 18092 16402
rect 17880 15570 17908 16374
rect 18052 16244 18104 16250
rect 18052 16186 18104 16192
rect 18064 16046 18092 16186
rect 18052 16040 18104 16046
rect 18052 15982 18104 15988
rect 18156 15892 18184 17274
rect 18236 16584 18288 16590
rect 18236 16526 18288 16532
rect 18064 15864 18184 15892
rect 17960 15700 18012 15706
rect 17960 15642 18012 15648
rect 17972 15570 18000 15642
rect 17868 15564 17920 15570
rect 17868 15506 17920 15512
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 17880 14890 17908 15506
rect 17868 14884 17920 14890
rect 17868 14826 17920 14832
rect 17684 14816 17736 14822
rect 17684 14758 17736 14764
rect 17590 14118 17592 14170
rect 17644 14118 17646 14170
rect 17500 13252 17552 13258
rect 17500 13194 17552 13200
rect 17590 13082 17646 14118
rect 17696 13734 17724 14758
rect 17684 13728 17736 13734
rect 17684 13670 17736 13676
rect 17776 13524 17828 13530
rect 17776 13466 17828 13472
rect 17788 13274 17816 13466
rect 17590 13030 17592 13082
rect 17644 13030 17646 13082
rect 17500 12776 17552 12782
rect 17500 12718 17552 12724
rect 17512 11830 17540 12718
rect 17590 11994 17646 13030
rect 17590 11942 17592 11994
rect 17644 11942 17646 11994
rect 17500 11824 17552 11830
rect 17500 11766 17552 11772
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 17512 11218 17540 11494
rect 17500 11212 17552 11218
rect 17500 11154 17552 11160
rect 17500 11008 17552 11014
rect 17500 10950 17552 10956
rect 17512 10674 17540 10950
rect 17590 10906 17646 11942
rect 17696 13246 17816 13274
rect 17696 11762 17724 13246
rect 17880 13240 17908 14826
rect 17960 13252 18012 13258
rect 17880 13212 17960 13240
rect 17960 13194 18012 13200
rect 17868 12844 17920 12850
rect 17868 12786 17920 12792
rect 17776 12368 17828 12374
rect 17776 12310 17828 12316
rect 17684 11756 17736 11762
rect 17684 11698 17736 11704
rect 17696 11286 17724 11698
rect 17684 11280 17736 11286
rect 17684 11222 17736 11228
rect 17590 10854 17592 10906
rect 17644 10854 17646 10906
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17590 9818 17646 10854
rect 17684 10600 17736 10606
rect 17684 10542 17736 10548
rect 17590 9766 17592 9818
rect 17644 9766 17646 9818
rect 17500 9580 17552 9586
rect 17500 9522 17552 9528
rect 17512 8974 17540 9522
rect 17500 8968 17552 8974
rect 17500 8910 17552 8916
rect 17512 8566 17540 8910
rect 17590 8730 17646 9766
rect 17590 8678 17592 8730
rect 17644 8678 17646 8730
rect 17500 8560 17552 8566
rect 17500 8502 17552 8508
rect 17500 7812 17552 7818
rect 17500 7754 17552 7760
rect 17512 1222 17540 7754
rect 17590 7642 17646 8678
rect 17696 7886 17724 10542
rect 17788 9586 17816 12310
rect 17880 11762 17908 12786
rect 17960 12436 18012 12442
rect 17960 12378 18012 12384
rect 17868 11756 17920 11762
rect 17868 11698 17920 11704
rect 17972 11014 18000 12378
rect 18064 11200 18092 15864
rect 18144 15156 18196 15162
rect 18144 15098 18196 15104
rect 18156 14958 18184 15098
rect 18144 14952 18196 14958
rect 18144 14894 18196 14900
rect 18248 14532 18276 16526
rect 18340 15706 18368 18090
rect 18524 15910 18552 18770
rect 18616 18358 18644 19654
rect 18708 18952 18736 19774
rect 18692 18924 18736 18952
rect 18692 18714 18720 18924
rect 18800 18834 18828 20964
rect 18972 20868 19024 20874
rect 18972 20810 19024 20816
rect 18880 20596 18932 20602
rect 18880 20538 18932 20544
rect 18892 19922 18920 20538
rect 18984 20466 19012 20810
rect 18972 20460 19024 20466
rect 18972 20402 19024 20408
rect 18880 19916 18932 19922
rect 18880 19858 18932 19864
rect 18972 19916 19024 19922
rect 18972 19858 19024 19864
rect 18880 19236 18932 19242
rect 18880 19178 18932 19184
rect 18788 18828 18840 18834
rect 18788 18770 18840 18776
rect 18692 18686 18736 18714
rect 18604 18352 18656 18358
rect 18604 18294 18656 18300
rect 18708 17338 18736 18686
rect 18892 18086 18920 19178
rect 18984 18902 19012 19858
rect 18972 18896 19024 18902
rect 18972 18838 19024 18844
rect 18880 18080 18932 18086
rect 18880 18022 18932 18028
rect 18984 17882 19012 18838
rect 18972 17876 19024 17882
rect 18972 17818 19024 17824
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 18696 17332 18748 17338
rect 18696 17274 18748 17280
rect 18880 17196 18932 17202
rect 18880 17138 18932 17144
rect 18892 16998 18920 17138
rect 18880 16992 18932 16998
rect 18880 16934 18932 16940
rect 18880 16652 18932 16658
rect 18880 16594 18932 16600
rect 18604 16448 18656 16454
rect 18604 16390 18656 16396
rect 18512 15904 18564 15910
rect 18512 15846 18564 15852
rect 18328 15700 18380 15706
rect 18328 15642 18380 15648
rect 18512 15020 18564 15026
rect 18512 14962 18564 14968
rect 18328 14884 18380 14890
rect 18328 14826 18380 14832
rect 18156 14504 18276 14532
rect 18156 14006 18184 14504
rect 18340 14464 18368 14826
rect 18248 14436 18368 14464
rect 18248 14278 18276 14436
rect 18236 14272 18288 14278
rect 18236 14214 18288 14220
rect 18144 14000 18196 14006
rect 18144 13942 18196 13948
rect 18328 13728 18380 13734
rect 18328 13670 18380 13676
rect 18340 13530 18368 13670
rect 18328 13524 18380 13530
rect 18328 13466 18380 13472
rect 18144 13456 18196 13462
rect 18144 13398 18196 13404
rect 18156 13258 18184 13398
rect 18144 13252 18196 13258
rect 18144 13194 18196 13200
rect 18144 12844 18196 12850
rect 18144 12786 18196 12792
rect 18156 12442 18184 12786
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 18328 12164 18380 12170
rect 18328 12106 18380 12112
rect 18340 11744 18368 12106
rect 18420 12096 18472 12102
rect 18524 12084 18552 14962
rect 18616 12918 18644 16390
rect 18892 16114 18920 16594
rect 18880 16108 18932 16114
rect 18880 16050 18932 16056
rect 18696 15564 18748 15570
rect 18696 15506 18748 15512
rect 18708 14550 18736 15506
rect 18788 15496 18840 15502
rect 18788 15438 18840 15444
rect 18696 14544 18748 14550
rect 18696 14486 18748 14492
rect 18696 14340 18748 14346
rect 18696 14282 18748 14288
rect 18708 13734 18736 14282
rect 18696 13728 18748 13734
rect 18696 13670 18748 13676
rect 18800 13326 18828 15438
rect 18880 15020 18932 15026
rect 18880 14962 18932 14968
rect 18788 13320 18840 13326
rect 18788 13262 18840 13268
rect 18604 12912 18656 12918
rect 18604 12854 18656 12860
rect 18472 12056 18736 12084
rect 18420 12038 18472 12044
rect 18340 11716 18644 11744
rect 18512 11620 18564 11626
rect 18512 11562 18564 11568
rect 18328 11212 18380 11218
rect 18064 11172 18184 11200
rect 17868 11008 17920 11014
rect 17868 10950 17920 10956
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 17880 10810 17908 10950
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 17972 10742 18000 10950
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 17972 10588 18000 10678
rect 17880 10560 18000 10588
rect 17880 9586 17908 10560
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 17868 9580 17920 9586
rect 17868 9522 17920 9528
rect 17776 9444 17828 9450
rect 17776 9386 17828 9392
rect 17788 9178 17816 9386
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17880 8974 17908 9522
rect 17960 9376 18012 9382
rect 17960 9318 18012 9324
rect 17972 9178 18000 9318
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17960 8356 18012 8362
rect 17960 8298 18012 8304
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 17590 7590 17592 7642
rect 17644 7590 17646 7642
rect 17590 6554 17646 7590
rect 17696 7410 17724 7822
rect 17972 7478 18000 8298
rect 17960 7472 18012 7478
rect 17960 7414 18012 7420
rect 17684 7404 17736 7410
rect 17684 7346 17736 7352
rect 17776 6996 17828 7002
rect 17776 6938 17828 6944
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 17590 6502 17592 6554
rect 17644 6502 17646 6554
rect 17590 5466 17646 6502
rect 17696 6322 17724 6734
rect 17684 6316 17736 6322
rect 17684 6258 17736 6264
rect 17590 5414 17592 5466
rect 17644 5414 17646 5466
rect 17590 4378 17646 5414
rect 17684 4548 17736 4554
rect 17684 4490 17736 4496
rect 17590 4326 17592 4378
rect 17644 4326 17646 4378
rect 17590 3290 17646 4326
rect 17696 4282 17724 4490
rect 17684 4276 17736 4282
rect 17684 4218 17736 4224
rect 17684 3936 17736 3942
rect 17684 3878 17736 3884
rect 17590 3238 17592 3290
rect 17644 3238 17646 3290
rect 17590 2202 17646 3238
rect 17696 3194 17724 3878
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 17590 2150 17592 2202
rect 17644 2150 17646 2202
rect 17500 1216 17552 1222
rect 17500 1158 17552 1164
rect 17590 1114 17646 2150
rect 17696 1766 17724 3130
rect 17788 2854 17816 6938
rect 17972 6882 18000 7414
rect 17880 6854 18000 6882
rect 17880 6798 17908 6854
rect 17868 6792 17920 6798
rect 17868 6734 17920 6740
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 17972 6458 18000 6734
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 17868 6248 17920 6254
rect 17868 6190 17920 6196
rect 17960 6248 18012 6254
rect 17960 6190 18012 6196
rect 17880 5642 17908 6190
rect 17972 6118 18000 6190
rect 17960 6112 18012 6118
rect 17960 6054 18012 6060
rect 17972 5778 18000 6054
rect 17960 5772 18012 5778
rect 17960 5714 18012 5720
rect 17868 5636 17920 5642
rect 17868 5578 17920 5584
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 17880 3534 17908 4082
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17880 2922 17908 3470
rect 17868 2916 17920 2922
rect 17868 2858 17920 2864
rect 17776 2848 17828 2854
rect 17776 2790 17828 2796
rect 17776 2304 17828 2310
rect 17776 2246 17828 2252
rect 17868 2304 17920 2310
rect 17868 2246 17920 2252
rect 17788 1970 17816 2246
rect 17880 2038 17908 2246
rect 17868 2032 17920 2038
rect 17868 1974 17920 1980
rect 17776 1964 17828 1970
rect 17776 1906 17828 1912
rect 17684 1760 17736 1766
rect 17684 1702 17736 1708
rect 17696 1426 17724 1702
rect 17684 1420 17736 1426
rect 17684 1362 17736 1368
rect 17972 1358 18000 5510
rect 18064 4826 18092 10950
rect 18156 9518 18184 11172
rect 18328 11154 18380 11160
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 18144 9512 18196 9518
rect 18144 9454 18196 9460
rect 18144 9376 18196 9382
rect 18144 9318 18196 9324
rect 18156 8906 18184 9318
rect 18248 9110 18276 11086
rect 18340 10266 18368 11154
rect 18524 11082 18552 11562
rect 18512 11076 18564 11082
rect 18512 11018 18564 11024
rect 18420 10804 18472 10810
rect 18420 10746 18472 10752
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18340 10062 18368 10202
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18432 9586 18460 10746
rect 18512 10192 18564 10198
rect 18512 10134 18564 10140
rect 18420 9580 18472 9586
rect 18420 9522 18472 9528
rect 18524 9518 18552 10134
rect 18616 10062 18644 11716
rect 18604 10056 18656 10062
rect 18604 9998 18656 10004
rect 18708 9518 18736 12056
rect 18512 9512 18564 9518
rect 18512 9454 18564 9460
rect 18696 9512 18748 9518
rect 18696 9454 18748 9460
rect 18236 9104 18288 9110
rect 18236 9046 18288 9052
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 18512 8968 18564 8974
rect 18512 8910 18564 8916
rect 18144 8900 18196 8906
rect 18144 8842 18196 8848
rect 18248 8498 18276 8910
rect 18328 8832 18380 8838
rect 18328 8774 18380 8780
rect 18236 8492 18288 8498
rect 18236 8434 18288 8440
rect 18340 7410 18368 8774
rect 18524 8362 18552 8910
rect 18696 8560 18748 8566
rect 18696 8502 18748 8508
rect 18512 8356 18564 8362
rect 18512 8298 18564 8304
rect 18708 7478 18736 8502
rect 18800 8090 18828 13262
rect 18892 8566 18920 14962
rect 18984 12374 19012 17478
rect 18972 12368 19024 12374
rect 18972 12310 19024 12316
rect 18972 12164 19024 12170
rect 18972 12106 19024 12112
rect 18984 11830 19012 12106
rect 18972 11824 19024 11830
rect 18972 11766 19024 11772
rect 19076 10742 19104 26794
rect 19444 25974 19472 29106
rect 19536 28150 19564 29718
rect 19524 28144 19576 28150
rect 19524 28086 19576 28092
rect 19432 25968 19484 25974
rect 19432 25910 19484 25916
rect 19536 25906 19564 28086
rect 19812 28014 19840 30058
rect 19800 28008 19852 28014
rect 19800 27950 19852 27956
rect 19708 26920 19760 26926
rect 19708 26862 19760 26868
rect 19904 26874 19932 42162
rect 20260 41132 20312 41138
rect 20260 41074 20312 41080
rect 20076 39296 20128 39302
rect 20076 39238 20128 39244
rect 20088 38282 20116 39238
rect 20076 38276 20128 38282
rect 20076 38218 20128 38224
rect 19984 37256 20036 37262
rect 19984 37198 20036 37204
rect 19996 36922 20024 37198
rect 19984 36916 20036 36922
rect 19984 36858 20036 36864
rect 19984 36168 20036 36174
rect 19984 36110 20036 36116
rect 19996 35494 20024 36110
rect 19984 35488 20036 35494
rect 19984 35430 20036 35436
rect 20168 35080 20220 35086
rect 20168 35022 20220 35028
rect 20076 34944 20128 34950
rect 20076 34886 20128 34892
rect 20088 34746 20116 34886
rect 20076 34740 20128 34746
rect 20076 34682 20128 34688
rect 19984 34672 20036 34678
rect 19984 34614 20036 34620
rect 19996 32570 20024 34614
rect 20180 33998 20208 35022
rect 20168 33992 20220 33998
rect 20168 33934 20220 33940
rect 20180 33658 20208 33934
rect 20168 33652 20220 33658
rect 20168 33594 20220 33600
rect 20168 33312 20220 33318
rect 20168 33254 20220 33260
rect 19984 32564 20036 32570
rect 19984 32506 20036 32512
rect 19996 30870 20024 32506
rect 20180 32366 20208 33254
rect 20168 32360 20220 32366
rect 20168 32302 20220 32308
rect 20272 31754 20300 41074
rect 20456 38962 20484 42162
rect 22742 41914 22798 42480
rect 23020 42084 23072 42090
rect 23020 42026 23072 42032
rect 22742 41862 22744 41914
rect 22796 41862 22798 41914
rect 21640 41608 21692 41614
rect 21640 41550 21692 41556
rect 21272 41132 21324 41138
rect 21272 41074 21324 41080
rect 21088 40928 21140 40934
rect 21088 40870 21140 40876
rect 20720 40520 20772 40526
rect 20720 40462 20772 40468
rect 20628 39364 20680 39370
rect 20628 39306 20680 39312
rect 20444 38956 20496 38962
rect 20444 38898 20496 38904
rect 20640 38894 20668 39306
rect 20628 38888 20680 38894
rect 20628 38830 20680 38836
rect 20536 37868 20588 37874
rect 20536 37810 20588 37816
rect 20548 37466 20576 37810
rect 20536 37460 20588 37466
rect 20536 37402 20588 37408
rect 20352 34944 20404 34950
rect 20352 34886 20404 34892
rect 20364 32978 20392 34886
rect 20640 34678 20668 38830
rect 20628 34672 20680 34678
rect 20628 34614 20680 34620
rect 20536 34400 20588 34406
rect 20536 34342 20588 34348
rect 20548 32978 20576 34342
rect 20628 33448 20680 33454
rect 20628 33390 20680 33396
rect 20352 32972 20404 32978
rect 20352 32914 20404 32920
rect 20536 32972 20588 32978
rect 20536 32914 20588 32920
rect 20444 32836 20496 32842
rect 20444 32778 20496 32784
rect 20352 32428 20404 32434
rect 20352 32370 20404 32376
rect 20364 32026 20392 32370
rect 20352 32020 20404 32026
rect 20352 31962 20404 31968
rect 20272 31726 20392 31754
rect 20260 31680 20312 31686
rect 20260 31622 20312 31628
rect 20272 31346 20300 31622
rect 20260 31340 20312 31346
rect 20260 31282 20312 31288
rect 19984 30864 20036 30870
rect 19984 30806 20036 30812
rect 20076 30116 20128 30122
rect 20076 30058 20128 30064
rect 20088 27878 20116 30058
rect 20260 28960 20312 28966
rect 20260 28902 20312 28908
rect 20272 28694 20300 28902
rect 20260 28688 20312 28694
rect 20260 28630 20312 28636
rect 20168 28484 20220 28490
rect 20168 28426 20220 28432
rect 20076 27872 20128 27878
rect 20076 27814 20128 27820
rect 20088 27470 20116 27814
rect 20076 27464 20128 27470
rect 20076 27406 20128 27412
rect 19984 27396 20036 27402
rect 19984 27338 20036 27344
rect 19996 27062 20024 27338
rect 19984 27056 20036 27062
rect 19984 26998 20036 27004
rect 20076 26988 20128 26994
rect 20076 26930 20128 26936
rect 19720 26450 19748 26862
rect 19904 26846 20024 26874
rect 19892 26784 19944 26790
rect 19892 26726 19944 26732
rect 19708 26444 19760 26450
rect 19708 26386 19760 26392
rect 19904 26314 19932 26726
rect 19892 26308 19944 26314
rect 19892 26250 19944 26256
rect 19524 25900 19576 25906
rect 19524 25842 19576 25848
rect 19432 25832 19484 25838
rect 19432 25774 19484 25780
rect 19444 25294 19472 25774
rect 19524 25492 19576 25498
rect 19524 25434 19576 25440
rect 19432 25288 19484 25294
rect 19432 25230 19484 25236
rect 19248 24948 19300 24954
rect 19248 24890 19300 24896
rect 19156 24608 19208 24614
rect 19156 24550 19208 24556
rect 19168 24342 19196 24550
rect 19260 24342 19288 24890
rect 19444 24818 19472 25230
rect 19432 24812 19484 24818
rect 19432 24754 19484 24760
rect 19156 24336 19208 24342
rect 19156 24278 19208 24284
rect 19248 24336 19300 24342
rect 19248 24278 19300 24284
rect 19340 24064 19392 24070
rect 19536 24018 19564 25434
rect 19708 25288 19760 25294
rect 19708 25230 19760 25236
rect 19720 24818 19748 25230
rect 19708 24812 19760 24818
rect 19708 24754 19760 24760
rect 19800 24744 19852 24750
rect 19800 24686 19852 24692
rect 19340 24006 19392 24012
rect 19352 23118 19380 24006
rect 19444 23990 19564 24018
rect 19444 23322 19472 23990
rect 19524 23860 19576 23866
rect 19524 23802 19576 23808
rect 19432 23316 19484 23322
rect 19432 23258 19484 23264
rect 19248 23112 19300 23118
rect 19248 23054 19300 23060
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 19156 21888 19208 21894
rect 19156 21830 19208 21836
rect 19168 21622 19196 21830
rect 19156 21616 19208 21622
rect 19156 21558 19208 21564
rect 19260 21486 19288 23054
rect 19536 22642 19564 23802
rect 19812 22982 19840 24686
rect 19892 23792 19944 23798
rect 19892 23734 19944 23740
rect 19904 23322 19932 23734
rect 19892 23316 19944 23322
rect 19892 23258 19944 23264
rect 19996 23050 20024 26846
rect 20088 26042 20116 26930
rect 20076 26036 20128 26042
rect 20076 25978 20128 25984
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 19984 23044 20036 23050
rect 19984 22986 20036 22992
rect 19800 22976 19852 22982
rect 19800 22918 19852 22924
rect 19812 22642 19840 22918
rect 19892 22772 19944 22778
rect 19892 22714 19944 22720
rect 19432 22636 19484 22642
rect 19432 22578 19484 22584
rect 19524 22636 19576 22642
rect 19524 22578 19576 22584
rect 19800 22636 19852 22642
rect 19800 22578 19852 22584
rect 19340 22568 19392 22574
rect 19340 22510 19392 22516
rect 19352 21622 19380 22510
rect 19444 22234 19472 22578
rect 19708 22568 19760 22574
rect 19708 22510 19760 22516
rect 19524 22432 19576 22438
rect 19524 22374 19576 22380
rect 19616 22432 19668 22438
rect 19616 22374 19668 22380
rect 19432 22228 19484 22234
rect 19432 22170 19484 22176
rect 19340 21616 19392 21622
rect 19340 21558 19392 21564
rect 19248 21480 19300 21486
rect 19248 21422 19300 21428
rect 19156 20868 19208 20874
rect 19156 20810 19208 20816
rect 19168 19922 19196 20810
rect 19260 19990 19288 21422
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19340 20800 19392 20806
rect 19340 20742 19392 20748
rect 19248 19984 19300 19990
rect 19248 19926 19300 19932
rect 19156 19916 19208 19922
rect 19156 19858 19208 19864
rect 19156 19372 19208 19378
rect 19156 19314 19208 19320
rect 19168 17338 19196 19314
rect 19260 18834 19288 19926
rect 19352 18952 19380 20742
rect 19444 19378 19472 20878
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19536 19310 19564 22374
rect 19628 22098 19656 22374
rect 19616 22092 19668 22098
rect 19616 22034 19668 22040
rect 19628 20874 19656 22034
rect 19616 20868 19668 20874
rect 19616 20810 19668 20816
rect 19616 20528 19668 20534
rect 19616 20470 19668 20476
rect 19628 19514 19656 20470
rect 19616 19508 19668 19514
rect 19616 19450 19668 19456
rect 19524 19304 19576 19310
rect 19524 19246 19576 19252
rect 19352 18924 19472 18952
rect 19248 18828 19300 18834
rect 19248 18770 19300 18776
rect 19340 18624 19392 18630
rect 19340 18566 19392 18572
rect 19248 18420 19300 18426
rect 19248 18362 19300 18368
rect 19260 18086 19288 18362
rect 19352 18290 19380 18566
rect 19340 18284 19392 18290
rect 19340 18226 19392 18232
rect 19248 18080 19300 18086
rect 19248 18022 19300 18028
rect 19340 18080 19392 18086
rect 19340 18022 19392 18028
rect 19156 17332 19208 17338
rect 19156 17274 19208 17280
rect 19156 16652 19208 16658
rect 19156 16594 19208 16600
rect 19168 16182 19196 16594
rect 19156 16176 19208 16182
rect 19156 16118 19208 16124
rect 19260 15434 19288 18022
rect 19352 17542 19380 18022
rect 19340 17536 19392 17542
rect 19340 17478 19392 17484
rect 19248 15428 19300 15434
rect 19248 15370 19300 15376
rect 19444 14414 19472 18924
rect 19524 18692 19576 18698
rect 19524 18634 19576 18640
rect 19536 18426 19564 18634
rect 19524 18420 19576 18426
rect 19524 18362 19576 18368
rect 19720 17082 19748 22510
rect 19812 22030 19840 22578
rect 19800 22024 19852 22030
rect 19800 21966 19852 21972
rect 19904 21672 19932 22714
rect 19812 21644 19932 21672
rect 19812 18086 19840 21644
rect 19892 21548 19944 21554
rect 19892 21490 19944 21496
rect 19800 18080 19852 18086
rect 19800 18022 19852 18028
rect 19800 17808 19852 17814
rect 19800 17750 19852 17756
rect 19812 17270 19840 17750
rect 19800 17264 19852 17270
rect 19800 17206 19852 17212
rect 19628 17054 19748 17082
rect 19524 16584 19576 16590
rect 19524 16526 19576 16532
rect 19536 15706 19564 16526
rect 19524 15700 19576 15706
rect 19524 15642 19576 15648
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19156 13320 19208 13326
rect 19156 13262 19208 13268
rect 19168 12918 19196 13262
rect 19260 13190 19288 14010
rect 19340 13524 19392 13530
rect 19536 13512 19564 15302
rect 19392 13484 19564 13512
rect 19340 13466 19392 13472
rect 19432 13388 19484 13394
rect 19352 13348 19432 13376
rect 19248 13184 19300 13190
rect 19248 13126 19300 13132
rect 19156 12912 19208 12918
rect 19156 12854 19208 12860
rect 19352 12442 19380 13348
rect 19432 13330 19484 13336
rect 19340 12436 19392 12442
rect 19340 12378 19392 12384
rect 19156 12232 19208 12238
rect 19156 12174 19208 12180
rect 19168 11694 19196 12174
rect 19156 11688 19208 11694
rect 19156 11630 19208 11636
rect 19628 11014 19656 17054
rect 19800 16516 19852 16522
rect 19800 16458 19852 16464
rect 19708 15496 19760 15502
rect 19708 15438 19760 15444
rect 19720 12238 19748 15438
rect 19812 13462 19840 16458
rect 19904 15706 19932 21490
rect 20088 20534 20116 24142
rect 20180 21894 20208 28426
rect 20260 25152 20312 25158
rect 20260 25094 20312 25100
rect 20272 24342 20300 25094
rect 20260 24336 20312 24342
rect 20260 24278 20312 24284
rect 20260 24132 20312 24138
rect 20260 24074 20312 24080
rect 20272 23730 20300 24074
rect 20260 23724 20312 23730
rect 20260 23666 20312 23672
rect 20168 21888 20220 21894
rect 20168 21830 20220 21836
rect 20076 20528 20128 20534
rect 20076 20470 20128 20476
rect 19984 20392 20036 20398
rect 19984 20334 20036 20340
rect 19996 20058 20024 20334
rect 20076 20256 20128 20262
rect 20076 20198 20128 20204
rect 19984 20052 20036 20058
rect 19984 19994 20036 20000
rect 19996 19854 20024 19994
rect 19984 19848 20036 19854
rect 19984 19790 20036 19796
rect 20088 19786 20116 20198
rect 20076 19780 20128 19786
rect 20076 19722 20128 19728
rect 19984 17672 20036 17678
rect 19984 17614 20036 17620
rect 19996 17338 20024 17614
rect 19984 17332 20036 17338
rect 19984 17274 20036 17280
rect 19984 17196 20036 17202
rect 19984 17138 20036 17144
rect 19892 15700 19944 15706
rect 19892 15642 19944 15648
rect 19904 14822 19932 15642
rect 19996 15502 20024 17138
rect 20088 16454 20116 19722
rect 20180 19310 20208 21830
rect 20272 20806 20300 23666
rect 20364 20992 20392 31726
rect 20456 31414 20484 32778
rect 20640 32366 20668 33390
rect 20732 33318 20760 40462
rect 20996 39500 21048 39506
rect 20996 39442 21048 39448
rect 20904 38820 20956 38826
rect 20904 38762 20956 38768
rect 20916 38214 20944 38762
rect 21008 38282 21036 39442
rect 20996 38276 21048 38282
rect 20996 38218 21048 38224
rect 20904 38208 20956 38214
rect 20904 38150 20956 38156
rect 21008 37262 21036 38218
rect 20996 37256 21048 37262
rect 20996 37198 21048 37204
rect 20904 36916 20956 36922
rect 20904 36858 20956 36864
rect 20812 36168 20864 36174
rect 20812 36110 20864 36116
rect 20824 35834 20852 36110
rect 20812 35828 20864 35834
rect 20812 35770 20864 35776
rect 20916 35698 20944 36858
rect 20904 35692 20956 35698
rect 20904 35634 20956 35640
rect 21008 35578 21036 37198
rect 20824 35550 21036 35578
rect 20824 35222 20852 35550
rect 20812 35216 20864 35222
rect 20812 35158 20864 35164
rect 20824 34134 20852 35158
rect 20904 35148 20956 35154
rect 20904 35090 20956 35096
rect 20916 34610 20944 35090
rect 20904 34604 20956 34610
rect 20904 34546 20956 34552
rect 20812 34128 20864 34134
rect 20812 34070 20864 34076
rect 20720 33312 20772 33318
rect 20720 33254 20772 33260
rect 20628 32360 20680 32366
rect 20628 32302 20680 32308
rect 20720 32224 20772 32230
rect 20720 32166 20772 32172
rect 20996 32224 21048 32230
rect 20996 32166 21048 32172
rect 20732 31822 20760 32166
rect 20720 31816 20772 31822
rect 20720 31758 20772 31764
rect 20444 31408 20496 31414
rect 20444 31350 20496 31356
rect 20536 31340 20588 31346
rect 20536 31282 20588 31288
rect 20444 30388 20496 30394
rect 20444 30330 20496 30336
rect 20456 29510 20484 30330
rect 20444 29504 20496 29510
rect 20444 29446 20496 29452
rect 20444 23520 20496 23526
rect 20444 23462 20496 23468
rect 20456 21622 20484 23462
rect 20548 22574 20576 31282
rect 20628 30660 20680 30666
rect 20628 30602 20680 30608
rect 20640 30394 20668 30602
rect 20628 30388 20680 30394
rect 20628 30330 20680 30336
rect 20628 30048 20680 30054
rect 20628 29990 20680 29996
rect 20640 29850 20668 29990
rect 20628 29844 20680 29850
rect 20628 29786 20680 29792
rect 20732 29646 20760 31758
rect 21008 31346 21036 32166
rect 21100 31754 21128 40870
rect 21180 39432 21232 39438
rect 21180 39374 21232 39380
rect 21192 38010 21220 39374
rect 21180 38004 21232 38010
rect 21180 37946 21232 37952
rect 21192 36922 21220 37946
rect 21180 36916 21232 36922
rect 21180 36858 21232 36864
rect 21192 36786 21220 36858
rect 21180 36780 21232 36786
rect 21180 36722 21232 36728
rect 21180 36576 21232 36582
rect 21180 36518 21232 36524
rect 21192 35630 21220 36518
rect 21180 35624 21232 35630
rect 21180 35566 21232 35572
rect 21180 35080 21232 35086
rect 21180 35022 21232 35028
rect 21192 34542 21220 35022
rect 21180 34536 21232 34542
rect 21180 34478 21232 34484
rect 21192 33522 21220 34478
rect 21180 33516 21232 33522
rect 21180 33458 21232 33464
rect 21180 32768 21232 32774
rect 21180 32710 21232 32716
rect 21192 32502 21220 32710
rect 21180 32496 21232 32502
rect 21180 32438 21232 32444
rect 21180 32360 21232 32366
rect 21180 32302 21232 32308
rect 21192 32026 21220 32302
rect 21180 32020 21232 32026
rect 21180 31962 21232 31968
rect 21100 31726 21220 31754
rect 21088 31680 21140 31686
rect 21088 31622 21140 31628
rect 20996 31340 21048 31346
rect 20996 31282 21048 31288
rect 20812 30252 20864 30258
rect 20812 30194 20864 30200
rect 20824 29850 20852 30194
rect 20996 30184 21048 30190
rect 20996 30126 21048 30132
rect 21008 29850 21036 30126
rect 20812 29844 20864 29850
rect 20812 29786 20864 29792
rect 20996 29844 21048 29850
rect 20996 29786 21048 29792
rect 20904 29776 20956 29782
rect 20824 29724 20904 29730
rect 20824 29718 20956 29724
rect 20824 29702 20944 29718
rect 20720 29640 20772 29646
rect 20720 29582 20772 29588
rect 20720 28756 20772 28762
rect 20720 28698 20772 28704
rect 20732 27470 20760 28698
rect 20720 27464 20772 27470
rect 20720 27406 20772 27412
rect 20732 26994 20760 27406
rect 20720 26988 20772 26994
rect 20720 26930 20772 26936
rect 20824 26926 20852 29702
rect 20904 29572 20956 29578
rect 21100 29560 21128 31622
rect 20956 29532 21128 29560
rect 20904 29514 20956 29520
rect 20996 29300 21048 29306
rect 20996 29242 21048 29248
rect 21008 29034 21036 29242
rect 20996 29028 21048 29034
rect 20996 28970 21048 28976
rect 21008 27554 21036 28970
rect 21192 28966 21220 31726
rect 21180 28960 21232 28966
rect 21180 28902 21232 28908
rect 21180 28552 21232 28558
rect 21180 28494 21232 28500
rect 21088 28076 21140 28082
rect 21088 28018 21140 28024
rect 21100 27674 21128 28018
rect 21192 28014 21220 28494
rect 21284 28098 21312 41074
rect 21652 41070 21680 41550
rect 21824 41540 21876 41546
rect 21824 41482 21876 41488
rect 21640 41064 21692 41070
rect 21640 41006 21692 41012
rect 21652 39302 21680 41006
rect 21836 40050 21864 41482
rect 22284 41268 22336 41274
rect 22284 41210 22336 41216
rect 22296 40526 22324 41210
rect 22742 40826 22798 41862
rect 22836 41064 22888 41070
rect 22836 41006 22888 41012
rect 22742 40774 22744 40826
rect 22796 40774 22798 40826
rect 22284 40520 22336 40526
rect 22284 40462 22336 40468
rect 22192 40452 22244 40458
rect 22192 40394 22244 40400
rect 22008 40384 22060 40390
rect 22008 40326 22060 40332
rect 21824 40044 21876 40050
rect 21824 39986 21876 39992
rect 21640 39296 21692 39302
rect 21640 39238 21692 39244
rect 21548 39024 21600 39030
rect 21548 38966 21600 38972
rect 21560 37262 21588 38966
rect 21652 38350 21680 39238
rect 21916 38820 21968 38826
rect 21916 38762 21968 38768
rect 21640 38344 21692 38350
rect 21640 38286 21692 38292
rect 21548 37256 21600 37262
rect 21548 37198 21600 37204
rect 21364 36644 21416 36650
rect 21364 36586 21416 36592
rect 21376 35086 21404 36586
rect 21548 36032 21600 36038
rect 21548 35974 21600 35980
rect 21560 35698 21588 35974
rect 21548 35692 21600 35698
rect 21548 35634 21600 35640
rect 21652 35630 21680 38286
rect 21732 37324 21784 37330
rect 21732 37266 21784 37272
rect 21744 35698 21772 37266
rect 21928 36582 21956 38762
rect 21916 36576 21968 36582
rect 21916 36518 21968 36524
rect 21916 36100 21968 36106
rect 21916 36042 21968 36048
rect 21732 35692 21784 35698
rect 21732 35634 21784 35640
rect 21640 35624 21692 35630
rect 21640 35566 21692 35572
rect 21548 35556 21600 35562
rect 21548 35498 21600 35504
rect 21456 35216 21508 35222
rect 21456 35158 21508 35164
rect 21364 35080 21416 35086
rect 21364 35022 21416 35028
rect 21364 33992 21416 33998
rect 21364 33934 21416 33940
rect 21376 33386 21404 33934
rect 21364 33380 21416 33386
rect 21364 33322 21416 33328
rect 21364 32360 21416 32366
rect 21364 32302 21416 32308
rect 21376 31686 21404 32302
rect 21364 31680 21416 31686
rect 21364 31622 21416 31628
rect 21376 29782 21404 31622
rect 21364 29776 21416 29782
rect 21364 29718 21416 29724
rect 21284 28070 21404 28098
rect 21180 28008 21232 28014
rect 21180 27950 21232 27956
rect 21088 27668 21140 27674
rect 21088 27610 21140 27616
rect 21008 27526 21128 27554
rect 20904 27396 20956 27402
rect 20904 27338 20956 27344
rect 20812 26920 20864 26926
rect 20812 26862 20864 26868
rect 20812 26376 20864 26382
rect 20812 26318 20864 26324
rect 20628 25900 20680 25906
rect 20628 25842 20680 25848
rect 20640 25362 20668 25842
rect 20628 25356 20680 25362
rect 20628 25298 20680 25304
rect 20824 24274 20852 26318
rect 20916 25430 20944 27338
rect 20996 26988 21048 26994
rect 20996 26930 21048 26936
rect 21008 26586 21036 26930
rect 21100 26790 21128 27526
rect 21192 26926 21220 27950
rect 21272 27940 21324 27946
rect 21272 27882 21324 27888
rect 21284 27606 21312 27882
rect 21272 27600 21324 27606
rect 21272 27542 21324 27548
rect 21180 26920 21232 26926
rect 21180 26862 21232 26868
rect 21088 26784 21140 26790
rect 21088 26726 21140 26732
rect 20996 26580 21048 26586
rect 20996 26522 21048 26528
rect 20904 25424 20956 25430
rect 20904 25366 20956 25372
rect 20916 24698 20944 25366
rect 20996 25152 21048 25158
rect 20996 25094 21048 25100
rect 21008 24818 21036 25094
rect 21100 24818 21128 26726
rect 21192 26246 21220 26862
rect 21180 26240 21232 26246
rect 21180 26182 21232 26188
rect 21192 25906 21220 26182
rect 21180 25900 21232 25906
rect 21180 25842 21232 25848
rect 20996 24812 21048 24818
rect 20996 24754 21048 24760
rect 21088 24812 21140 24818
rect 21088 24754 21140 24760
rect 20916 24670 21036 24698
rect 20904 24608 20956 24614
rect 20904 24550 20956 24556
rect 20812 24268 20864 24274
rect 20812 24210 20864 24216
rect 20720 23792 20772 23798
rect 20720 23734 20772 23740
rect 20824 23746 20852 24210
rect 20916 24206 20944 24550
rect 20904 24200 20956 24206
rect 20904 24142 20956 24148
rect 20628 23724 20680 23730
rect 20628 23666 20680 23672
rect 20536 22568 20588 22574
rect 20536 22510 20588 22516
rect 20444 21616 20496 21622
rect 20444 21558 20496 21564
rect 20640 21146 20668 23666
rect 20732 23168 20760 23734
rect 20824 23718 20944 23746
rect 20916 23186 20944 23718
rect 20904 23180 20956 23186
rect 20732 23140 20852 23168
rect 20720 23044 20772 23050
rect 20720 22986 20772 22992
rect 20732 22778 20760 22986
rect 20720 22772 20772 22778
rect 20720 22714 20772 22720
rect 20628 21140 20680 21146
rect 20628 21082 20680 21088
rect 20720 21140 20772 21146
rect 20720 21082 20772 21088
rect 20364 20964 20576 20992
rect 20444 20868 20496 20874
rect 20444 20810 20496 20816
rect 20260 20800 20312 20806
rect 20260 20742 20312 20748
rect 20260 20324 20312 20330
rect 20260 20266 20312 20272
rect 20168 19304 20220 19310
rect 20168 19246 20220 19252
rect 20272 18358 20300 20266
rect 20352 19848 20404 19854
rect 20352 19790 20404 19796
rect 20364 19378 20392 19790
rect 20352 19372 20404 19378
rect 20352 19314 20404 19320
rect 20260 18352 20312 18358
rect 20260 18294 20312 18300
rect 20364 18222 20392 19314
rect 20260 18216 20312 18222
rect 20260 18158 20312 18164
rect 20352 18216 20404 18222
rect 20352 18158 20404 18164
rect 20168 18080 20220 18086
rect 20168 18022 20220 18028
rect 20180 17678 20208 18022
rect 20168 17672 20220 17678
rect 20168 17614 20220 17620
rect 20180 17066 20208 17614
rect 20168 17060 20220 17066
rect 20168 17002 20220 17008
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 20272 16250 20300 18158
rect 20352 17536 20404 17542
rect 20352 17478 20404 17484
rect 20364 17202 20392 17478
rect 20352 17196 20404 17202
rect 20352 17138 20404 17144
rect 20260 16244 20312 16250
rect 20260 16186 20312 16192
rect 20272 16114 20300 16186
rect 20260 16108 20312 16114
rect 20260 16050 20312 16056
rect 20272 15502 20300 16050
rect 20364 15570 20392 17138
rect 20352 15564 20404 15570
rect 20352 15506 20404 15512
rect 19984 15496 20036 15502
rect 20260 15496 20312 15502
rect 20036 15456 20116 15484
rect 19984 15438 20036 15444
rect 19892 14816 19944 14822
rect 19892 14758 19944 14764
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 19892 13932 19944 13938
rect 19892 13874 19944 13880
rect 19800 13456 19852 13462
rect 19800 13398 19852 13404
rect 19812 12646 19840 13398
rect 19904 12918 19932 13874
rect 19996 13394 20024 14010
rect 19984 13388 20036 13394
rect 19984 13330 20036 13336
rect 19892 12912 19944 12918
rect 19892 12854 19944 12860
rect 19800 12640 19852 12646
rect 19800 12582 19852 12588
rect 20088 12238 20116 15456
rect 20260 15438 20312 15444
rect 20272 15094 20300 15438
rect 20260 15088 20312 15094
rect 20260 15030 20312 15036
rect 20456 13002 20484 20810
rect 20548 14226 20576 20964
rect 20732 20618 20760 21082
rect 20824 20806 20852 23140
rect 20904 23122 20956 23128
rect 20904 22636 20956 22642
rect 20904 22578 20956 22584
rect 20916 22030 20944 22578
rect 21008 22522 21036 24670
rect 21284 23882 21312 27542
rect 21192 23854 21312 23882
rect 21088 23180 21140 23186
rect 21088 23122 21140 23128
rect 21100 22642 21128 23122
rect 21192 22778 21220 23854
rect 21272 23792 21324 23798
rect 21272 23734 21324 23740
rect 21180 22772 21232 22778
rect 21180 22714 21232 22720
rect 21088 22636 21140 22642
rect 21088 22578 21140 22584
rect 21008 22494 21128 22522
rect 20996 22092 21048 22098
rect 20996 22034 21048 22040
rect 20904 22024 20956 22030
rect 20904 21966 20956 21972
rect 20904 21888 20956 21894
rect 20904 21830 20956 21836
rect 20916 21418 20944 21830
rect 21008 21690 21036 22034
rect 20996 21684 21048 21690
rect 20996 21626 21048 21632
rect 20904 21412 20956 21418
rect 20904 21354 20956 21360
rect 21008 20942 21036 21626
rect 20996 20936 21048 20942
rect 20996 20878 21048 20884
rect 20812 20800 20864 20806
rect 20812 20742 20864 20748
rect 20640 20590 20760 20618
rect 20640 20262 20668 20590
rect 20720 20460 20772 20466
rect 20720 20402 20772 20408
rect 20628 20256 20680 20262
rect 20628 20198 20680 20204
rect 20628 19780 20680 19786
rect 20628 19722 20680 19728
rect 20640 17542 20668 19722
rect 20732 18630 20760 20402
rect 20720 18624 20772 18630
rect 20720 18566 20772 18572
rect 20628 17536 20680 17542
rect 20628 17478 20680 17484
rect 20640 14414 20668 17478
rect 20720 17128 20772 17134
rect 20720 17070 20772 17076
rect 20732 14822 20760 17070
rect 20824 15502 20852 20742
rect 20996 20392 21048 20398
rect 20996 20334 21048 20340
rect 21008 18834 21036 20334
rect 20996 18828 21048 18834
rect 20996 18770 21048 18776
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 20916 17134 20944 18702
rect 20996 18284 21048 18290
rect 20996 18226 21048 18232
rect 21008 17882 21036 18226
rect 20996 17876 21048 17882
rect 20996 17818 21048 17824
rect 20904 17128 20956 17134
rect 20904 17070 20956 17076
rect 20996 16720 21048 16726
rect 20996 16662 21048 16668
rect 20904 16652 20956 16658
rect 20904 16594 20956 16600
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 20916 15026 20944 16594
rect 21008 15910 21036 16662
rect 20996 15904 21048 15910
rect 20996 15846 21048 15852
rect 21008 15162 21036 15846
rect 20996 15156 21048 15162
rect 20996 15098 21048 15104
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 20628 14408 20680 14414
rect 20628 14350 20680 14356
rect 20548 14198 20668 14226
rect 20180 12986 20484 13002
rect 20168 12980 20484 12986
rect 20220 12974 20484 12980
rect 20168 12922 20220 12928
rect 20536 12844 20588 12850
rect 20536 12786 20588 12792
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 20444 12776 20496 12782
rect 20444 12718 20496 12724
rect 20272 12238 20300 12718
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 19708 12232 19760 12238
rect 19708 12174 19760 12180
rect 20076 12232 20128 12238
rect 20076 12174 20128 12180
rect 20260 12232 20312 12238
rect 20260 12174 20312 12180
rect 20168 11824 20220 11830
rect 20168 11766 20220 11772
rect 19616 11008 19668 11014
rect 19616 10950 19668 10956
rect 19064 10736 19116 10742
rect 19064 10678 19116 10684
rect 19432 10736 19484 10742
rect 19432 10678 19484 10684
rect 19340 10600 19392 10606
rect 19340 10542 19392 10548
rect 19352 9994 19380 10542
rect 19340 9988 19392 9994
rect 19340 9930 19392 9936
rect 19352 9586 19380 9930
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19156 9512 19208 9518
rect 19156 9454 19208 9460
rect 19064 9444 19116 9450
rect 19064 9386 19116 9392
rect 18880 8560 18932 8566
rect 18880 8502 18932 8508
rect 18788 8084 18840 8090
rect 18788 8026 18840 8032
rect 18696 7472 18748 7478
rect 18696 7414 18748 7420
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 18328 7404 18380 7410
rect 18328 7346 18380 7352
rect 18156 6458 18184 7346
rect 18144 6452 18196 6458
rect 18144 6394 18196 6400
rect 18156 5166 18184 6394
rect 18236 5296 18288 5302
rect 18236 5238 18288 5244
rect 18420 5296 18472 5302
rect 18420 5238 18472 5244
rect 18144 5160 18196 5166
rect 18144 5102 18196 5108
rect 18052 4820 18104 4826
rect 18052 4762 18104 4768
rect 18156 2446 18184 5102
rect 18248 3618 18276 5238
rect 18328 4684 18380 4690
rect 18432 4672 18460 5238
rect 18788 5024 18840 5030
rect 18788 4966 18840 4972
rect 18604 4684 18656 4690
rect 18380 4644 18460 4672
rect 18524 4644 18604 4672
rect 18328 4626 18380 4632
rect 18328 4548 18380 4554
rect 18328 4490 18380 4496
rect 18340 4282 18368 4490
rect 18328 4276 18380 4282
rect 18328 4218 18380 4224
rect 18248 3602 18368 3618
rect 18248 3596 18380 3602
rect 18248 3590 18328 3596
rect 18328 3538 18380 3544
rect 18420 3392 18472 3398
rect 18420 3334 18472 3340
rect 18236 2848 18288 2854
rect 18236 2790 18288 2796
rect 18144 2440 18196 2446
rect 18144 2382 18196 2388
rect 18156 2038 18184 2382
rect 18144 2032 18196 2038
rect 18144 1974 18196 1980
rect 18248 1358 18276 2790
rect 18432 2446 18460 3334
rect 18420 2440 18472 2446
rect 18524 2428 18552 4644
rect 18604 4626 18656 4632
rect 18800 4146 18828 4966
rect 18972 4208 19024 4214
rect 18972 4150 19024 4156
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 18788 4140 18840 4146
rect 18788 4082 18840 4088
rect 18616 3466 18644 4082
rect 18696 3528 18748 3534
rect 18696 3470 18748 3476
rect 18604 3460 18656 3466
rect 18604 3402 18656 3408
rect 18616 3058 18644 3402
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18708 2650 18736 3470
rect 18696 2644 18748 2650
rect 18696 2586 18748 2592
rect 18604 2440 18656 2446
rect 18524 2400 18604 2428
rect 18420 2382 18472 2388
rect 18604 2382 18656 2388
rect 18328 1964 18380 1970
rect 18328 1906 18380 1912
rect 18340 1562 18368 1906
rect 18616 1562 18644 2382
rect 18328 1556 18380 1562
rect 18328 1498 18380 1504
rect 18604 1556 18656 1562
rect 18604 1498 18656 1504
rect 18708 1358 18736 2586
rect 18800 2514 18828 4082
rect 18984 2990 19012 4150
rect 18972 2984 19024 2990
rect 18972 2926 19024 2932
rect 18788 2508 18840 2514
rect 18788 2450 18840 2456
rect 17960 1352 18012 1358
rect 17960 1294 18012 1300
rect 18236 1352 18288 1358
rect 18236 1294 18288 1300
rect 18696 1352 18748 1358
rect 18696 1294 18748 1300
rect 19076 1222 19104 9386
rect 19168 8498 19196 9454
rect 19444 8922 19472 10678
rect 19524 9920 19576 9926
rect 19524 9862 19576 9868
rect 19536 9450 19564 9862
rect 19524 9444 19576 9450
rect 19524 9386 19576 9392
rect 19616 9376 19668 9382
rect 19616 9318 19668 9324
rect 19628 9042 19656 9318
rect 19708 9104 19760 9110
rect 19708 9046 19760 9052
rect 19616 9036 19668 9042
rect 19616 8978 19668 8984
rect 19720 8974 19748 9046
rect 20180 8974 20208 11766
rect 20364 11762 20392 12582
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 20456 11558 20484 12718
rect 20548 12442 20576 12786
rect 20536 12436 20588 12442
rect 20536 12378 20588 12384
rect 20536 12232 20588 12238
rect 20536 12174 20588 12180
rect 20444 11552 20496 11558
rect 20444 11494 20496 11500
rect 20548 11506 20576 12174
rect 20640 11694 20668 14198
rect 21008 14074 21036 15098
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 20996 13728 21048 13734
rect 20996 13670 21048 13676
rect 21008 13394 21036 13670
rect 20996 13388 21048 13394
rect 20996 13330 21048 13336
rect 20720 12980 20772 12986
rect 20720 12922 20772 12928
rect 20732 12374 20760 12922
rect 20812 12640 20864 12646
rect 20812 12582 20864 12588
rect 20720 12368 20772 12374
rect 20720 12310 20772 12316
rect 20628 11688 20680 11694
rect 20628 11630 20680 11636
rect 20628 11552 20680 11558
rect 20548 11500 20628 11506
rect 20548 11494 20680 11500
rect 20456 11218 20484 11494
rect 20548 11478 20668 11494
rect 20444 11212 20496 11218
rect 20444 11154 20496 11160
rect 20456 10470 20484 11154
rect 20640 10742 20668 11478
rect 20824 11218 20852 12582
rect 20904 12436 20956 12442
rect 20904 12378 20956 12384
rect 20812 11212 20864 11218
rect 20812 11154 20864 11160
rect 20628 10736 20680 10742
rect 20628 10678 20680 10684
rect 20444 10464 20496 10470
rect 20444 10406 20496 10412
rect 20824 10130 20852 11154
rect 20916 11150 20944 12378
rect 20904 11144 20956 11150
rect 20904 11086 20956 11092
rect 20916 10810 20944 11086
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 20812 10124 20864 10130
rect 20812 10066 20864 10072
rect 21100 10062 21128 22494
rect 21180 21888 21232 21894
rect 21180 21830 21232 21836
rect 21192 19378 21220 21830
rect 21284 21146 21312 23734
rect 21272 21140 21324 21146
rect 21272 21082 21324 21088
rect 21272 20052 21324 20058
rect 21272 19994 21324 20000
rect 21180 19372 21232 19378
rect 21180 19314 21232 19320
rect 21180 18964 21232 18970
rect 21180 18906 21232 18912
rect 21192 18290 21220 18906
rect 21180 18284 21232 18290
rect 21180 18226 21232 18232
rect 21284 16250 21312 19994
rect 21376 18290 21404 28070
rect 21468 23746 21496 35158
rect 21560 33590 21588 35498
rect 21640 35488 21692 35494
rect 21640 35430 21692 35436
rect 21652 35086 21680 35430
rect 21640 35080 21692 35086
rect 21640 35022 21692 35028
rect 21640 34740 21692 34746
rect 21640 34682 21692 34688
rect 21548 33584 21600 33590
rect 21548 33526 21600 33532
rect 21548 33380 21600 33386
rect 21548 33322 21600 33328
rect 21560 31958 21588 33322
rect 21548 31952 21600 31958
rect 21548 31894 21600 31900
rect 21548 31816 21600 31822
rect 21548 31758 21600 31764
rect 21560 31482 21588 31758
rect 21548 31476 21600 31482
rect 21548 31418 21600 31424
rect 21548 29640 21600 29646
rect 21548 29582 21600 29588
rect 21560 28762 21588 29582
rect 21548 28756 21600 28762
rect 21548 28698 21600 28704
rect 21548 28008 21600 28014
rect 21548 27950 21600 27956
rect 21560 24138 21588 27950
rect 21652 26450 21680 34682
rect 21744 34202 21772 35634
rect 21732 34196 21784 34202
rect 21732 34138 21784 34144
rect 21928 33658 21956 36042
rect 22020 35578 22048 40326
rect 22204 40118 22232 40394
rect 22192 40112 22244 40118
rect 22192 40054 22244 40060
rect 22204 39982 22232 40054
rect 22192 39976 22244 39982
rect 22192 39918 22244 39924
rect 22204 39658 22232 39918
rect 22468 39840 22520 39846
rect 22468 39782 22520 39788
rect 22204 39630 22324 39658
rect 22296 38962 22324 39630
rect 22284 38956 22336 38962
rect 22284 38898 22336 38904
rect 22284 38752 22336 38758
rect 22284 38694 22336 38700
rect 22100 38276 22152 38282
rect 22100 38218 22152 38224
rect 22112 38010 22140 38218
rect 22100 38004 22152 38010
rect 22100 37946 22152 37952
rect 22296 37874 22324 38694
rect 22480 37874 22508 39782
rect 22742 39738 22798 40774
rect 22848 40730 22876 41006
rect 22836 40724 22888 40730
rect 22836 40666 22888 40672
rect 23032 40594 23060 42026
rect 23572 42016 23624 42022
rect 23572 41958 23624 41964
rect 23664 42016 23716 42022
rect 23664 41958 23716 41964
rect 23584 41682 23612 41958
rect 23572 41676 23624 41682
rect 23572 41618 23624 41624
rect 23296 41540 23348 41546
rect 23296 41482 23348 41488
rect 23308 40730 23336 41482
rect 23572 41472 23624 41478
rect 23572 41414 23624 41420
rect 23584 41002 23612 41414
rect 23572 40996 23624 41002
rect 23572 40938 23624 40944
rect 23296 40724 23348 40730
rect 23296 40666 23348 40672
rect 23676 40610 23704 41958
rect 24400 41608 24452 41614
rect 24400 41550 24452 41556
rect 23848 41472 23900 41478
rect 23848 41414 23900 41420
rect 23756 40928 23808 40934
rect 23756 40870 23808 40876
rect 23020 40588 23072 40594
rect 23020 40530 23072 40536
rect 23584 40582 23704 40610
rect 23032 40050 23060 40530
rect 23584 40526 23612 40582
rect 23768 40526 23796 40870
rect 23480 40520 23532 40526
rect 23480 40462 23532 40468
rect 23572 40520 23624 40526
rect 23572 40462 23624 40468
rect 23756 40520 23808 40526
rect 23756 40462 23808 40468
rect 23492 40186 23520 40462
rect 23480 40180 23532 40186
rect 23480 40122 23532 40128
rect 22836 40044 22888 40050
rect 22836 39986 22888 39992
rect 23020 40044 23072 40050
rect 23020 39986 23072 39992
rect 23296 40044 23348 40050
rect 23296 39986 23348 39992
rect 22742 39686 22744 39738
rect 22796 39686 22798 39738
rect 22742 38650 22798 39686
rect 22848 39642 22876 39986
rect 22928 39976 22980 39982
rect 22928 39918 22980 39924
rect 22836 39636 22888 39642
rect 22836 39578 22888 39584
rect 22940 39030 22968 39918
rect 23032 39438 23060 39986
rect 23308 39438 23336 39986
rect 23584 39846 23612 40462
rect 23664 39976 23716 39982
rect 23664 39918 23716 39924
rect 23572 39840 23624 39846
rect 23572 39782 23624 39788
rect 23584 39574 23612 39782
rect 23572 39568 23624 39574
rect 23572 39510 23624 39516
rect 23020 39432 23072 39438
rect 23020 39374 23072 39380
rect 23296 39432 23348 39438
rect 23348 39380 23428 39386
rect 23296 39374 23428 39380
rect 22928 39024 22980 39030
rect 22928 38966 22980 38972
rect 22742 38598 22744 38650
rect 22796 38598 22798 38650
rect 22284 37868 22336 37874
rect 22284 37810 22336 37816
rect 22468 37868 22520 37874
rect 22468 37810 22520 37816
rect 22742 37562 22798 38598
rect 22940 38554 22968 38966
rect 23032 38962 23060 39374
rect 23308 39358 23428 39374
rect 23296 39092 23348 39098
rect 23296 39034 23348 39040
rect 23020 38956 23072 38962
rect 23020 38898 23072 38904
rect 22928 38548 22980 38554
rect 22928 38490 22980 38496
rect 22940 37942 22968 38490
rect 22928 37936 22980 37942
rect 22928 37878 22980 37884
rect 22928 37800 22980 37806
rect 22928 37742 22980 37748
rect 22742 37510 22744 37562
rect 22796 37510 22798 37562
rect 22652 36780 22704 36786
rect 22652 36722 22704 36728
rect 22376 36712 22428 36718
rect 22376 36654 22428 36660
rect 22192 36372 22244 36378
rect 22192 36314 22244 36320
rect 22204 36088 22232 36314
rect 22284 36100 22336 36106
rect 22204 36060 22284 36088
rect 22020 35550 22140 35578
rect 22112 35290 22140 35550
rect 22008 35284 22060 35290
rect 22008 35226 22060 35232
rect 22100 35284 22152 35290
rect 22100 35226 22152 35232
rect 22020 33930 22048 35226
rect 22204 35170 22232 36060
rect 22284 36042 22336 36048
rect 22388 35494 22416 36654
rect 22664 36174 22692 36722
rect 22742 36474 22798 37510
rect 22742 36422 22744 36474
rect 22796 36422 22798 36474
rect 22560 36168 22612 36174
rect 22560 36110 22612 36116
rect 22652 36168 22704 36174
rect 22652 36110 22704 36116
rect 22376 35488 22428 35494
rect 22376 35430 22428 35436
rect 22112 35142 22232 35170
rect 22008 33924 22060 33930
rect 22008 33866 22060 33872
rect 22112 33862 22140 35142
rect 22284 35012 22336 35018
rect 22284 34954 22336 34960
rect 22192 34468 22244 34474
rect 22192 34410 22244 34416
rect 22204 33998 22232 34410
rect 22192 33992 22244 33998
rect 22192 33934 22244 33940
rect 22100 33856 22152 33862
rect 22100 33798 22152 33804
rect 21916 33652 21968 33658
rect 21916 33594 21968 33600
rect 22100 33448 22152 33454
rect 22100 33390 22152 33396
rect 22008 33312 22060 33318
rect 22008 33254 22060 33260
rect 21732 33040 21784 33046
rect 21732 32982 21784 32988
rect 21744 32910 21772 32982
rect 21824 32972 21876 32978
rect 21824 32914 21876 32920
rect 21732 32904 21784 32910
rect 21732 32846 21784 32852
rect 21744 31822 21772 32846
rect 21732 31816 21784 31822
rect 21732 31758 21784 31764
rect 21836 31482 21864 32914
rect 21916 32836 21968 32842
rect 21916 32778 21968 32784
rect 21928 32366 21956 32778
rect 21916 32360 21968 32366
rect 21916 32302 21968 32308
rect 21916 32224 21968 32230
rect 21916 32166 21968 32172
rect 21824 31476 21876 31482
rect 21824 31418 21876 31424
rect 21732 31408 21784 31414
rect 21732 31350 21784 31356
rect 21744 30870 21772 31350
rect 21732 30864 21784 30870
rect 21732 30806 21784 30812
rect 21928 30716 21956 32166
rect 21744 30688 21956 30716
rect 21744 27402 21772 30688
rect 21824 30592 21876 30598
rect 21824 30534 21876 30540
rect 21732 27396 21784 27402
rect 21732 27338 21784 27344
rect 21836 26994 21864 30534
rect 21916 29572 21968 29578
rect 21916 29514 21968 29520
rect 21928 29306 21956 29514
rect 21916 29300 21968 29306
rect 21916 29242 21968 29248
rect 21916 28620 21968 28626
rect 21916 28562 21968 28568
rect 21928 27470 21956 28562
rect 22020 28422 22048 33254
rect 22112 32434 22140 33390
rect 22100 32428 22152 32434
rect 22100 32370 22152 32376
rect 22100 31476 22152 31482
rect 22100 31418 22152 31424
rect 22112 31142 22140 31418
rect 22100 31136 22152 31142
rect 22100 31078 22152 31084
rect 22100 30932 22152 30938
rect 22100 30874 22152 30880
rect 22112 30258 22140 30874
rect 22204 30802 22232 33934
rect 22296 33318 22324 34954
rect 22468 34604 22520 34610
rect 22468 34546 22520 34552
rect 22376 34400 22428 34406
rect 22376 34342 22428 34348
rect 22388 33998 22416 34342
rect 22376 33992 22428 33998
rect 22376 33934 22428 33940
rect 22376 33856 22428 33862
rect 22376 33798 22428 33804
rect 22284 33312 22336 33318
rect 22284 33254 22336 33260
rect 22388 33130 22416 33798
rect 22296 33102 22416 33130
rect 22192 30796 22244 30802
rect 22192 30738 22244 30744
rect 22192 30660 22244 30666
rect 22192 30602 22244 30608
rect 22204 30394 22232 30602
rect 22192 30388 22244 30394
rect 22192 30330 22244 30336
rect 22100 30252 22152 30258
rect 22100 30194 22152 30200
rect 22100 30116 22152 30122
rect 22100 30058 22152 30064
rect 22008 28416 22060 28422
rect 22008 28358 22060 28364
rect 21916 27464 21968 27470
rect 21916 27406 21968 27412
rect 21824 26988 21876 26994
rect 21824 26930 21876 26936
rect 21640 26444 21692 26450
rect 21640 26386 21692 26392
rect 21652 25838 21680 26386
rect 21732 26376 21784 26382
rect 21836 26330 21864 26930
rect 21784 26324 21864 26330
rect 21732 26318 21864 26324
rect 21744 26302 21864 26318
rect 21836 26042 21864 26302
rect 21824 26036 21876 26042
rect 21824 25978 21876 25984
rect 21640 25832 21692 25838
rect 21640 25774 21692 25780
rect 21652 25226 21680 25774
rect 22112 25294 22140 30058
rect 22192 29504 22244 29510
rect 22192 29446 22244 29452
rect 22204 29306 22232 29446
rect 22192 29300 22244 29306
rect 22192 29242 22244 29248
rect 22192 28960 22244 28966
rect 22192 28902 22244 28908
rect 22204 26790 22232 28902
rect 22192 26784 22244 26790
rect 22192 26726 22244 26732
rect 22192 25832 22244 25838
rect 22192 25774 22244 25780
rect 22100 25288 22152 25294
rect 22100 25230 22152 25236
rect 21640 25220 21692 25226
rect 21640 25162 21692 25168
rect 22112 24818 22140 25230
rect 22204 24954 22232 25774
rect 22192 24948 22244 24954
rect 22192 24890 22244 24896
rect 22100 24812 22152 24818
rect 22100 24754 22152 24760
rect 22008 24676 22060 24682
rect 22008 24618 22060 24624
rect 21548 24132 21600 24138
rect 21548 24074 21600 24080
rect 21916 23792 21968 23798
rect 21468 23718 21588 23746
rect 21916 23734 21968 23740
rect 21456 22772 21508 22778
rect 21456 22714 21508 22720
rect 21468 20534 21496 22714
rect 21560 21026 21588 23718
rect 21928 22778 21956 23734
rect 22020 23526 22048 24618
rect 22112 24392 22140 24754
rect 22192 24404 22244 24410
rect 22112 24364 22192 24392
rect 22192 24346 22244 24352
rect 22100 23588 22152 23594
rect 22100 23530 22152 23536
rect 22008 23520 22060 23526
rect 22008 23462 22060 23468
rect 21916 22772 21968 22778
rect 21916 22714 21968 22720
rect 22008 22636 22060 22642
rect 22008 22578 22060 22584
rect 21916 21956 21968 21962
rect 21916 21898 21968 21904
rect 21824 21616 21876 21622
rect 21824 21558 21876 21564
rect 21560 20998 21680 21026
rect 21548 20936 21600 20942
rect 21548 20878 21600 20884
rect 21456 20528 21508 20534
rect 21456 20470 21508 20476
rect 21560 19310 21588 20878
rect 21652 20058 21680 20998
rect 21836 20806 21864 21558
rect 21928 21010 21956 21898
rect 22020 21690 22048 22578
rect 22112 22094 22140 23530
rect 22112 22066 22232 22094
rect 22100 22024 22152 22030
rect 22100 21966 22152 21972
rect 22008 21684 22060 21690
rect 22008 21626 22060 21632
rect 21916 21004 21968 21010
rect 21916 20946 21968 20952
rect 21824 20800 21876 20806
rect 21824 20742 21876 20748
rect 21824 20460 21876 20466
rect 21824 20402 21876 20408
rect 21732 20392 21784 20398
rect 21732 20334 21784 20340
rect 21640 20052 21692 20058
rect 21640 19994 21692 20000
rect 21548 19304 21600 19310
rect 21548 19246 21600 19252
rect 21744 18766 21772 20334
rect 21836 19514 21864 20402
rect 21928 20330 21956 20946
rect 21916 20324 21968 20330
rect 21916 20266 21968 20272
rect 22008 20256 22060 20262
rect 22008 20198 22060 20204
rect 21916 19984 21968 19990
rect 21916 19926 21968 19932
rect 21824 19508 21876 19514
rect 21824 19450 21876 19456
rect 21824 19168 21876 19174
rect 21824 19110 21876 19116
rect 21732 18760 21784 18766
rect 21732 18702 21784 18708
rect 21640 18692 21692 18698
rect 21640 18634 21692 18640
rect 21364 18284 21416 18290
rect 21364 18226 21416 18232
rect 21652 18086 21680 18634
rect 21640 18080 21692 18086
rect 21640 18022 21692 18028
rect 21272 16244 21324 16250
rect 21272 16186 21324 16192
rect 21456 16176 21508 16182
rect 21456 16118 21508 16124
rect 21272 15904 21324 15910
rect 21272 15846 21324 15852
rect 21284 15026 21312 15846
rect 21272 15020 21324 15026
rect 21272 14962 21324 14968
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 21364 14272 21416 14278
rect 21364 14214 21416 14220
rect 21192 13938 21220 14214
rect 21376 14006 21404 14214
rect 21364 14000 21416 14006
rect 21364 13942 21416 13948
rect 21180 13932 21232 13938
rect 21180 13874 21232 13880
rect 21376 13870 21404 13942
rect 21364 13864 21416 13870
rect 21364 13806 21416 13812
rect 21376 12714 21404 13806
rect 21364 12708 21416 12714
rect 21364 12650 21416 12656
rect 21468 12238 21496 16118
rect 21548 12776 21600 12782
rect 21548 12718 21600 12724
rect 21456 12232 21508 12238
rect 21456 12174 21508 12180
rect 21364 12164 21416 12170
rect 21364 12106 21416 12112
rect 21376 11830 21404 12106
rect 21364 11824 21416 11830
rect 21364 11766 21416 11772
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 21192 10674 21220 11290
rect 21180 10668 21232 10674
rect 21180 10610 21232 10616
rect 21088 10056 21140 10062
rect 21088 9998 21140 10004
rect 20536 9580 20588 9586
rect 20536 9522 20588 9528
rect 20260 9512 20312 9518
rect 20260 9454 20312 9460
rect 19708 8968 19760 8974
rect 19444 8894 19564 8922
rect 19708 8910 19760 8916
rect 20168 8968 20220 8974
rect 20168 8910 20220 8916
rect 19432 8832 19484 8838
rect 19352 8792 19432 8820
rect 19352 8786 19380 8792
rect 19306 8758 19380 8786
rect 19432 8774 19484 8780
rect 19306 8634 19334 8758
rect 19294 8628 19346 8634
rect 19294 8570 19346 8576
rect 19156 8492 19208 8498
rect 19156 8434 19208 8440
rect 19536 8412 19564 8894
rect 19352 8384 19564 8412
rect 19156 7268 19208 7274
rect 19156 7210 19208 7216
rect 19168 5846 19196 7210
rect 19248 7200 19300 7206
rect 19248 7142 19300 7148
rect 19156 5840 19208 5846
rect 19156 5782 19208 5788
rect 19156 4548 19208 4554
rect 19156 4490 19208 4496
rect 19168 4078 19196 4490
rect 19260 4078 19288 7142
rect 19352 5234 19380 8384
rect 19616 8356 19668 8362
rect 19536 8316 19616 8344
rect 19432 7812 19484 7818
rect 19432 7754 19484 7760
rect 19444 7002 19472 7754
rect 19432 6996 19484 7002
rect 19432 6938 19484 6944
rect 19536 6798 19564 8316
rect 19616 8298 19668 8304
rect 19616 7336 19668 7342
rect 19616 7278 19668 7284
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19340 5228 19392 5234
rect 19340 5170 19392 5176
rect 19340 4140 19392 4146
rect 19340 4082 19392 4088
rect 19156 4072 19208 4078
rect 19156 4014 19208 4020
rect 19248 4072 19300 4078
rect 19248 4014 19300 4020
rect 19248 3936 19300 3942
rect 19248 3878 19300 3884
rect 19260 3602 19288 3878
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19352 3534 19380 4082
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19352 2666 19380 3470
rect 19260 2638 19380 2666
rect 19260 2582 19288 2638
rect 19248 2576 19300 2582
rect 19248 2518 19300 2524
rect 19340 1352 19392 1358
rect 19340 1294 19392 1300
rect 19064 1216 19116 1222
rect 19064 1158 19116 1164
rect 17590 1062 17592 1114
rect 17644 1062 17646 1114
rect 17590 1040 17646 1062
rect 17408 1012 17460 1018
rect 17408 954 17460 960
rect 13820 944 13872 950
rect 13820 886 13872 892
rect 13832 800 13860 886
rect 19352 800 19380 1294
rect 19628 882 19656 7278
rect 19720 6866 19748 8910
rect 19984 8832 20036 8838
rect 19984 8774 20036 8780
rect 19996 8634 20024 8774
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 19800 8492 19852 8498
rect 19800 8434 19852 8440
rect 19812 7206 19840 8434
rect 20180 7886 20208 8910
rect 20272 8498 20300 9454
rect 20548 8498 20576 9522
rect 20628 9444 20680 9450
rect 20628 9386 20680 9392
rect 20260 8492 20312 8498
rect 20260 8434 20312 8440
rect 20536 8492 20588 8498
rect 20536 8434 20588 8440
rect 20640 8362 20668 9386
rect 21100 8974 21128 9998
rect 21272 9580 21324 9586
rect 21272 9522 21324 9528
rect 21284 9110 21312 9522
rect 21272 9104 21324 9110
rect 21272 9046 21324 9052
rect 21088 8968 21140 8974
rect 21088 8910 21140 8916
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20732 8498 20760 8774
rect 20720 8492 20772 8498
rect 20720 8434 20772 8440
rect 20628 8356 20680 8362
rect 20628 8298 20680 8304
rect 20732 8090 20760 8434
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 21284 7886 21312 9046
rect 20168 7880 20220 7886
rect 20168 7822 20220 7828
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 21088 7744 21140 7750
rect 21088 7686 21140 7692
rect 20628 7404 20680 7410
rect 20628 7346 20680 7352
rect 19800 7200 19852 7206
rect 19800 7142 19852 7148
rect 19708 6860 19760 6866
rect 19708 6802 19760 6808
rect 19812 6798 19840 7142
rect 19800 6792 19852 6798
rect 19800 6734 19852 6740
rect 19708 5636 19760 5642
rect 19708 5578 19760 5584
rect 19720 1222 19748 5578
rect 19812 5302 19840 6734
rect 19892 6724 19944 6730
rect 19892 6666 19944 6672
rect 19904 6458 19932 6666
rect 19892 6452 19944 6458
rect 19892 6394 19944 6400
rect 20640 5846 20668 7346
rect 20996 7336 21048 7342
rect 20996 7278 21048 7284
rect 20904 7200 20956 7206
rect 20904 7142 20956 7148
rect 20916 6186 20944 7142
rect 20904 6180 20956 6186
rect 20904 6122 20956 6128
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 20628 5840 20680 5846
rect 20628 5782 20680 5788
rect 20260 5568 20312 5574
rect 20260 5510 20312 5516
rect 19800 5296 19852 5302
rect 19800 5238 19852 5244
rect 19892 5228 19944 5234
rect 19892 5170 19944 5176
rect 19904 3738 19932 5170
rect 20272 5030 20300 5510
rect 20444 5160 20496 5166
rect 20444 5102 20496 5108
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 20260 5024 20312 5030
rect 20260 4966 20312 4972
rect 19892 3732 19944 3738
rect 19892 3674 19944 3680
rect 19800 3392 19852 3398
rect 19800 3334 19852 3340
rect 19812 3058 19840 3334
rect 19800 3052 19852 3058
rect 19800 2994 19852 3000
rect 19800 2848 19852 2854
rect 19800 2790 19852 2796
rect 19812 2378 19840 2790
rect 19800 2372 19852 2378
rect 19800 2314 19852 2320
rect 19996 1970 20024 4966
rect 20272 4690 20300 4966
rect 20260 4684 20312 4690
rect 20260 4626 20312 4632
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 20088 3194 20116 4558
rect 20168 4480 20220 4486
rect 20168 4422 20220 4428
rect 20180 4146 20208 4422
rect 20456 4282 20484 5102
rect 20640 4690 20668 5782
rect 20628 4684 20680 4690
rect 20628 4626 20680 4632
rect 20628 4548 20680 4554
rect 20628 4490 20680 4496
rect 20444 4276 20496 4282
rect 20444 4218 20496 4224
rect 20168 4140 20220 4146
rect 20168 4082 20220 4088
rect 20260 3528 20312 3534
rect 20260 3470 20312 3476
rect 20076 3188 20128 3194
rect 20076 3130 20128 3136
rect 20272 3058 20300 3470
rect 20260 3052 20312 3058
rect 20260 2994 20312 3000
rect 20456 2854 20484 4218
rect 20640 3534 20668 4490
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 20444 2848 20496 2854
rect 20444 2790 20496 2796
rect 20640 2106 20668 3470
rect 20628 2100 20680 2106
rect 20628 2042 20680 2048
rect 19984 1964 20036 1970
rect 19984 1906 20036 1912
rect 20732 1358 20760 6054
rect 21008 5114 21036 7278
rect 21100 6662 21128 7686
rect 21284 7460 21312 7822
rect 21364 7472 21416 7478
rect 21284 7432 21364 7460
rect 21364 7414 21416 7420
rect 21088 6656 21140 6662
rect 21088 6598 21140 6604
rect 21100 5302 21128 6598
rect 21088 5296 21140 5302
rect 21088 5238 21140 5244
rect 21272 5160 21324 5166
rect 21008 5086 21128 5114
rect 21272 5102 21324 5108
rect 20996 4616 21048 4622
rect 20996 4558 21048 4564
rect 21008 3738 21036 4558
rect 20996 3732 21048 3738
rect 20996 3674 21048 3680
rect 20904 3664 20956 3670
rect 20904 3606 20956 3612
rect 20916 3466 20944 3606
rect 20904 3460 20956 3466
rect 20904 3402 20956 3408
rect 20916 3058 20944 3402
rect 20904 3052 20956 3058
rect 20904 2994 20956 3000
rect 21100 2774 21128 5086
rect 21284 4826 21312 5102
rect 21272 4820 21324 4826
rect 21272 4762 21324 4768
rect 21180 4616 21232 4622
rect 21180 4558 21232 4564
rect 21192 4078 21220 4558
rect 21180 4072 21232 4078
rect 21180 4014 21232 4020
rect 21192 2904 21220 4014
rect 21468 3618 21496 12174
rect 21560 10470 21588 12718
rect 21652 12442 21680 18022
rect 21744 17882 21772 18702
rect 21836 18358 21864 19110
rect 21824 18352 21876 18358
rect 21824 18294 21876 18300
rect 21928 18222 21956 19926
rect 22020 19854 22048 20198
rect 22008 19848 22060 19854
rect 22008 19790 22060 19796
rect 22112 19786 22140 21966
rect 22204 21690 22232 22066
rect 22192 21684 22244 21690
rect 22192 21626 22244 21632
rect 22192 21344 22244 21350
rect 22192 21286 22244 21292
rect 22100 19780 22152 19786
rect 22100 19722 22152 19728
rect 22112 19378 22140 19722
rect 22100 19372 22152 19378
rect 22100 19314 22152 19320
rect 22008 19168 22060 19174
rect 22204 19122 22232 21286
rect 22296 20262 22324 33102
rect 22480 32298 22508 34546
rect 22572 33454 22600 36110
rect 22664 35222 22692 36110
rect 22742 35386 22798 36422
rect 22742 35334 22744 35386
rect 22796 35334 22798 35386
rect 22652 35216 22704 35222
rect 22652 35158 22704 35164
rect 22742 34298 22798 35334
rect 22742 34246 22744 34298
rect 22796 34246 22798 34298
rect 22560 33448 22612 33454
rect 22560 33390 22612 33396
rect 22572 32434 22600 33390
rect 22742 33210 22798 34246
rect 22940 33674 22968 37742
rect 23308 37670 23336 39034
rect 23400 38962 23428 39358
rect 23388 38956 23440 38962
rect 23388 38898 23440 38904
rect 23676 38826 23704 39918
rect 23664 38820 23716 38826
rect 23664 38762 23716 38768
rect 23676 38350 23704 38762
rect 23768 38418 23796 40462
rect 23860 40050 23888 41414
rect 24308 41064 24360 41070
rect 24308 41006 24360 41012
rect 24032 40928 24084 40934
rect 24032 40870 24084 40876
rect 24044 40594 24072 40870
rect 24032 40588 24084 40594
rect 24032 40530 24084 40536
rect 23848 40044 23900 40050
rect 23848 39986 23900 39992
rect 23860 39506 23888 39986
rect 23848 39500 23900 39506
rect 23848 39442 23900 39448
rect 24320 39438 24348 41006
rect 24412 40526 24440 41550
rect 24768 41540 24820 41546
rect 24768 41482 24820 41488
rect 24400 40520 24452 40526
rect 24400 40462 24452 40468
rect 24492 40452 24544 40458
rect 24492 40394 24544 40400
rect 24504 39642 24532 40394
rect 24584 40112 24636 40118
rect 24584 40054 24636 40060
rect 24492 39636 24544 39642
rect 24492 39578 24544 39584
rect 24596 39438 24624 40054
rect 24676 39500 24728 39506
rect 24676 39442 24728 39448
rect 24308 39432 24360 39438
rect 24308 39374 24360 39380
rect 24584 39432 24636 39438
rect 24584 39374 24636 39380
rect 24216 38752 24268 38758
rect 24216 38694 24268 38700
rect 23756 38412 23808 38418
rect 23756 38354 23808 38360
rect 23664 38344 23716 38350
rect 23664 38286 23716 38292
rect 24228 37874 24256 38694
rect 24320 37874 24348 39374
rect 24584 38956 24636 38962
rect 24584 38898 24636 38904
rect 24400 38344 24452 38350
rect 24400 38286 24452 38292
rect 24412 38010 24440 38286
rect 24492 38208 24544 38214
rect 24492 38150 24544 38156
rect 24400 38004 24452 38010
rect 24400 37946 24452 37952
rect 24504 37874 24532 38150
rect 24216 37868 24268 37874
rect 24216 37810 24268 37816
rect 24308 37868 24360 37874
rect 24308 37810 24360 37816
rect 24492 37868 24544 37874
rect 24492 37810 24544 37816
rect 23296 37664 23348 37670
rect 23296 37606 23348 37612
rect 23308 37466 23336 37606
rect 23296 37460 23348 37466
rect 23296 37402 23348 37408
rect 23480 37460 23532 37466
rect 23480 37402 23532 37408
rect 23020 37256 23072 37262
rect 23020 37198 23072 37204
rect 23032 36786 23060 37198
rect 23388 37188 23440 37194
rect 23388 37130 23440 37136
rect 23400 36854 23428 37130
rect 23388 36848 23440 36854
rect 23388 36790 23440 36796
rect 23020 36780 23072 36786
rect 23020 36722 23072 36728
rect 23492 36174 23520 37402
rect 24228 37330 24256 37810
rect 24400 37664 24452 37670
rect 24400 37606 24452 37612
rect 24216 37324 24268 37330
rect 24216 37266 24268 37272
rect 24032 37256 24084 37262
rect 24032 37198 24084 37204
rect 24044 37126 24072 37198
rect 24032 37120 24084 37126
rect 24032 37062 24084 37068
rect 24044 36718 24072 37062
rect 24032 36712 24084 36718
rect 24032 36654 24084 36660
rect 23480 36168 23532 36174
rect 23480 36110 23532 36116
rect 23204 36100 23256 36106
rect 23204 36042 23256 36048
rect 23020 35692 23072 35698
rect 23020 35634 23072 35640
rect 23032 35290 23060 35634
rect 23020 35284 23072 35290
rect 23020 35226 23072 35232
rect 23112 35216 23164 35222
rect 23112 35158 23164 35164
rect 23124 34610 23152 35158
rect 23216 35086 23244 36042
rect 23204 35080 23256 35086
rect 23204 35022 23256 35028
rect 23112 34604 23164 34610
rect 23112 34546 23164 34552
rect 23204 34536 23256 34542
rect 23204 34478 23256 34484
rect 22940 33646 23060 33674
rect 22928 33584 22980 33590
rect 22928 33526 22980 33532
rect 22836 33516 22888 33522
rect 22836 33458 22888 33464
rect 22742 33158 22744 33210
rect 22796 33158 22798 33210
rect 22560 32428 22612 32434
rect 22560 32370 22612 32376
rect 22468 32292 22520 32298
rect 22468 32234 22520 32240
rect 22742 32122 22798 33158
rect 22848 33114 22876 33458
rect 22836 33108 22888 33114
rect 22836 33050 22888 33056
rect 22940 32910 22968 33526
rect 22928 32904 22980 32910
rect 22928 32846 22980 32852
rect 22836 32768 22888 32774
rect 22836 32710 22888 32716
rect 22742 32070 22744 32122
rect 22796 32070 22798 32122
rect 22376 31952 22428 31958
rect 22428 31900 22692 31906
rect 22376 31894 22692 31900
rect 22388 31890 22692 31894
rect 22388 31884 22704 31890
rect 22388 31878 22652 31884
rect 22652 31826 22704 31832
rect 22376 31816 22428 31822
rect 22376 31758 22428 31764
rect 22388 28762 22416 31758
rect 22468 31748 22520 31754
rect 22468 31690 22520 31696
rect 22480 31414 22508 31690
rect 22468 31408 22520 31414
rect 22468 31350 22520 31356
rect 22468 31136 22520 31142
rect 22468 31078 22520 31084
rect 22480 30258 22508 31078
rect 22742 31034 22798 32070
rect 22848 31822 22876 32710
rect 23032 32586 23060 33646
rect 23216 32978 23244 34478
rect 23492 33386 23520 36110
rect 23848 36032 23900 36038
rect 23848 35974 23900 35980
rect 23860 35562 23888 35974
rect 23848 35556 23900 35562
rect 23848 35498 23900 35504
rect 23664 35080 23716 35086
rect 23664 35022 23716 35028
rect 23676 34610 23704 35022
rect 23664 34604 23716 34610
rect 23664 34546 23716 34552
rect 23572 34400 23624 34406
rect 23572 34342 23624 34348
rect 23480 33380 23532 33386
rect 23480 33322 23532 33328
rect 23296 33312 23348 33318
rect 23296 33254 23348 33260
rect 23204 32972 23256 32978
rect 23204 32914 23256 32920
rect 23032 32558 23152 32586
rect 22928 32020 22980 32026
rect 22928 31962 22980 31968
rect 22836 31816 22888 31822
rect 22836 31758 22888 31764
rect 22742 30982 22744 31034
rect 22796 30982 22798 31034
rect 22468 30252 22520 30258
rect 22468 30194 22520 30200
rect 22480 29170 22508 30194
rect 22742 29946 22798 30982
rect 22836 30184 22888 30190
rect 22836 30126 22888 30132
rect 22742 29894 22744 29946
rect 22796 29894 22798 29946
rect 22468 29164 22520 29170
rect 22468 29106 22520 29112
rect 22560 29164 22612 29170
rect 22560 29106 22612 29112
rect 22468 28960 22520 28966
rect 22468 28902 22520 28908
rect 22376 28756 22428 28762
rect 22376 28698 22428 28704
rect 22480 28626 22508 28902
rect 22468 28620 22520 28626
rect 22468 28562 22520 28568
rect 22468 28416 22520 28422
rect 22468 28358 22520 28364
rect 22480 28218 22508 28358
rect 22468 28212 22520 28218
rect 22468 28154 22520 28160
rect 22572 28082 22600 29106
rect 22652 29096 22704 29102
rect 22652 29038 22704 29044
rect 22664 28558 22692 29038
rect 22742 28858 22798 29894
rect 22848 29782 22876 30126
rect 22836 29776 22888 29782
rect 22836 29718 22888 29724
rect 22848 29288 22876 29718
rect 22940 29510 22968 31962
rect 23020 31680 23072 31686
rect 23020 31622 23072 31628
rect 22928 29504 22980 29510
rect 22928 29446 22980 29452
rect 22928 29300 22980 29306
rect 22848 29260 22928 29288
rect 22928 29242 22980 29248
rect 22742 28806 22744 28858
rect 22796 28806 22798 28858
rect 22652 28552 22704 28558
rect 22652 28494 22704 28500
rect 22560 28076 22612 28082
rect 22560 28018 22612 28024
rect 22664 28014 22692 28494
rect 22652 28008 22704 28014
rect 22652 27950 22704 27956
rect 22468 27940 22520 27946
rect 22468 27882 22520 27888
rect 22376 27464 22428 27470
rect 22376 27406 22428 27412
rect 22388 26994 22416 27406
rect 22376 26988 22428 26994
rect 22376 26930 22428 26936
rect 22480 26314 22508 27882
rect 22560 27600 22612 27606
rect 22560 27542 22612 27548
rect 22468 26308 22520 26314
rect 22468 26250 22520 26256
rect 22480 25362 22508 26250
rect 22468 25356 22520 25362
rect 22468 25298 22520 25304
rect 22572 25294 22600 27542
rect 22664 27538 22692 27950
rect 22742 27770 22798 28806
rect 22940 28694 22968 29242
rect 23032 29102 23060 31622
rect 23124 29578 23152 32558
rect 23308 32502 23336 33254
rect 23584 32978 23612 34342
rect 23676 34202 23704 34546
rect 23860 34474 23888 35498
rect 23848 34468 23900 34474
rect 23848 34410 23900 34416
rect 23664 34196 23716 34202
rect 23664 34138 23716 34144
rect 23676 33318 23704 34138
rect 23860 33522 23888 34410
rect 23848 33516 23900 33522
rect 23848 33458 23900 33464
rect 23860 33402 23888 33458
rect 23768 33374 23888 33402
rect 23664 33312 23716 33318
rect 23664 33254 23716 33260
rect 23572 32972 23624 32978
rect 23572 32914 23624 32920
rect 23664 32972 23716 32978
rect 23768 32960 23796 33374
rect 23848 33312 23900 33318
rect 23848 33254 23900 33260
rect 23716 32932 23796 32960
rect 23664 32914 23716 32920
rect 23388 32768 23440 32774
rect 23388 32710 23440 32716
rect 23296 32496 23348 32502
rect 23296 32438 23348 32444
rect 23400 31346 23428 32710
rect 23584 32434 23612 32914
rect 23860 32910 23888 33254
rect 23848 32904 23900 32910
rect 23848 32846 23900 32852
rect 23940 32836 23992 32842
rect 23940 32778 23992 32784
rect 23572 32428 23624 32434
rect 23572 32370 23624 32376
rect 23952 32298 23980 32778
rect 23940 32292 23992 32298
rect 23940 32234 23992 32240
rect 23480 32224 23532 32230
rect 23480 32166 23532 32172
rect 23492 31822 23520 32166
rect 23480 31816 23532 31822
rect 23480 31758 23532 31764
rect 24044 31686 24072 36654
rect 24124 33380 24176 33386
rect 24124 33322 24176 33328
rect 24032 31680 24084 31686
rect 24032 31622 24084 31628
rect 23848 31476 23900 31482
rect 23848 31418 23900 31424
rect 23388 31340 23440 31346
rect 23388 31282 23440 31288
rect 23664 31136 23716 31142
rect 23664 31078 23716 31084
rect 23572 30932 23624 30938
rect 23572 30874 23624 30880
rect 23112 29572 23164 29578
rect 23112 29514 23164 29520
rect 23480 29572 23532 29578
rect 23480 29514 23532 29520
rect 23112 29164 23164 29170
rect 23112 29106 23164 29112
rect 23020 29096 23072 29102
rect 23020 29038 23072 29044
rect 22928 28688 22980 28694
rect 22928 28630 22980 28636
rect 22836 28484 22888 28490
rect 22888 28444 22968 28472
rect 22836 28426 22888 28432
rect 22742 27718 22744 27770
rect 22796 27718 22798 27770
rect 22652 27532 22704 27538
rect 22652 27474 22704 27480
rect 22664 26382 22692 27474
rect 22742 26682 22798 27718
rect 22940 27554 22968 28444
rect 23032 28098 23060 29038
rect 23124 28762 23152 29106
rect 23112 28756 23164 28762
rect 23112 28698 23164 28704
rect 23124 28234 23152 28698
rect 23124 28206 23244 28234
rect 23032 28070 23141 28098
rect 23216 28082 23244 28206
rect 23113 27996 23141 28070
rect 23204 28076 23256 28082
rect 23204 28018 23256 28024
rect 23388 28008 23440 28014
rect 23113 27968 23152 27996
rect 23124 27962 23152 27968
rect 23124 27956 23388 27962
rect 23124 27950 23440 27956
rect 23124 27934 23428 27950
rect 23124 27928 23152 27934
rect 23032 27900 23152 27928
rect 23032 27674 23060 27900
rect 23020 27668 23072 27674
rect 23020 27610 23072 27616
rect 23296 27668 23348 27674
rect 23296 27610 23348 27616
rect 23204 27600 23256 27606
rect 22940 27526 23060 27554
rect 23204 27542 23256 27548
rect 22928 27464 22980 27470
rect 22928 27406 22980 27412
rect 22940 27130 22968 27406
rect 22928 27124 22980 27130
rect 22928 27066 22980 27072
rect 22836 26988 22888 26994
rect 22836 26930 22888 26936
rect 22742 26630 22744 26682
rect 22796 26630 22798 26682
rect 22652 26376 22704 26382
rect 22652 26318 22704 26324
rect 22742 25594 22798 26630
rect 22848 26246 22876 26930
rect 22940 26382 22968 27066
rect 23032 26586 23060 27526
rect 23020 26580 23072 26586
rect 23020 26522 23072 26528
rect 22928 26376 22980 26382
rect 22928 26318 22980 26324
rect 22836 26240 22888 26246
rect 22836 26182 22888 26188
rect 22742 25542 22744 25594
rect 22796 25542 22798 25594
rect 22560 25288 22612 25294
rect 22560 25230 22612 25236
rect 22468 25152 22520 25158
rect 22468 25094 22520 25100
rect 22480 24886 22508 25094
rect 22560 24948 22612 24954
rect 22560 24890 22612 24896
rect 22468 24880 22520 24886
rect 22468 24822 22520 24828
rect 22572 24750 22600 24890
rect 22652 24880 22704 24886
rect 22652 24822 22704 24828
rect 22560 24744 22612 24750
rect 22560 24686 22612 24692
rect 22664 24342 22692 24822
rect 22742 24506 22798 25542
rect 22742 24454 22744 24506
rect 22796 24454 22798 24506
rect 22652 24336 22704 24342
rect 22652 24278 22704 24284
rect 22652 24200 22704 24206
rect 22652 24142 22704 24148
rect 22468 23656 22520 23662
rect 22468 23598 22520 23604
rect 22480 22982 22508 23598
rect 22468 22976 22520 22982
rect 22468 22918 22520 22924
rect 22376 22704 22428 22710
rect 22376 22646 22428 22652
rect 22388 22030 22416 22646
rect 22376 22024 22428 22030
rect 22376 21966 22428 21972
rect 22480 21894 22508 22918
rect 22560 22160 22612 22166
rect 22560 22102 22612 22108
rect 22376 21888 22428 21894
rect 22376 21830 22428 21836
rect 22468 21888 22520 21894
rect 22468 21830 22520 21836
rect 22388 21010 22416 21830
rect 22376 21004 22428 21010
rect 22376 20946 22428 20952
rect 22480 20942 22508 21830
rect 22572 21554 22600 22102
rect 22560 21548 22612 21554
rect 22560 21490 22612 21496
rect 22468 20936 22520 20942
rect 22468 20878 22520 20884
rect 22376 20868 22428 20874
rect 22376 20810 22428 20816
rect 22284 20256 22336 20262
rect 22284 20198 22336 20204
rect 22284 20052 22336 20058
rect 22284 19994 22336 20000
rect 22008 19110 22060 19116
rect 22020 18426 22048 19110
rect 22112 19094 22232 19122
rect 22112 18426 22140 19094
rect 22192 18964 22244 18970
rect 22192 18906 22244 18912
rect 22008 18420 22060 18426
rect 22008 18362 22060 18368
rect 22100 18420 22152 18426
rect 22100 18362 22152 18368
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 21916 18216 21968 18222
rect 21916 18158 21968 18164
rect 21824 18080 21876 18086
rect 21824 18022 21876 18028
rect 21732 17876 21784 17882
rect 21732 17818 21784 17824
rect 21744 17202 21772 17818
rect 21836 17270 21864 18022
rect 21928 17678 21956 18158
rect 21916 17672 21968 17678
rect 21916 17614 21968 17620
rect 21824 17264 21876 17270
rect 21824 17206 21876 17212
rect 21732 17196 21784 17202
rect 21732 17138 21784 17144
rect 21928 16114 21956 17614
rect 22112 16998 22140 18226
rect 22204 17202 22232 18906
rect 22192 17196 22244 17202
rect 22192 17138 22244 17144
rect 22100 16992 22152 16998
rect 22152 16952 22232 16980
rect 22100 16934 22152 16940
rect 21916 16108 21968 16114
rect 21916 16050 21968 16056
rect 22100 16108 22152 16114
rect 22100 16050 22152 16056
rect 22008 15360 22060 15366
rect 22008 15302 22060 15308
rect 21824 14272 21876 14278
rect 21824 14214 21876 14220
rect 21732 14068 21784 14074
rect 21732 14010 21784 14016
rect 21744 13530 21772 14010
rect 21732 13524 21784 13530
rect 21732 13466 21784 13472
rect 21836 13326 21864 14214
rect 22020 13734 22048 15302
rect 22112 15162 22140 16050
rect 22100 15156 22152 15162
rect 22100 15098 22152 15104
rect 22204 15094 22232 16952
rect 22296 16590 22324 19994
rect 22388 18630 22416 20810
rect 22560 20324 22612 20330
rect 22560 20266 22612 20272
rect 22468 20256 22520 20262
rect 22468 20198 22520 20204
rect 22376 18624 22428 18630
rect 22376 18566 22428 18572
rect 22376 18420 22428 18426
rect 22376 18362 22428 18368
rect 22388 16794 22416 18362
rect 22376 16788 22428 16794
rect 22376 16730 22428 16736
rect 22388 16590 22416 16730
rect 22284 16584 22336 16590
rect 22284 16526 22336 16532
rect 22376 16584 22428 16590
rect 22376 16526 22428 16532
rect 22284 16448 22336 16454
rect 22284 16390 22336 16396
rect 22192 15088 22244 15094
rect 22112 15036 22192 15042
rect 22112 15030 22244 15036
rect 22112 15014 22232 15030
rect 22296 15026 22324 16390
rect 22284 15020 22336 15026
rect 22008 13728 22060 13734
rect 22008 13670 22060 13676
rect 21824 13320 21876 13326
rect 21824 13262 21876 13268
rect 21916 13184 21968 13190
rect 21916 13126 21968 13132
rect 21928 12850 21956 13126
rect 21916 12844 21968 12850
rect 21916 12786 21968 12792
rect 21640 12436 21692 12442
rect 21640 12378 21692 12384
rect 21640 11620 21692 11626
rect 21640 11562 21692 11568
rect 21548 10464 21600 10470
rect 21548 10406 21600 10412
rect 21560 9042 21588 10406
rect 21652 10062 21680 11562
rect 21916 11212 21968 11218
rect 21916 11154 21968 11160
rect 21732 11076 21784 11082
rect 21732 11018 21784 11024
rect 21640 10056 21692 10062
rect 21640 9998 21692 10004
rect 21744 9450 21772 11018
rect 21824 10464 21876 10470
rect 21824 10406 21876 10412
rect 21836 9586 21864 10406
rect 21928 10198 21956 11154
rect 21916 10192 21968 10198
rect 21916 10134 21968 10140
rect 21916 9648 21968 9654
rect 21916 9590 21968 9596
rect 21824 9580 21876 9586
rect 21824 9522 21876 9528
rect 21732 9444 21784 9450
rect 21732 9386 21784 9392
rect 21548 9036 21600 9042
rect 21548 8978 21600 8984
rect 21824 9036 21876 9042
rect 21824 8978 21876 8984
rect 21732 8492 21784 8498
rect 21732 8434 21784 8440
rect 21744 8090 21772 8434
rect 21640 8084 21692 8090
rect 21640 8026 21692 8032
rect 21732 8084 21784 8090
rect 21732 8026 21784 8032
rect 21652 7342 21680 8026
rect 21836 7970 21864 8978
rect 21744 7942 21864 7970
rect 21928 7954 21956 9590
rect 21916 7948 21968 7954
rect 21640 7336 21692 7342
rect 21640 7278 21692 7284
rect 21640 7200 21692 7206
rect 21640 7142 21692 7148
rect 21652 7002 21680 7142
rect 21640 6996 21692 7002
rect 21640 6938 21692 6944
rect 21744 6882 21772 7942
rect 21916 7890 21968 7896
rect 22020 7886 22048 13670
rect 22112 13530 22140 15014
rect 22284 14962 22336 14968
rect 22192 14952 22244 14958
rect 22192 14894 22244 14900
rect 22100 13524 22152 13530
rect 22100 13466 22152 13472
rect 22112 11626 22140 13466
rect 22100 11620 22152 11626
rect 22100 11562 22152 11568
rect 22204 11286 22232 14894
rect 22388 14414 22416 16526
rect 22376 14408 22428 14414
rect 22376 14350 22428 14356
rect 22376 13388 22428 13394
rect 22376 13330 22428 13336
rect 22388 12918 22416 13330
rect 22376 12912 22428 12918
rect 22376 12854 22428 12860
rect 22480 12434 22508 20198
rect 22572 19310 22600 20266
rect 22560 19304 22612 19310
rect 22560 19246 22612 19252
rect 22572 18086 22600 19246
rect 22560 18080 22612 18086
rect 22560 18022 22612 18028
rect 22560 17672 22612 17678
rect 22560 17614 22612 17620
rect 22572 17338 22600 17614
rect 22560 17332 22612 17338
rect 22560 17274 22612 17280
rect 22560 16448 22612 16454
rect 22560 16390 22612 16396
rect 22572 14414 22600 16390
rect 22560 14408 22612 14414
rect 22560 14350 22612 14356
rect 22572 13394 22600 14350
rect 22560 13388 22612 13394
rect 22560 13330 22612 13336
rect 22560 13252 22612 13258
rect 22560 13194 22612 13200
rect 22572 12646 22600 13194
rect 22560 12640 22612 12646
rect 22560 12582 22612 12588
rect 22388 12406 22508 12434
rect 22192 11280 22244 11286
rect 22192 11222 22244 11228
rect 22284 11076 22336 11082
rect 22284 11018 22336 11024
rect 22100 10804 22152 10810
rect 22100 10746 22152 10752
rect 22112 10674 22140 10746
rect 22296 10674 22324 11018
rect 22100 10668 22152 10674
rect 22100 10610 22152 10616
rect 22284 10668 22336 10674
rect 22284 10610 22336 10616
rect 22112 9518 22140 10610
rect 22388 10554 22416 12406
rect 22572 12238 22600 12582
rect 22560 12232 22612 12238
rect 22560 12174 22612 12180
rect 22560 11144 22612 11150
rect 22560 11086 22612 11092
rect 22468 11008 22520 11014
rect 22468 10950 22520 10956
rect 22480 10674 22508 10950
rect 22572 10810 22600 11086
rect 22560 10804 22612 10810
rect 22560 10746 22612 10752
rect 22664 10690 22692 24142
rect 22468 10668 22520 10674
rect 22468 10610 22520 10616
rect 22572 10662 22692 10690
rect 22742 23418 22798 24454
rect 22848 24206 22876 26182
rect 23216 25838 23244 27542
rect 23204 25832 23256 25838
rect 23204 25774 23256 25780
rect 23308 24818 23336 27610
rect 23388 27464 23440 27470
rect 23388 27406 23440 27412
rect 23400 27062 23428 27406
rect 23492 27130 23520 29514
rect 23584 27674 23612 30874
rect 23676 30258 23704 31078
rect 23664 30252 23716 30258
rect 23664 30194 23716 30200
rect 23664 30116 23716 30122
rect 23664 30058 23716 30064
rect 23676 29850 23704 30058
rect 23664 29844 23716 29850
rect 23664 29786 23716 29792
rect 23572 27668 23624 27674
rect 23572 27610 23624 27616
rect 23572 27328 23624 27334
rect 23572 27270 23624 27276
rect 23480 27124 23532 27130
rect 23480 27066 23532 27072
rect 23388 27056 23440 27062
rect 23388 26998 23440 27004
rect 23480 26988 23532 26994
rect 23480 26930 23532 26936
rect 23492 26586 23520 26930
rect 23480 26580 23532 26586
rect 23480 26522 23532 26528
rect 23584 25702 23612 27270
rect 23572 25696 23624 25702
rect 23572 25638 23624 25644
rect 23388 25288 23440 25294
rect 23388 25230 23440 25236
rect 23296 24812 23348 24818
rect 23296 24754 23348 24760
rect 23308 24274 23336 24754
rect 23400 24750 23428 25230
rect 23584 25158 23612 25638
rect 23572 25152 23624 25158
rect 23572 25094 23624 25100
rect 23676 24970 23704 29786
rect 23756 29504 23808 29510
rect 23756 29446 23808 29452
rect 23768 27878 23796 29446
rect 23860 28558 23888 31418
rect 23940 31340 23992 31346
rect 23940 31282 23992 31288
rect 23848 28552 23900 28558
rect 23848 28494 23900 28500
rect 23756 27872 23808 27878
rect 23756 27814 23808 27820
rect 23860 27538 23888 28494
rect 23952 28370 23980 31282
rect 24032 31272 24084 31278
rect 24032 31214 24084 31220
rect 24044 29050 24072 31214
rect 24136 29306 24164 33322
rect 24412 33046 24440 37606
rect 24596 37398 24624 38898
rect 24688 38418 24716 39442
rect 24780 38826 24808 41482
rect 24872 39914 24900 42720
rect 25780 42628 25832 42634
rect 25780 42570 25832 42576
rect 29736 42628 29788 42634
rect 29736 42570 29788 42576
rect 25596 42560 25648 42566
rect 25596 42502 25648 42508
rect 25412 42220 25464 42226
rect 25412 42162 25464 42168
rect 25044 41064 25096 41070
rect 25044 41006 25096 41012
rect 25056 40526 25084 41006
rect 25044 40520 25096 40526
rect 25044 40462 25096 40468
rect 24860 39908 24912 39914
rect 24860 39850 24912 39856
rect 24768 38820 24820 38826
rect 24768 38762 24820 38768
rect 24676 38412 24728 38418
rect 24676 38354 24728 38360
rect 24860 38344 24912 38350
rect 24780 38304 24860 38332
rect 24780 38298 24808 38304
rect 24688 38270 24808 38298
rect 24860 38286 24912 38292
rect 25320 38276 25372 38282
rect 24688 37466 24716 38270
rect 25320 38218 25372 38224
rect 24768 37936 24820 37942
rect 24768 37878 24820 37884
rect 24676 37460 24728 37466
rect 24676 37402 24728 37408
rect 24584 37392 24636 37398
rect 24584 37334 24636 37340
rect 24780 37194 24808 37878
rect 25332 37874 25360 38218
rect 25320 37868 25372 37874
rect 25320 37810 25372 37816
rect 24768 37188 24820 37194
rect 24768 37130 24820 37136
rect 24676 36576 24728 36582
rect 24676 36518 24728 36524
rect 24688 35698 24716 36518
rect 24780 36378 24808 37130
rect 25228 36780 25280 36786
rect 25228 36722 25280 36728
rect 24768 36372 24820 36378
rect 24768 36314 24820 36320
rect 24952 36236 25004 36242
rect 24952 36178 25004 36184
rect 24860 36168 24912 36174
rect 24860 36110 24912 36116
rect 24676 35692 24728 35698
rect 24676 35634 24728 35640
rect 24872 35018 24900 36110
rect 24964 35766 24992 36178
rect 25136 36100 25188 36106
rect 25136 36042 25188 36048
rect 24952 35760 25004 35766
rect 24952 35702 25004 35708
rect 25044 35760 25096 35766
rect 25044 35702 25096 35708
rect 24860 35012 24912 35018
rect 24860 34954 24912 34960
rect 24768 34400 24820 34406
rect 24768 34342 24820 34348
rect 24676 33924 24728 33930
rect 24676 33866 24728 33872
rect 24688 33658 24716 33866
rect 24676 33652 24728 33658
rect 24676 33594 24728 33600
rect 24780 33522 24808 34342
rect 24964 33998 24992 35702
rect 25056 35494 25084 35702
rect 25148 35494 25176 36042
rect 25044 35488 25096 35494
rect 25044 35430 25096 35436
rect 25136 35488 25188 35494
rect 25136 35430 25188 35436
rect 25148 35086 25176 35430
rect 25240 35290 25268 36722
rect 25228 35284 25280 35290
rect 25228 35226 25280 35232
rect 25136 35080 25188 35086
rect 25056 35040 25136 35068
rect 25056 34610 25084 35040
rect 25136 35022 25188 35028
rect 25228 35012 25280 35018
rect 25228 34954 25280 34960
rect 25240 34610 25268 34954
rect 25332 34950 25360 37810
rect 25320 34944 25372 34950
rect 25320 34886 25372 34892
rect 25044 34604 25096 34610
rect 25044 34546 25096 34552
rect 25228 34604 25280 34610
rect 25228 34546 25280 34552
rect 24952 33992 25004 33998
rect 24952 33934 25004 33940
rect 24768 33516 24820 33522
rect 24768 33458 24820 33464
rect 25136 33312 25188 33318
rect 25136 33254 25188 33260
rect 24400 33040 24452 33046
rect 24400 32982 24452 32988
rect 24952 32904 25004 32910
rect 24952 32846 25004 32852
rect 24676 32768 24728 32774
rect 24676 32710 24728 32716
rect 24688 32434 24716 32710
rect 24676 32428 24728 32434
rect 24676 32370 24728 32376
rect 24964 32026 24992 32846
rect 24952 32020 25004 32026
rect 24952 31962 25004 31968
rect 24492 31680 24544 31686
rect 24492 31622 24544 31628
rect 24400 29504 24452 29510
rect 24400 29446 24452 29452
rect 24124 29300 24176 29306
rect 24124 29242 24176 29248
rect 24136 29170 24348 29186
rect 24124 29164 24348 29170
rect 24176 29158 24348 29164
rect 24124 29106 24176 29112
rect 24216 29096 24268 29102
rect 24044 29044 24216 29050
rect 24044 29038 24268 29044
rect 24044 29022 24256 29038
rect 23952 28342 24072 28370
rect 23848 27532 23900 27538
rect 23848 27474 23900 27480
rect 23756 26784 23808 26790
rect 23756 26726 23808 26732
rect 23768 26518 23796 26726
rect 23756 26512 23808 26518
rect 23756 26454 23808 26460
rect 23756 25968 23808 25974
rect 23756 25910 23808 25916
rect 23768 25498 23796 25910
rect 23756 25492 23808 25498
rect 23756 25434 23808 25440
rect 23584 24942 23704 24970
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 23388 24744 23440 24750
rect 23388 24686 23440 24692
rect 23296 24268 23348 24274
rect 23296 24210 23348 24216
rect 22836 24200 22888 24206
rect 22836 24142 22888 24148
rect 23204 24200 23256 24206
rect 23204 24142 23256 24148
rect 23112 24064 23164 24070
rect 23112 24006 23164 24012
rect 22836 23656 22888 23662
rect 22836 23598 22888 23604
rect 22742 23366 22744 23418
rect 22796 23366 22798 23418
rect 22742 22330 22798 23366
rect 22742 22278 22744 22330
rect 22796 22278 22798 22330
rect 22742 21242 22798 22278
rect 22742 21190 22744 21242
rect 22796 21190 22798 21242
rect 22742 20154 22798 21190
rect 22742 20102 22744 20154
rect 22796 20102 22798 20154
rect 22742 19066 22798 20102
rect 22742 19014 22744 19066
rect 22796 19014 22798 19066
rect 22742 17978 22798 19014
rect 22742 17926 22744 17978
rect 22796 17926 22798 17978
rect 22742 16890 22798 17926
rect 22742 16838 22744 16890
rect 22796 16838 22798 16890
rect 22742 15802 22798 16838
rect 22742 15750 22744 15802
rect 22796 15750 22798 15802
rect 22742 14714 22798 15750
rect 22848 15366 22876 23598
rect 22928 22092 22980 22098
rect 22928 22034 22980 22040
rect 22940 21962 22968 22034
rect 22928 21956 22980 21962
rect 22928 21898 22980 21904
rect 22928 21344 22980 21350
rect 22928 21286 22980 21292
rect 22940 20466 22968 21286
rect 23124 21010 23152 24006
rect 23216 21690 23244 24142
rect 23400 23050 23428 24686
rect 23492 23322 23520 24754
rect 23480 23316 23532 23322
rect 23480 23258 23532 23264
rect 23388 23044 23440 23050
rect 23388 22986 23440 22992
rect 23388 22704 23440 22710
rect 23388 22646 23440 22652
rect 23400 22030 23428 22646
rect 23388 22024 23440 22030
rect 23388 21966 23440 21972
rect 23204 21684 23256 21690
rect 23204 21626 23256 21632
rect 23388 21480 23440 21486
rect 23388 21422 23440 21428
rect 23112 21004 23164 21010
rect 23164 20964 23244 20992
rect 23112 20946 23164 20952
rect 22928 20460 22980 20466
rect 22928 20402 22980 20408
rect 22940 17066 22968 20402
rect 23020 20324 23072 20330
rect 23020 20266 23072 20272
rect 23032 18970 23060 20266
rect 23020 18964 23072 18970
rect 23020 18906 23072 18912
rect 23020 18624 23072 18630
rect 23020 18566 23072 18572
rect 23032 17746 23060 18566
rect 23112 18284 23164 18290
rect 23112 18226 23164 18232
rect 23020 17740 23072 17746
rect 23020 17682 23072 17688
rect 23020 17536 23072 17542
rect 23020 17478 23072 17484
rect 22928 17060 22980 17066
rect 22928 17002 22980 17008
rect 22928 16788 22980 16794
rect 22928 16730 22980 16736
rect 22940 15570 22968 16730
rect 22928 15564 22980 15570
rect 22928 15506 22980 15512
rect 22836 15360 22888 15366
rect 22836 15302 22888 15308
rect 22928 14952 22980 14958
rect 22928 14894 22980 14900
rect 22742 14662 22744 14714
rect 22796 14662 22798 14714
rect 22742 13626 22798 14662
rect 22836 14476 22888 14482
rect 22836 14418 22888 14424
rect 22848 13802 22876 14418
rect 22940 14414 22968 14894
rect 22928 14408 22980 14414
rect 22928 14350 22980 14356
rect 22940 14074 22968 14350
rect 22928 14068 22980 14074
rect 22928 14010 22980 14016
rect 22928 13932 22980 13938
rect 22928 13874 22980 13880
rect 22836 13796 22888 13802
rect 22836 13738 22888 13744
rect 22742 13574 22744 13626
rect 22796 13574 22798 13626
rect 22742 12538 22798 13574
rect 22940 13258 22968 13874
rect 22928 13252 22980 13258
rect 22928 13194 22980 13200
rect 22742 12486 22744 12538
rect 22796 12486 22798 12538
rect 22742 11450 22798 12486
rect 23032 12434 23060 17478
rect 23124 17338 23152 18226
rect 23216 18170 23244 20964
rect 23400 20262 23428 21422
rect 23492 20602 23520 23258
rect 23480 20596 23532 20602
rect 23480 20538 23532 20544
rect 23388 20256 23440 20262
rect 23388 20198 23440 20204
rect 23400 20040 23428 20198
rect 23480 20052 23532 20058
rect 23400 20012 23480 20040
rect 23296 19508 23348 19514
rect 23296 19450 23348 19456
rect 23308 18766 23336 19450
rect 23400 19446 23428 20012
rect 23480 19994 23532 20000
rect 23480 19712 23532 19718
rect 23480 19654 23532 19660
rect 23388 19440 23440 19446
rect 23388 19382 23440 19388
rect 23388 19304 23440 19310
rect 23388 19246 23440 19252
rect 23296 18760 23348 18766
rect 23296 18702 23348 18708
rect 23400 18426 23428 19246
rect 23388 18420 23440 18426
rect 23388 18362 23440 18368
rect 23216 18142 23336 18170
rect 23204 18080 23256 18086
rect 23204 18022 23256 18028
rect 23216 17338 23244 18022
rect 23112 17332 23164 17338
rect 23112 17274 23164 17280
rect 23204 17332 23256 17338
rect 23204 17274 23256 17280
rect 23204 17060 23256 17066
rect 23204 17002 23256 17008
rect 23112 16584 23164 16590
rect 23112 16526 23164 16532
rect 23124 15910 23152 16526
rect 23216 16182 23244 17002
rect 23204 16176 23256 16182
rect 23204 16118 23256 16124
rect 23112 15904 23164 15910
rect 23112 15846 23164 15852
rect 23112 15564 23164 15570
rect 23112 15506 23164 15512
rect 22742 11398 22744 11450
rect 22796 11398 22798 11450
rect 22296 10526 22416 10554
rect 22100 9512 22152 9518
rect 22100 9454 22152 9460
rect 22296 9024 22324 10526
rect 22468 9920 22520 9926
rect 22468 9862 22520 9868
rect 22480 9586 22508 9862
rect 22468 9580 22520 9586
rect 22468 9522 22520 9528
rect 22468 9104 22520 9110
rect 22468 9046 22520 9052
rect 22296 8996 22416 9024
rect 22284 8900 22336 8906
rect 22284 8842 22336 8848
rect 22296 8294 22324 8842
rect 22284 8288 22336 8294
rect 22284 8230 22336 8236
rect 22008 7880 22060 7886
rect 22008 7822 22060 7828
rect 22100 7880 22152 7886
rect 22100 7822 22152 7828
rect 21824 7812 21876 7818
rect 21824 7754 21876 7760
rect 21836 7546 21864 7754
rect 21824 7540 21876 7546
rect 21824 7482 21876 7488
rect 21652 6854 21772 6882
rect 21548 3664 21600 3670
rect 21468 3612 21548 3618
rect 21468 3606 21600 3612
rect 21468 3590 21588 3606
rect 21272 2916 21324 2922
rect 21192 2876 21272 2904
rect 21272 2858 21324 2864
rect 20916 2746 21128 2774
rect 20720 1352 20772 1358
rect 20720 1294 20772 1300
rect 20916 1222 20944 2746
rect 21468 2310 21496 3590
rect 21652 2774 21680 6854
rect 22112 6798 22140 7822
rect 22192 7336 22244 7342
rect 22192 7278 22244 7284
rect 22100 6792 22152 6798
rect 22100 6734 22152 6740
rect 21824 6724 21876 6730
rect 21824 6666 21876 6672
rect 21732 6316 21784 6322
rect 21732 6258 21784 6264
rect 21744 4622 21772 6258
rect 21732 4616 21784 4622
rect 21732 4558 21784 4564
rect 21836 3942 21864 6666
rect 22204 6458 22232 7278
rect 22296 7002 22324 8230
rect 22388 8090 22416 8996
rect 22376 8084 22428 8090
rect 22376 8026 22428 8032
rect 22388 7342 22416 8026
rect 22376 7336 22428 7342
rect 22376 7278 22428 7284
rect 22284 6996 22336 7002
rect 22336 6956 22416 6984
rect 22284 6938 22336 6944
rect 22192 6452 22244 6458
rect 22192 6394 22244 6400
rect 22100 6112 22152 6118
rect 22100 6054 22152 6060
rect 22112 5710 22140 6054
rect 21916 5704 21968 5710
rect 22100 5704 22152 5710
rect 21968 5664 22048 5692
rect 21916 5646 21968 5652
rect 22020 5166 22048 5664
rect 22100 5646 22152 5652
rect 22388 5302 22416 6956
rect 22480 6322 22508 9046
rect 22572 8566 22600 10662
rect 22742 10362 22798 11398
rect 22742 10310 22744 10362
rect 22796 10310 22798 10362
rect 22652 9988 22704 9994
rect 22652 9930 22704 9936
rect 22664 9722 22692 9930
rect 22652 9716 22704 9722
rect 22652 9658 22704 9664
rect 22742 9274 22798 10310
rect 22742 9222 22744 9274
rect 22796 9222 22798 9274
rect 22652 8900 22704 8906
rect 22652 8842 22704 8848
rect 22560 8560 22612 8566
rect 22560 8502 22612 8508
rect 22560 8424 22612 8430
rect 22664 8412 22692 8842
rect 22612 8384 22692 8412
rect 22560 8366 22612 8372
rect 22742 8186 22798 9222
rect 22848 12406 23060 12434
rect 22848 8786 22876 12406
rect 23124 12306 23152 15506
rect 23308 14550 23336 18142
rect 23400 17660 23428 18362
rect 23492 17814 23520 19654
rect 23480 17808 23532 17814
rect 23480 17750 23532 17756
rect 23400 17632 23520 17660
rect 23388 16992 23440 16998
rect 23388 16934 23440 16940
rect 23400 16794 23428 16934
rect 23388 16788 23440 16794
rect 23388 16730 23440 16736
rect 23492 16674 23520 17632
rect 23400 16646 23520 16674
rect 23400 16130 23428 16646
rect 23480 16516 23532 16522
rect 23480 16458 23532 16464
rect 23492 16250 23520 16458
rect 23480 16244 23532 16250
rect 23480 16186 23532 16192
rect 23400 16102 23520 16130
rect 23584 16114 23612 24942
rect 23664 23724 23716 23730
rect 23664 23666 23716 23672
rect 23676 16250 23704 23666
rect 23940 22976 23992 22982
rect 23940 22918 23992 22924
rect 23756 22432 23808 22438
rect 23756 22374 23808 22380
rect 23768 22030 23796 22374
rect 23756 22024 23808 22030
rect 23756 21966 23808 21972
rect 23768 20466 23796 21966
rect 23756 20460 23808 20466
rect 23756 20402 23808 20408
rect 23848 19304 23900 19310
rect 23848 19246 23900 19252
rect 23860 18970 23888 19246
rect 23848 18964 23900 18970
rect 23848 18906 23900 18912
rect 23756 18828 23808 18834
rect 23756 18770 23808 18776
rect 23768 18290 23796 18770
rect 23848 18624 23900 18630
rect 23848 18566 23900 18572
rect 23756 18284 23808 18290
rect 23756 18226 23808 18232
rect 23768 17882 23796 18226
rect 23756 17876 23808 17882
rect 23756 17818 23808 17824
rect 23756 16992 23808 16998
rect 23756 16934 23808 16940
rect 23664 16244 23716 16250
rect 23664 16186 23716 16192
rect 23388 16040 23440 16046
rect 23388 15982 23440 15988
rect 23400 15434 23428 15982
rect 23492 15858 23520 16102
rect 23572 16108 23624 16114
rect 23572 16050 23624 16056
rect 23664 15904 23716 15910
rect 23492 15830 23612 15858
rect 23664 15846 23716 15852
rect 23388 15428 23440 15434
rect 23388 15370 23440 15376
rect 23388 15020 23440 15026
rect 23388 14962 23440 14968
rect 23400 14618 23428 14962
rect 23388 14612 23440 14618
rect 23388 14554 23440 14560
rect 23296 14544 23348 14550
rect 23296 14486 23348 14492
rect 23308 14278 23336 14486
rect 23388 14340 23440 14346
rect 23388 14282 23440 14288
rect 23296 14272 23348 14278
rect 23296 14214 23348 14220
rect 23400 13326 23428 14282
rect 23584 13530 23612 15830
rect 23676 15706 23704 15846
rect 23664 15700 23716 15706
rect 23664 15642 23716 15648
rect 23768 15502 23796 16934
rect 23756 15496 23808 15502
rect 23756 15438 23808 15444
rect 23664 15428 23716 15434
rect 23664 15370 23716 15376
rect 23676 15162 23704 15370
rect 23664 15156 23716 15162
rect 23664 15098 23716 15104
rect 23664 14408 23716 14414
rect 23768 14396 23796 15438
rect 23716 14368 23796 14396
rect 23664 14350 23716 14356
rect 23676 13852 23704 14350
rect 23756 13864 23808 13870
rect 23676 13824 23756 13852
rect 23572 13524 23624 13530
rect 23572 13466 23624 13472
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 23572 13184 23624 13190
rect 23572 13126 23624 13132
rect 23296 12844 23348 12850
rect 23296 12786 23348 12792
rect 23308 12442 23336 12786
rect 23296 12436 23348 12442
rect 23296 12378 23348 12384
rect 23480 12436 23532 12442
rect 23480 12378 23532 12384
rect 23492 12306 23520 12378
rect 23112 12300 23164 12306
rect 23112 12242 23164 12248
rect 23480 12300 23532 12306
rect 23480 12242 23532 12248
rect 23584 12238 23612 13126
rect 23676 12306 23704 13824
rect 23756 13806 23808 13812
rect 23860 12434 23888 18566
rect 23952 16114 23980 22918
rect 24044 21146 24072 28342
rect 24136 28098 24164 29022
rect 24216 28960 24268 28966
rect 24216 28902 24268 28908
rect 24228 28626 24256 28902
rect 24320 28694 24348 29158
rect 24308 28688 24360 28694
rect 24308 28630 24360 28636
rect 24216 28620 24268 28626
rect 24216 28562 24268 28568
rect 24412 28472 24440 29446
rect 24504 28506 24532 31622
rect 25148 31346 25176 33254
rect 25424 33114 25452 42162
rect 25608 42022 25636 42502
rect 25792 42226 25820 42570
rect 27894 42458 27950 42480
rect 27894 42406 27896 42458
rect 27948 42406 27950 42458
rect 25780 42220 25832 42226
rect 25780 42162 25832 42168
rect 27160 42220 27212 42226
rect 27160 42162 27212 42168
rect 26608 42152 26660 42158
rect 26608 42094 26660 42100
rect 25596 42016 25648 42022
rect 25596 41958 25648 41964
rect 26240 42016 26292 42022
rect 26240 41958 26292 41964
rect 25596 41676 25648 41682
rect 25596 41618 25648 41624
rect 25608 40662 25636 41618
rect 26056 41472 26108 41478
rect 26056 41414 26108 41420
rect 26068 41206 26096 41414
rect 26056 41200 26108 41206
rect 26056 41142 26108 41148
rect 25780 41132 25832 41138
rect 25780 41074 25832 41080
rect 25596 40656 25648 40662
rect 25596 40598 25648 40604
rect 25792 40526 25820 41074
rect 26056 40656 26108 40662
rect 26056 40598 26108 40604
rect 25780 40520 25832 40526
rect 25780 40462 25832 40468
rect 25596 39364 25648 39370
rect 25596 39306 25648 39312
rect 25608 39030 25636 39306
rect 25596 39024 25648 39030
rect 25596 38966 25648 38972
rect 25608 37126 25636 38966
rect 25792 38758 25820 40462
rect 25872 40384 25924 40390
rect 25872 40326 25924 40332
rect 25884 40032 25912 40326
rect 25964 40044 26016 40050
rect 25884 40004 25964 40032
rect 25884 39438 25912 40004
rect 25964 39986 26016 39992
rect 25964 39568 26016 39574
rect 25964 39510 26016 39516
rect 25872 39432 25924 39438
rect 25872 39374 25924 39380
rect 25884 38894 25912 39374
rect 25872 38888 25924 38894
rect 25872 38830 25924 38836
rect 25780 38752 25832 38758
rect 25780 38694 25832 38700
rect 25688 38208 25740 38214
rect 25688 38150 25740 38156
rect 25596 37120 25648 37126
rect 25596 37062 25648 37068
rect 25596 36644 25648 36650
rect 25596 36586 25648 36592
rect 25504 35080 25556 35086
rect 25504 35022 25556 35028
rect 25516 33590 25544 35022
rect 25504 33584 25556 33590
rect 25504 33526 25556 33532
rect 25412 33108 25464 33114
rect 25412 33050 25464 33056
rect 25504 31884 25556 31890
rect 25504 31826 25556 31832
rect 25136 31340 25188 31346
rect 25136 31282 25188 31288
rect 25136 31204 25188 31210
rect 25136 31146 25188 31152
rect 25228 31204 25280 31210
rect 25228 31146 25280 31152
rect 25044 31136 25096 31142
rect 25044 31078 25096 31084
rect 25056 30734 25084 31078
rect 25148 30734 25176 31146
rect 25044 30728 25096 30734
rect 25044 30670 25096 30676
rect 25136 30728 25188 30734
rect 25136 30670 25188 30676
rect 25240 30054 25268 31146
rect 25320 30592 25372 30598
rect 25320 30534 25372 30540
rect 25332 30190 25360 30534
rect 25320 30184 25372 30190
rect 25320 30126 25372 30132
rect 25228 30048 25280 30054
rect 25228 29990 25280 29996
rect 25332 29782 25360 30126
rect 25320 29776 25372 29782
rect 25320 29718 25372 29724
rect 24584 29708 24636 29714
rect 24584 29650 24636 29656
rect 24596 28966 24624 29650
rect 24676 29504 24728 29510
rect 24676 29446 24728 29452
rect 24688 29170 24716 29446
rect 24676 29164 24728 29170
rect 24676 29106 24728 29112
rect 24952 29096 25004 29102
rect 24952 29038 25004 29044
rect 25136 29096 25188 29102
rect 25136 29038 25188 29044
rect 24676 29028 24728 29034
rect 24676 28970 24728 28976
rect 24584 28960 24636 28966
rect 24584 28902 24636 28908
rect 24504 28478 24624 28506
rect 24228 28444 24440 28472
rect 24228 28218 24256 28444
rect 24492 28416 24544 28422
rect 24492 28358 24544 28364
rect 24216 28212 24268 28218
rect 24216 28154 24268 28160
rect 24308 28212 24360 28218
rect 24308 28154 24360 28160
rect 24136 28070 24256 28098
rect 24124 28008 24176 28014
rect 24124 27950 24176 27956
rect 24136 27470 24164 27950
rect 24124 27464 24176 27470
rect 24124 27406 24176 27412
rect 24124 26920 24176 26926
rect 24124 26862 24176 26868
rect 24136 26450 24164 26862
rect 24124 26444 24176 26450
rect 24124 26386 24176 26392
rect 24228 26058 24256 28070
rect 24320 27606 24348 28154
rect 24400 28144 24452 28150
rect 24400 28086 24452 28092
rect 24308 27600 24360 27606
rect 24308 27542 24360 27548
rect 24412 27470 24440 28086
rect 24504 27674 24532 28358
rect 24596 28218 24624 28478
rect 24584 28212 24636 28218
rect 24584 28154 24636 28160
rect 24688 28082 24716 28970
rect 24768 28620 24820 28626
rect 24768 28562 24820 28568
rect 24780 28422 24808 28562
rect 24768 28416 24820 28422
rect 24768 28358 24820 28364
rect 24860 28416 24912 28422
rect 24860 28358 24912 28364
rect 24768 28212 24820 28218
rect 24768 28154 24820 28160
rect 24584 28076 24636 28082
rect 24584 28018 24636 28024
rect 24676 28076 24728 28082
rect 24676 28018 24728 28024
rect 24596 27962 24624 28018
rect 24596 27934 24716 27962
rect 24688 27878 24716 27934
rect 24584 27872 24636 27878
rect 24584 27814 24636 27820
rect 24676 27872 24728 27878
rect 24676 27814 24728 27820
rect 24492 27668 24544 27674
rect 24492 27610 24544 27616
rect 24400 27464 24452 27470
rect 24400 27406 24452 27412
rect 24492 26376 24544 26382
rect 24492 26318 24544 26324
rect 24228 26030 24440 26058
rect 24504 26042 24532 26318
rect 24124 25220 24176 25226
rect 24124 25162 24176 25168
rect 24136 23594 24164 25162
rect 24308 25152 24360 25158
rect 24308 25094 24360 25100
rect 24216 24200 24268 24206
rect 24216 24142 24268 24148
rect 24124 23588 24176 23594
rect 24124 23530 24176 23536
rect 24124 23180 24176 23186
rect 24124 23122 24176 23128
rect 24032 21140 24084 21146
rect 24032 21082 24084 21088
rect 24032 18760 24084 18766
rect 24032 18702 24084 18708
rect 24044 18154 24072 18702
rect 24136 18630 24164 23122
rect 24228 22642 24256 24142
rect 24320 23050 24348 25094
rect 24308 23044 24360 23050
rect 24308 22986 24360 22992
rect 24308 22772 24360 22778
rect 24308 22714 24360 22720
rect 24216 22636 24268 22642
rect 24216 22578 24268 22584
rect 24216 20392 24268 20398
rect 24216 20334 24268 20340
rect 24124 18624 24176 18630
rect 24124 18566 24176 18572
rect 24228 18426 24256 20334
rect 24320 20262 24348 22714
rect 24308 20256 24360 20262
rect 24308 20198 24360 20204
rect 24308 19372 24360 19378
rect 24308 19314 24360 19320
rect 24216 18420 24268 18426
rect 24216 18362 24268 18368
rect 24124 18352 24176 18358
rect 24124 18294 24176 18300
rect 24032 18148 24084 18154
rect 24032 18090 24084 18096
rect 24136 17882 24164 18294
rect 24124 17876 24176 17882
rect 24124 17818 24176 17824
rect 24032 17808 24084 17814
rect 24032 17750 24084 17756
rect 24044 16794 24072 17750
rect 24216 17536 24268 17542
rect 24216 17478 24268 17484
rect 24228 17202 24256 17478
rect 24320 17338 24348 19314
rect 24308 17332 24360 17338
rect 24308 17274 24360 17280
rect 24216 17196 24268 17202
rect 24216 17138 24268 17144
rect 24412 16946 24440 26030
rect 24492 26036 24544 26042
rect 24492 25978 24544 25984
rect 24504 25498 24532 25978
rect 24492 25492 24544 25498
rect 24492 25434 24544 25440
rect 24596 22778 24624 27814
rect 24780 27334 24808 28154
rect 24872 27878 24900 28358
rect 24964 27946 24992 29038
rect 25044 28552 25096 28558
rect 25044 28494 25096 28500
rect 25056 28218 25084 28494
rect 25044 28212 25096 28218
rect 25044 28154 25096 28160
rect 24952 27940 25004 27946
rect 24952 27882 25004 27888
rect 24860 27872 24912 27878
rect 24860 27814 24912 27820
rect 25148 27402 25176 29038
rect 25516 28762 25544 31826
rect 25504 28756 25556 28762
rect 25504 28698 25556 28704
rect 25320 28688 25372 28694
rect 25320 28630 25372 28636
rect 25228 28484 25280 28490
rect 25228 28426 25280 28432
rect 25240 28218 25268 28426
rect 25228 28212 25280 28218
rect 25228 28154 25280 28160
rect 25136 27396 25188 27402
rect 25136 27338 25188 27344
rect 24768 27328 24820 27334
rect 24768 27270 24820 27276
rect 25044 27124 25096 27130
rect 25044 27066 25096 27072
rect 24768 26784 24820 26790
rect 24768 26726 24820 26732
rect 24780 25362 24808 26726
rect 25056 26382 25084 27066
rect 25044 26376 25096 26382
rect 25044 26318 25096 26324
rect 24768 25356 24820 25362
rect 24768 25298 24820 25304
rect 24676 24880 24728 24886
rect 24676 24822 24728 24828
rect 24688 24138 24716 24822
rect 24780 24614 24808 25298
rect 24952 25220 25004 25226
rect 25056 25208 25084 26318
rect 25004 25180 25084 25208
rect 24952 25162 25004 25168
rect 24768 24608 24820 24614
rect 24768 24550 24820 24556
rect 24676 24132 24728 24138
rect 24676 24074 24728 24080
rect 25148 23594 25176 27338
rect 25228 26784 25280 26790
rect 25228 26726 25280 26732
rect 25240 26246 25268 26726
rect 25228 26240 25280 26246
rect 25228 26182 25280 26188
rect 25240 25294 25268 26182
rect 25228 25288 25280 25294
rect 25228 25230 25280 25236
rect 25240 24818 25268 25230
rect 25332 25158 25360 28630
rect 25412 28552 25464 28558
rect 25412 28494 25464 28500
rect 25320 25152 25372 25158
rect 25320 25094 25372 25100
rect 25228 24812 25280 24818
rect 25228 24754 25280 24760
rect 25240 23730 25268 24754
rect 25228 23724 25280 23730
rect 25228 23666 25280 23672
rect 25136 23588 25188 23594
rect 25136 23530 25188 23536
rect 24768 23520 24820 23526
rect 24768 23462 24820 23468
rect 24676 23316 24728 23322
rect 24676 23258 24728 23264
rect 24584 22772 24636 22778
rect 24584 22714 24636 22720
rect 24688 22710 24716 23258
rect 24676 22704 24728 22710
rect 24676 22646 24728 22652
rect 24492 22636 24544 22642
rect 24492 22578 24544 22584
rect 24504 21690 24532 22578
rect 24584 22024 24636 22030
rect 24584 21966 24636 21972
rect 24492 21684 24544 21690
rect 24492 21626 24544 21632
rect 24596 20602 24624 21966
rect 24584 20596 24636 20602
rect 24584 20538 24636 20544
rect 24688 20346 24716 22646
rect 24780 21554 24808 23462
rect 24952 23316 25004 23322
rect 24952 23258 25004 23264
rect 24860 22024 24912 22030
rect 24860 21966 24912 21972
rect 24872 21622 24900 21966
rect 24964 21894 24992 23258
rect 25136 23112 25188 23118
rect 25136 23054 25188 23060
rect 25044 22976 25096 22982
rect 25044 22918 25096 22924
rect 24952 21888 25004 21894
rect 24952 21830 25004 21836
rect 24860 21616 24912 21622
rect 24860 21558 24912 21564
rect 24768 21548 24820 21554
rect 24768 21490 24820 21496
rect 24768 21412 24820 21418
rect 24768 21354 24820 21360
rect 24780 20942 24808 21354
rect 24964 20942 24992 21830
rect 25056 21350 25084 22918
rect 25044 21344 25096 21350
rect 25044 21286 25096 21292
rect 24768 20936 24820 20942
rect 24952 20936 25004 20942
rect 24820 20896 24900 20924
rect 24768 20878 24820 20884
rect 24872 20466 24900 20896
rect 24952 20878 25004 20884
rect 24768 20460 24820 20466
rect 24768 20402 24820 20408
rect 24860 20460 24912 20466
rect 24860 20402 24912 20408
rect 24504 20318 24716 20346
rect 24504 18970 24532 20318
rect 24676 20256 24728 20262
rect 24676 20198 24728 20204
rect 24688 19938 24716 20198
rect 24780 20058 24808 20402
rect 24860 20324 24912 20330
rect 24860 20266 24912 20272
rect 24768 20052 24820 20058
rect 24768 19994 24820 20000
rect 24688 19910 24808 19938
rect 24872 19922 24900 20266
rect 24676 19780 24728 19786
rect 24676 19722 24728 19728
rect 24492 18964 24544 18970
rect 24492 18906 24544 18912
rect 24584 18760 24636 18766
rect 24584 18702 24636 18708
rect 24492 18624 24544 18630
rect 24492 18566 24544 18572
rect 24504 18358 24532 18566
rect 24492 18352 24544 18358
rect 24492 18294 24544 18300
rect 24492 18148 24544 18154
rect 24492 18090 24544 18096
rect 24504 17202 24532 18090
rect 24596 17678 24624 18702
rect 24688 18698 24716 19722
rect 24676 18692 24728 18698
rect 24676 18634 24728 18640
rect 24584 17672 24636 17678
rect 24584 17614 24636 17620
rect 24492 17196 24544 17202
rect 24492 17138 24544 17144
rect 24136 16918 24440 16946
rect 24492 16992 24544 16998
rect 24492 16934 24544 16940
rect 24032 16788 24084 16794
rect 24032 16730 24084 16736
rect 24032 16448 24084 16454
rect 24032 16390 24084 16396
rect 23940 16108 23992 16114
rect 23940 16050 23992 16056
rect 23940 15700 23992 15706
rect 23940 15642 23992 15648
rect 23952 15094 23980 15642
rect 24044 15162 24072 16390
rect 24032 15156 24084 15162
rect 24032 15098 24084 15104
rect 23940 15088 23992 15094
rect 23940 15030 23992 15036
rect 24032 14272 24084 14278
rect 24032 14214 24084 14220
rect 23940 13320 23992 13326
rect 23940 13262 23992 13268
rect 23952 12646 23980 13262
rect 23940 12640 23992 12646
rect 23940 12582 23992 12588
rect 23768 12406 23888 12434
rect 23664 12300 23716 12306
rect 23664 12242 23716 12248
rect 23572 12232 23624 12238
rect 23572 12174 23624 12180
rect 23676 12170 23704 12242
rect 23664 12164 23716 12170
rect 23664 12106 23716 12112
rect 23388 12096 23440 12102
rect 23388 12038 23440 12044
rect 23572 12096 23624 12102
rect 23572 12038 23624 12044
rect 23020 11620 23072 11626
rect 23020 11562 23072 11568
rect 23204 11620 23256 11626
rect 23204 11562 23256 11568
rect 22928 11076 22980 11082
rect 22928 11018 22980 11024
rect 22940 9450 22968 11018
rect 23032 9738 23060 11562
rect 23216 11150 23244 11562
rect 23296 11552 23348 11558
rect 23296 11494 23348 11500
rect 23204 11144 23256 11150
rect 23124 11104 23204 11132
rect 23124 10606 23152 11104
rect 23204 11086 23256 11092
rect 23204 11008 23256 11014
rect 23204 10950 23256 10956
rect 23216 10674 23244 10950
rect 23204 10668 23256 10674
rect 23204 10610 23256 10616
rect 23308 10606 23336 11494
rect 23400 11082 23428 12038
rect 23584 11762 23612 12038
rect 23664 11892 23716 11898
rect 23664 11834 23716 11840
rect 23572 11756 23624 11762
rect 23572 11698 23624 11704
rect 23480 11280 23532 11286
rect 23480 11222 23532 11228
rect 23388 11076 23440 11082
rect 23388 11018 23440 11024
rect 23492 10690 23520 11222
rect 23400 10662 23520 10690
rect 23112 10600 23164 10606
rect 23112 10542 23164 10548
rect 23296 10600 23348 10606
rect 23296 10542 23348 10548
rect 23124 9926 23152 10542
rect 23308 9994 23336 10542
rect 23296 9988 23348 9994
rect 23296 9930 23348 9936
rect 23112 9920 23164 9926
rect 23112 9862 23164 9868
rect 23032 9710 23244 9738
rect 23020 9648 23072 9654
rect 23020 9590 23072 9596
rect 22928 9444 22980 9450
rect 22928 9386 22980 9392
rect 23032 8838 23060 9590
rect 23216 9382 23244 9710
rect 23308 9586 23336 9930
rect 23296 9580 23348 9586
rect 23296 9522 23348 9528
rect 23204 9376 23256 9382
rect 23204 9318 23256 9324
rect 23296 9376 23348 9382
rect 23296 9318 23348 9324
rect 23216 9110 23244 9318
rect 23204 9104 23256 9110
rect 23204 9046 23256 9052
rect 23204 8968 23256 8974
rect 23204 8910 23256 8916
rect 23020 8832 23072 8838
rect 22848 8758 22968 8786
rect 23020 8774 23072 8780
rect 22836 8424 22888 8430
rect 22836 8366 22888 8372
rect 22742 8134 22744 8186
rect 22796 8134 22798 8186
rect 22652 7404 22704 7410
rect 22652 7346 22704 7352
rect 22664 7002 22692 7346
rect 22742 7098 22798 8134
rect 22848 7546 22876 8366
rect 22836 7540 22888 7546
rect 22836 7482 22888 7488
rect 22742 7046 22744 7098
rect 22796 7046 22798 7098
rect 22652 6996 22704 7002
rect 22652 6938 22704 6944
rect 22468 6316 22520 6322
rect 22468 6258 22520 6264
rect 22652 6112 22704 6118
rect 22652 6054 22704 6060
rect 22560 5636 22612 5642
rect 22560 5578 22612 5584
rect 22376 5296 22428 5302
rect 22376 5238 22428 5244
rect 22008 5160 22060 5166
rect 22060 5120 22140 5148
rect 22008 5102 22060 5108
rect 22008 5024 22060 5030
rect 22008 4966 22060 4972
rect 22020 4146 22048 4966
rect 22112 4758 22140 5120
rect 22192 5024 22244 5030
rect 22192 4966 22244 4972
rect 22100 4752 22152 4758
rect 22100 4694 22152 4700
rect 22112 4214 22140 4694
rect 22100 4208 22152 4214
rect 22100 4150 22152 4156
rect 22008 4140 22060 4146
rect 22008 4082 22060 4088
rect 21824 3936 21876 3942
rect 21824 3878 21876 3884
rect 22204 3534 22232 4966
rect 22572 4622 22600 5578
rect 22560 4616 22612 4622
rect 22560 4558 22612 4564
rect 22572 4146 22600 4558
rect 22560 4140 22612 4146
rect 22560 4082 22612 4088
rect 22664 4078 22692 6054
rect 22742 6010 22798 7046
rect 22940 6866 22968 8758
rect 23216 8650 23244 8910
rect 23124 8622 23244 8650
rect 23020 8560 23072 8566
rect 23020 8502 23072 8508
rect 22928 6860 22980 6866
rect 22928 6802 22980 6808
rect 22836 6656 22888 6662
rect 22836 6598 22888 6604
rect 22848 6254 22876 6598
rect 22836 6248 22888 6254
rect 22836 6190 22888 6196
rect 22742 5958 22744 6010
rect 22796 5958 22798 6010
rect 22742 4922 22798 5958
rect 22742 4870 22744 4922
rect 22796 4870 22798 4922
rect 22652 4072 22704 4078
rect 22652 4014 22704 4020
rect 22742 3834 22798 4870
rect 22742 3782 22744 3834
rect 22796 3782 22798 3834
rect 22192 3528 22244 3534
rect 22192 3470 22244 3476
rect 22284 3528 22336 3534
rect 22284 3470 22336 3476
rect 22560 3528 22612 3534
rect 22560 3470 22612 3476
rect 22296 3058 22324 3470
rect 22572 3058 22600 3470
rect 22284 3052 22336 3058
rect 22284 2994 22336 3000
rect 22560 3052 22612 3058
rect 22560 2994 22612 3000
rect 22652 2848 22704 2854
rect 22652 2790 22704 2796
rect 21560 2746 21680 2774
rect 21456 2304 21508 2310
rect 21456 2246 21508 2252
rect 21560 1426 21588 2746
rect 21916 2440 21968 2446
rect 21916 2382 21968 2388
rect 21928 1970 21956 2382
rect 21916 1964 21968 1970
rect 21916 1906 21968 1912
rect 22468 1964 22520 1970
rect 22468 1906 22520 1912
rect 22480 1562 22508 1906
rect 22468 1556 22520 1562
rect 22468 1498 22520 1504
rect 21548 1420 21600 1426
rect 21548 1362 21600 1368
rect 22664 1358 22692 2790
rect 22742 2746 22798 3782
rect 22848 3534 22876 6190
rect 22836 3528 22888 3534
rect 22836 3470 22888 3476
rect 22742 2694 22744 2746
rect 22796 2694 22798 2746
rect 22742 1658 22798 2694
rect 22848 2650 22876 3470
rect 23032 3058 23060 8502
rect 23124 8498 23152 8622
rect 23112 8492 23164 8498
rect 23112 8434 23164 8440
rect 23204 8492 23256 8498
rect 23204 8434 23256 8440
rect 23216 7002 23244 8434
rect 23308 8294 23336 9318
rect 23296 8288 23348 8294
rect 23296 8230 23348 8236
rect 23400 7478 23428 10662
rect 23676 10062 23704 11834
rect 23768 10674 23796 12406
rect 24044 12170 24072 14214
rect 24136 12374 24164 16918
rect 24216 16788 24268 16794
rect 24216 16730 24268 16736
rect 24400 16788 24452 16794
rect 24400 16730 24452 16736
rect 24228 13818 24256 16730
rect 24308 16584 24360 16590
rect 24308 16526 24360 16532
rect 24320 16096 24348 16526
rect 24412 16250 24440 16730
rect 24504 16590 24532 16934
rect 24596 16590 24624 17614
rect 24676 17264 24728 17270
rect 24676 17206 24728 17212
rect 24688 16794 24716 17206
rect 24780 16998 24808 19910
rect 24860 19916 24912 19922
rect 24860 19858 24912 19864
rect 24964 19378 24992 20878
rect 25148 20874 25176 23054
rect 25320 21480 25372 21486
rect 25320 21422 25372 21428
rect 25136 20868 25188 20874
rect 25136 20810 25188 20816
rect 25148 20346 25176 20810
rect 25148 20318 25268 20346
rect 25136 20256 25188 20262
rect 25136 20198 25188 20204
rect 25148 19786 25176 20198
rect 25240 19990 25268 20318
rect 25228 19984 25280 19990
rect 25228 19926 25280 19932
rect 25136 19780 25188 19786
rect 25136 19722 25188 19728
rect 25044 19508 25096 19514
rect 25044 19450 25096 19456
rect 24952 19372 25004 19378
rect 24952 19314 25004 19320
rect 25056 17678 25084 19450
rect 25148 18358 25176 19722
rect 25136 18352 25188 18358
rect 25136 18294 25188 18300
rect 25240 18204 25268 19926
rect 25148 18176 25268 18204
rect 25044 17672 25096 17678
rect 25044 17614 25096 17620
rect 24952 17536 25004 17542
rect 24952 17478 25004 17484
rect 24860 17196 24912 17202
rect 24860 17138 24912 17144
rect 24768 16992 24820 16998
rect 24768 16934 24820 16940
rect 24676 16788 24728 16794
rect 24676 16730 24728 16736
rect 24492 16584 24544 16590
rect 24492 16526 24544 16532
rect 24584 16584 24636 16590
rect 24636 16544 24716 16572
rect 24584 16526 24636 16532
rect 24400 16244 24452 16250
rect 24400 16186 24452 16192
rect 24688 16130 24716 16544
rect 24400 16108 24452 16114
rect 24320 16068 24400 16096
rect 24628 16102 24716 16130
rect 24628 16096 24656 16102
rect 24400 16050 24452 16056
rect 24504 16068 24656 16096
rect 24400 15972 24452 15978
rect 24320 15932 24400 15960
rect 24320 15502 24348 15932
rect 24400 15914 24452 15920
rect 24308 15496 24360 15502
rect 24308 15438 24360 15444
rect 24320 14414 24348 15438
rect 24504 14958 24532 16068
rect 24676 16040 24728 16046
rect 24728 16000 24808 16028
rect 24676 15982 24728 15988
rect 24584 15972 24636 15978
rect 24584 15914 24636 15920
rect 24596 15722 24624 15914
rect 24596 15694 24716 15722
rect 24688 15586 24716 15694
rect 24780 15638 24808 16000
rect 24628 15558 24716 15586
rect 24768 15632 24820 15638
rect 24768 15574 24820 15580
rect 24628 15484 24656 15558
rect 24596 15456 24656 15484
rect 24768 15496 24820 15502
rect 24492 14952 24544 14958
rect 24492 14894 24544 14900
rect 24308 14408 24360 14414
rect 24308 14350 24360 14356
rect 24504 14346 24532 14894
rect 24492 14340 24544 14346
rect 24492 14282 24544 14288
rect 24228 13790 24440 13818
rect 24216 13728 24268 13734
rect 24216 13670 24268 13676
rect 24228 13326 24256 13670
rect 24308 13524 24360 13530
rect 24308 13466 24360 13472
rect 24216 13320 24268 13326
rect 24216 13262 24268 13268
rect 24124 12368 24176 12374
rect 24124 12310 24176 12316
rect 24032 12164 24084 12170
rect 24032 12106 24084 12112
rect 23940 11756 23992 11762
rect 23940 11698 23992 11704
rect 23952 10810 23980 11698
rect 23940 10804 23992 10810
rect 23940 10746 23992 10752
rect 24032 10736 24084 10742
rect 24032 10678 24084 10684
rect 23756 10668 23808 10674
rect 23756 10610 23808 10616
rect 23848 10668 23900 10674
rect 23848 10610 23900 10616
rect 23664 10056 23716 10062
rect 23664 9998 23716 10004
rect 23572 9444 23624 9450
rect 23572 9386 23624 9392
rect 23388 7472 23440 7478
rect 23388 7414 23440 7420
rect 23296 7336 23348 7342
rect 23296 7278 23348 7284
rect 23204 6996 23256 7002
rect 23204 6938 23256 6944
rect 23216 5574 23244 6938
rect 23308 6798 23336 7278
rect 23296 6792 23348 6798
rect 23296 6734 23348 6740
rect 23204 5568 23256 5574
rect 23204 5510 23256 5516
rect 23112 4752 23164 4758
rect 23112 4694 23164 4700
rect 23124 3058 23152 4694
rect 23216 4690 23244 5510
rect 23308 5098 23336 6734
rect 23480 6112 23532 6118
rect 23480 6054 23532 6060
rect 23492 5302 23520 6054
rect 23480 5296 23532 5302
rect 23480 5238 23532 5244
rect 23296 5092 23348 5098
rect 23296 5034 23348 5040
rect 23584 4690 23612 9386
rect 23768 9382 23796 10610
rect 23860 10266 23888 10610
rect 24044 10266 24072 10678
rect 23848 10260 23900 10266
rect 23848 10202 23900 10208
rect 24032 10260 24084 10266
rect 24032 10202 24084 10208
rect 24136 9654 24164 12310
rect 24320 12102 24348 13466
rect 24308 12096 24360 12102
rect 24308 12038 24360 12044
rect 24216 10464 24268 10470
rect 24216 10406 24268 10412
rect 24228 9994 24256 10406
rect 24216 9988 24268 9994
rect 24216 9930 24268 9936
rect 24124 9648 24176 9654
rect 24124 9590 24176 9596
rect 23756 9376 23808 9382
rect 23756 9318 23808 9324
rect 24124 9376 24176 9382
rect 24124 9318 24176 9324
rect 23756 8832 23808 8838
rect 23756 8774 23808 8780
rect 23768 8362 23796 8774
rect 23756 8356 23808 8362
rect 23756 8298 23808 8304
rect 23664 7744 23716 7750
rect 23664 7686 23716 7692
rect 23676 7410 23704 7686
rect 23768 7410 23796 8298
rect 24136 7886 24164 9318
rect 24124 7880 24176 7886
rect 24124 7822 24176 7828
rect 23664 7404 23716 7410
rect 23664 7346 23716 7352
rect 23756 7404 23808 7410
rect 23756 7346 23808 7352
rect 23756 6112 23808 6118
rect 23756 6054 23808 6060
rect 23664 5636 23716 5642
rect 23664 5578 23716 5584
rect 23204 4684 23256 4690
rect 23204 4626 23256 4632
rect 23572 4684 23624 4690
rect 23572 4626 23624 4632
rect 23204 4072 23256 4078
rect 23204 4014 23256 4020
rect 23020 3052 23072 3058
rect 23020 2994 23072 3000
rect 23112 3052 23164 3058
rect 23112 2994 23164 3000
rect 23032 2922 23060 2994
rect 23020 2916 23072 2922
rect 23020 2858 23072 2864
rect 22836 2644 22888 2650
rect 22836 2586 22888 2592
rect 22928 2372 22980 2378
rect 22928 2314 22980 2320
rect 22742 1606 22744 1658
rect 22796 1606 22798 1658
rect 22008 1352 22060 1358
rect 22008 1294 22060 1300
rect 22652 1352 22704 1358
rect 22652 1294 22704 1300
rect 19708 1216 19760 1222
rect 19708 1158 19760 1164
rect 20904 1216 20956 1222
rect 20904 1158 20956 1164
rect 22020 950 22048 1294
rect 22742 1040 22798 1606
rect 22940 1358 22968 2314
rect 23032 2106 23060 2858
rect 23124 2446 23152 2994
rect 23112 2440 23164 2446
rect 23112 2382 23164 2388
rect 23020 2100 23072 2106
rect 23020 2042 23072 2048
rect 23216 1426 23244 4014
rect 23572 3936 23624 3942
rect 23572 3878 23624 3884
rect 23584 3534 23612 3878
rect 23676 3738 23704 5578
rect 23768 3738 23796 6054
rect 24032 5704 24084 5710
rect 24032 5646 24084 5652
rect 24044 5234 24072 5646
rect 24032 5228 24084 5234
rect 24032 5170 24084 5176
rect 23848 4684 23900 4690
rect 23848 4626 23900 4632
rect 23860 4146 23888 4626
rect 23848 4140 23900 4146
rect 23848 4082 23900 4088
rect 23664 3732 23716 3738
rect 23664 3674 23716 3680
rect 23756 3732 23808 3738
rect 23756 3674 23808 3680
rect 23572 3528 23624 3534
rect 23572 3470 23624 3476
rect 23296 3052 23348 3058
rect 23296 2994 23348 3000
rect 23204 1420 23256 1426
rect 23204 1362 23256 1368
rect 22928 1352 22980 1358
rect 22928 1294 22980 1300
rect 23308 1222 23336 2994
rect 24044 2446 24072 5170
rect 24124 4072 24176 4078
rect 24124 4014 24176 4020
rect 24136 3602 24164 4014
rect 24124 3596 24176 3602
rect 24124 3538 24176 3544
rect 24032 2440 24084 2446
rect 24032 2382 24084 2388
rect 23572 2304 23624 2310
rect 23572 2246 23624 2252
rect 23584 1358 23612 2246
rect 24044 1970 24072 2382
rect 24032 1964 24084 1970
rect 24032 1906 24084 1912
rect 23572 1352 23624 1358
rect 23572 1294 23624 1300
rect 23296 1216 23348 1222
rect 23296 1158 23348 1164
rect 22008 944 22060 950
rect 22008 886 22060 892
rect 19616 876 19668 882
rect 19616 818 19668 824
rect 24320 814 24348 12038
rect 24412 11014 24440 13790
rect 24492 12912 24544 12918
rect 24492 12854 24544 12860
rect 24504 11778 24532 12854
rect 24596 12832 24624 15456
rect 24768 15438 24820 15444
rect 24780 15144 24808 15438
rect 24872 15434 24900 17138
rect 24964 17134 24992 17478
rect 24952 17128 25004 17134
rect 24952 17070 25004 17076
rect 24860 15428 24912 15434
rect 24860 15370 24912 15376
rect 24688 15116 24900 15144
rect 24688 14074 24716 15116
rect 24768 15020 24820 15026
rect 24768 14962 24820 14968
rect 24676 14068 24728 14074
rect 24676 14010 24728 14016
rect 24676 13864 24728 13870
rect 24676 13806 24728 13812
rect 24688 13258 24716 13806
rect 24780 13394 24808 14962
rect 24872 14278 24900 15116
rect 24964 15094 24992 17070
rect 25044 16652 25096 16658
rect 25044 16594 25096 16600
rect 24952 15088 25004 15094
rect 24952 15030 25004 15036
rect 25056 14906 25084 16594
rect 24964 14878 25084 14906
rect 24964 14550 24992 14878
rect 25044 14816 25096 14822
rect 25044 14758 25096 14764
rect 25056 14550 25084 14758
rect 24952 14544 25004 14550
rect 24952 14486 25004 14492
rect 25044 14544 25096 14550
rect 25044 14486 25096 14492
rect 24860 14272 24912 14278
rect 24860 14214 24912 14220
rect 24860 14068 24912 14074
rect 24860 14010 24912 14016
rect 24768 13388 24820 13394
rect 24768 13330 24820 13336
rect 24676 13252 24728 13258
rect 24676 13194 24728 13200
rect 24596 12804 24716 12832
rect 24584 11824 24636 11830
rect 24504 11772 24584 11778
rect 24504 11766 24636 11772
rect 24504 11750 24624 11766
rect 24400 11008 24452 11014
rect 24400 10950 24452 10956
rect 24412 8498 24440 10950
rect 24400 8492 24452 8498
rect 24400 8434 24452 8440
rect 24504 8294 24532 11750
rect 24584 8356 24636 8362
rect 24584 8298 24636 8304
rect 24492 8288 24544 8294
rect 24492 8230 24544 8236
rect 24492 7336 24544 7342
rect 24492 7278 24544 7284
rect 24504 7002 24532 7278
rect 24492 6996 24544 7002
rect 24492 6938 24544 6944
rect 24596 6798 24624 8298
rect 24584 6792 24636 6798
rect 24584 6734 24636 6740
rect 24492 6316 24544 6322
rect 24492 6258 24544 6264
rect 24504 5914 24532 6258
rect 24584 6180 24636 6186
rect 24584 6122 24636 6128
rect 24492 5908 24544 5914
rect 24492 5850 24544 5856
rect 24492 3052 24544 3058
rect 24492 2994 24544 3000
rect 24504 2582 24532 2994
rect 24596 2922 24624 6122
rect 24584 2916 24636 2922
rect 24584 2858 24636 2864
rect 24492 2576 24544 2582
rect 24492 2518 24544 2524
rect 24596 2378 24624 2858
rect 24688 2774 24716 12804
rect 24768 12096 24820 12102
rect 24768 12038 24820 12044
rect 24780 11898 24808 12038
rect 24768 11892 24820 11898
rect 24768 11834 24820 11840
rect 24872 9654 24900 14010
rect 25056 12850 25084 14486
rect 25148 14074 25176 18176
rect 25228 16992 25280 16998
rect 25228 16934 25280 16940
rect 25240 16590 25268 16934
rect 25228 16584 25280 16590
rect 25228 16526 25280 16532
rect 25228 16176 25280 16182
rect 25228 16118 25280 16124
rect 25240 15026 25268 16118
rect 25228 15020 25280 15026
rect 25228 14962 25280 14968
rect 25228 14884 25280 14890
rect 25228 14826 25280 14832
rect 25136 14068 25188 14074
rect 25136 14010 25188 14016
rect 25240 13938 25268 14826
rect 25228 13932 25280 13938
rect 25228 13874 25280 13880
rect 25044 12844 25096 12850
rect 25044 12786 25096 12792
rect 24952 12776 25004 12782
rect 24952 12718 25004 12724
rect 24964 12238 24992 12718
rect 25056 12238 25084 12786
rect 25228 12640 25280 12646
rect 25228 12582 25280 12588
rect 24952 12232 25004 12238
rect 24952 12174 25004 12180
rect 25044 12232 25096 12238
rect 25044 12174 25096 12180
rect 25240 11558 25268 12582
rect 25228 11552 25280 11558
rect 25228 11494 25280 11500
rect 24952 10532 25004 10538
rect 24952 10474 25004 10480
rect 24860 9648 24912 9654
rect 24860 9590 24912 9596
rect 24872 8906 24900 9590
rect 24964 9330 24992 10474
rect 25044 9580 25096 9586
rect 25096 9540 25268 9568
rect 25044 9522 25096 9528
rect 24964 9302 25084 9330
rect 24952 9172 25004 9178
rect 24952 9114 25004 9120
rect 24860 8900 24912 8906
rect 24860 8842 24912 8848
rect 24964 7886 24992 9114
rect 25056 8838 25084 9302
rect 25044 8832 25096 8838
rect 25096 8792 25176 8820
rect 25044 8774 25096 8780
rect 25148 8566 25176 8792
rect 25044 8560 25096 8566
rect 25044 8502 25096 8508
rect 25136 8560 25188 8566
rect 25136 8502 25188 8508
rect 24952 7880 25004 7886
rect 24952 7822 25004 7828
rect 25056 6662 25084 8502
rect 25240 8498 25268 9540
rect 25228 8492 25280 8498
rect 25228 8434 25280 8440
rect 25332 7426 25360 21422
rect 25424 20398 25452 28494
rect 25516 27470 25544 28698
rect 25608 28558 25636 36586
rect 25700 33658 25728 38150
rect 25792 36242 25820 38694
rect 25872 38276 25924 38282
rect 25872 38218 25924 38224
rect 25884 37806 25912 38218
rect 25976 37874 26004 39510
rect 25964 37868 26016 37874
rect 25964 37810 26016 37816
rect 25872 37800 25924 37806
rect 25872 37742 25924 37748
rect 25976 37262 26004 37810
rect 26068 37262 26096 40598
rect 26252 40526 26280 41958
rect 26424 41608 26476 41614
rect 26424 41550 26476 41556
rect 26332 40928 26384 40934
rect 26332 40870 26384 40876
rect 26240 40520 26292 40526
rect 26240 40462 26292 40468
rect 26252 40186 26280 40462
rect 26240 40180 26292 40186
rect 26240 40122 26292 40128
rect 26240 39432 26292 39438
rect 26240 39374 26292 39380
rect 26252 38486 26280 39374
rect 26344 39370 26372 40870
rect 26436 40730 26464 41550
rect 26620 41414 26648 42094
rect 26620 41386 27016 41414
rect 26424 40724 26476 40730
rect 26424 40666 26476 40672
rect 26332 39364 26384 39370
rect 26332 39306 26384 39312
rect 26240 38480 26292 38486
rect 26240 38422 26292 38428
rect 26148 38344 26200 38350
rect 26148 38286 26200 38292
rect 26160 38010 26188 38286
rect 26148 38004 26200 38010
rect 26148 37946 26200 37952
rect 26252 37398 26280 38422
rect 26332 38208 26384 38214
rect 26332 38150 26384 38156
rect 26344 37942 26372 38150
rect 26516 38004 26568 38010
rect 26516 37946 26568 37952
rect 26332 37936 26384 37942
rect 26332 37878 26384 37884
rect 26240 37392 26292 37398
rect 26240 37334 26292 37340
rect 25964 37256 26016 37262
rect 25964 37198 26016 37204
rect 26056 37256 26108 37262
rect 26056 37198 26108 37204
rect 26148 36780 26200 36786
rect 26148 36722 26200 36728
rect 26056 36576 26108 36582
rect 26056 36518 26108 36524
rect 26068 36258 26096 36518
rect 26160 36378 26188 36722
rect 26148 36372 26200 36378
rect 26148 36314 26200 36320
rect 25780 36236 25832 36242
rect 26068 36230 26188 36258
rect 25780 36178 25832 36184
rect 26056 36100 26108 36106
rect 26056 36042 26108 36048
rect 25780 35488 25832 35494
rect 25780 35430 25832 35436
rect 25792 35086 25820 35430
rect 26068 35290 26096 36042
rect 26160 35290 26188 36230
rect 26528 36038 26556 37946
rect 26516 36032 26568 36038
rect 26516 35974 26568 35980
rect 26332 35488 26384 35494
rect 26332 35430 26384 35436
rect 26056 35284 26108 35290
rect 26056 35226 26108 35232
rect 26148 35284 26200 35290
rect 26148 35226 26200 35232
rect 25964 35148 26016 35154
rect 25964 35090 26016 35096
rect 25780 35080 25832 35086
rect 25780 35022 25832 35028
rect 25976 34678 26004 35090
rect 25964 34672 26016 34678
rect 25964 34614 26016 34620
rect 25780 34604 25832 34610
rect 25780 34546 25832 34552
rect 25792 34202 25820 34546
rect 25780 34196 25832 34202
rect 25780 34138 25832 34144
rect 25780 33992 25832 33998
rect 25780 33934 25832 33940
rect 25688 33652 25740 33658
rect 25688 33594 25740 33600
rect 25792 33114 25820 33934
rect 26160 33318 26188 35226
rect 26240 35216 26292 35222
rect 26240 35158 26292 35164
rect 26252 34610 26280 35158
rect 26344 35086 26372 35430
rect 26528 35086 26556 35974
rect 26620 35698 26648 41386
rect 26988 40662 27016 41386
rect 26976 40656 27028 40662
rect 26976 40598 27028 40604
rect 26700 40520 26752 40526
rect 26976 40520 27028 40526
rect 26700 40462 26752 40468
rect 26896 40468 26976 40474
rect 26896 40462 27028 40468
rect 26712 40118 26740 40462
rect 26896 40446 27016 40462
rect 26896 40186 26924 40446
rect 27172 40186 27200 42162
rect 27344 42152 27396 42158
rect 27344 42094 27396 42100
rect 27252 42016 27304 42022
rect 27252 41958 27304 41964
rect 27264 41206 27292 41958
rect 27252 41200 27304 41206
rect 27252 41142 27304 41148
rect 27356 40934 27384 42094
rect 27620 42084 27672 42090
rect 27620 42026 27672 42032
rect 27632 41818 27660 42026
rect 27620 41812 27672 41818
rect 27620 41754 27672 41760
rect 27620 41608 27672 41614
rect 27620 41550 27672 41556
rect 27632 41138 27660 41550
rect 27894 41370 27950 42406
rect 29748 42226 29776 42570
rect 30104 42560 30156 42566
rect 30104 42502 30156 42508
rect 28632 42220 28684 42226
rect 28632 42162 28684 42168
rect 29736 42220 29788 42226
rect 29736 42162 29788 42168
rect 28540 42084 28592 42090
rect 28540 42026 28592 42032
rect 28448 42016 28500 42022
rect 28448 41958 28500 41964
rect 28460 41614 28488 41958
rect 28448 41608 28500 41614
rect 28448 41550 28500 41556
rect 28356 41540 28408 41546
rect 28356 41482 28408 41488
rect 27894 41318 27896 41370
rect 27948 41318 27950 41370
rect 27620 41132 27672 41138
rect 27620 41074 27672 41080
rect 27344 40928 27396 40934
rect 27344 40870 27396 40876
rect 27712 40928 27764 40934
rect 27712 40870 27764 40876
rect 27356 40594 27384 40870
rect 27344 40588 27396 40594
rect 27344 40530 27396 40536
rect 26884 40180 26936 40186
rect 26884 40122 26936 40128
rect 27160 40180 27212 40186
rect 27160 40122 27212 40128
rect 26700 40112 26752 40118
rect 26700 40054 26752 40060
rect 27724 40050 27752 40870
rect 27804 40520 27856 40526
rect 27804 40462 27856 40468
rect 27816 40118 27844 40462
rect 27894 40282 27950 41318
rect 28264 40520 28316 40526
rect 28264 40462 28316 40468
rect 28080 40452 28132 40458
rect 28080 40394 28132 40400
rect 27894 40230 27896 40282
rect 27948 40230 27950 40282
rect 27804 40112 27856 40118
rect 27804 40054 27856 40060
rect 27712 40044 27764 40050
rect 27712 39986 27764 39992
rect 27160 39296 27212 39302
rect 27160 39238 27212 39244
rect 27172 38350 27200 39238
rect 27620 38956 27672 38962
rect 27620 38898 27672 38904
rect 27632 38554 27660 38898
rect 27620 38548 27672 38554
rect 27620 38490 27672 38496
rect 27068 38344 27120 38350
rect 27068 38286 27120 38292
rect 27160 38344 27212 38350
rect 27160 38286 27212 38292
rect 26976 37868 27028 37874
rect 26976 37810 27028 37816
rect 26988 37346 27016 37810
rect 27080 37466 27108 38286
rect 27436 38208 27488 38214
rect 27436 38150 27488 38156
rect 27448 38010 27476 38150
rect 27436 38004 27488 38010
rect 27436 37946 27488 37952
rect 27344 37902 27396 37908
rect 27252 37868 27304 37874
rect 27632 37874 27660 38490
rect 27724 38486 27752 39986
rect 27816 39506 27844 40054
rect 27804 39500 27856 39506
rect 27804 39442 27856 39448
rect 27894 39194 27950 40230
rect 28092 40186 28120 40394
rect 28080 40180 28132 40186
rect 28080 40122 28132 40128
rect 28276 39914 28304 40462
rect 28264 39908 28316 39914
rect 28264 39850 28316 39856
rect 27894 39142 27896 39194
rect 27948 39142 27950 39194
rect 27804 38752 27856 38758
rect 27804 38694 27856 38700
rect 27816 38554 27844 38694
rect 27804 38548 27856 38554
rect 27804 38490 27856 38496
rect 27712 38480 27764 38486
rect 27712 38422 27764 38428
rect 27804 38344 27856 38350
rect 27804 38286 27856 38292
rect 27344 37844 27396 37850
rect 27620 37868 27672 37874
rect 27252 37810 27304 37816
rect 27068 37460 27120 37466
rect 27068 37402 27120 37408
rect 27160 37460 27212 37466
rect 27160 37402 27212 37408
rect 27172 37346 27200 37402
rect 27264 37398 27292 37810
rect 26988 37318 27200 37346
rect 27252 37392 27304 37398
rect 27252 37334 27304 37340
rect 26792 37256 26844 37262
rect 26792 37198 26844 37204
rect 26804 36718 26832 37198
rect 27160 37120 27212 37126
rect 27160 37062 27212 37068
rect 27172 36786 27200 37062
rect 27356 36922 27384 37844
rect 27620 37810 27672 37816
rect 27816 37806 27844 38286
rect 27894 38106 27950 39142
rect 28368 38826 28396 41482
rect 28552 41414 28580 42026
rect 28460 41386 28580 41414
rect 28460 40526 28488 41386
rect 28448 40520 28500 40526
rect 28448 40462 28500 40468
rect 28448 40384 28500 40390
rect 28448 40326 28500 40332
rect 28460 38962 28488 40326
rect 28644 40186 28672 42162
rect 28816 42152 28868 42158
rect 28816 42094 28868 42100
rect 28828 41290 28856 42094
rect 29368 42084 29420 42090
rect 29368 42026 29420 42032
rect 28828 41262 29040 41290
rect 28724 41132 28776 41138
rect 28724 41074 28776 41080
rect 28908 41132 28960 41138
rect 28908 41074 28960 41080
rect 28736 40594 28764 41074
rect 28816 40928 28868 40934
rect 28816 40870 28868 40876
rect 28828 40610 28856 40870
rect 28920 40730 28948 41074
rect 29012 40934 29040 41262
rect 29000 40928 29052 40934
rect 29000 40870 29052 40876
rect 28908 40724 28960 40730
rect 28908 40666 28960 40672
rect 28724 40588 28776 40594
rect 28828 40582 28948 40610
rect 28724 40530 28776 40536
rect 28920 40526 28948 40582
rect 28816 40520 28868 40526
rect 28816 40462 28868 40468
rect 28908 40520 28960 40526
rect 28908 40462 28960 40468
rect 28632 40180 28684 40186
rect 28632 40122 28684 40128
rect 28724 40044 28776 40050
rect 28724 39986 28776 39992
rect 28632 39432 28684 39438
rect 28632 39374 28684 39380
rect 28448 38956 28500 38962
rect 28448 38898 28500 38904
rect 28356 38820 28408 38826
rect 28356 38762 28408 38768
rect 27988 38344 28040 38350
rect 28644 38332 28672 39374
rect 28736 39098 28764 39986
rect 28828 39914 28856 40462
rect 29012 40372 29040 40870
rect 28920 40344 29040 40372
rect 28920 40050 28948 40344
rect 28908 40044 28960 40050
rect 28908 39986 28960 39992
rect 28816 39908 28868 39914
rect 28816 39850 28868 39856
rect 28724 39092 28776 39098
rect 28724 39034 28776 39040
rect 28828 38962 28856 39850
rect 29184 39364 29236 39370
rect 29184 39306 29236 39312
rect 28816 38956 28868 38962
rect 28816 38898 28868 38904
rect 29196 38894 29224 39306
rect 29184 38888 29236 38894
rect 29184 38830 29236 38836
rect 28724 38344 28776 38350
rect 28644 38304 28724 38332
rect 27988 38286 28040 38292
rect 28724 38286 28776 38292
rect 27894 38054 27896 38106
rect 27948 38054 27950 38106
rect 27804 37800 27856 37806
rect 27804 37742 27856 37748
rect 27620 37392 27672 37398
rect 27620 37334 27672 37340
rect 27436 37256 27488 37262
rect 27436 37198 27488 37204
rect 27344 36916 27396 36922
rect 27344 36858 27396 36864
rect 27160 36780 27212 36786
rect 27160 36722 27212 36728
rect 26792 36712 26844 36718
rect 26792 36654 26844 36660
rect 26792 36576 26844 36582
rect 26792 36518 26844 36524
rect 26804 36242 26832 36518
rect 27356 36310 27384 36858
rect 27448 36582 27476 37198
rect 27632 37194 27660 37334
rect 27620 37188 27672 37194
rect 27620 37130 27672 37136
rect 27804 37188 27856 37194
rect 27804 37130 27856 37136
rect 27436 36576 27488 36582
rect 27436 36518 27488 36524
rect 27344 36304 27396 36310
rect 27344 36246 27396 36252
rect 26792 36236 26844 36242
rect 26792 36178 26844 36184
rect 27160 36168 27212 36174
rect 27160 36110 27212 36116
rect 27172 35698 27200 36110
rect 27356 35766 27384 36246
rect 27436 36100 27488 36106
rect 27436 36042 27488 36048
rect 27344 35760 27396 35766
rect 27344 35702 27396 35708
rect 27448 35698 27476 36042
rect 27816 35894 27844 37130
rect 27724 35866 27844 35894
rect 27894 37018 27950 38054
rect 28000 37330 28028 38286
rect 28736 37670 28764 38286
rect 28724 37664 28776 37670
rect 28724 37606 28776 37612
rect 29000 37664 29052 37670
rect 29000 37606 29052 37612
rect 28724 37392 28776 37398
rect 29012 37380 29040 37606
rect 29196 37466 29224 38830
rect 29184 37460 29236 37466
rect 29184 37402 29236 37408
rect 28776 37352 29040 37380
rect 28724 37334 28776 37340
rect 27988 37324 28040 37330
rect 27988 37266 28040 37272
rect 29012 37262 29040 37352
rect 28816 37256 28868 37262
rect 28816 37198 28868 37204
rect 29000 37256 29052 37262
rect 29000 37198 29052 37204
rect 27894 36966 27896 37018
rect 27948 36966 27950 37018
rect 27894 35930 27950 36966
rect 28828 36922 28856 37198
rect 28954 37120 29006 37126
rect 29006 37080 29316 37108
rect 28954 37062 29006 37068
rect 28816 36916 28868 36922
rect 28816 36858 28868 36864
rect 29000 36848 29052 36854
rect 29000 36790 29052 36796
rect 28908 36644 28960 36650
rect 28908 36586 28960 36592
rect 28632 36576 28684 36582
rect 28552 36536 28632 36564
rect 28552 36174 28580 36536
rect 28632 36518 28684 36524
rect 28920 36378 28948 36586
rect 28908 36372 28960 36378
rect 28908 36314 28960 36320
rect 28540 36168 28592 36174
rect 28540 36110 28592 36116
rect 28632 36168 28684 36174
rect 28632 36110 28684 36116
rect 28264 36032 28316 36038
rect 28264 35974 28316 35980
rect 27894 35878 27896 35930
rect 27948 35878 27950 35930
rect 26608 35692 26660 35698
rect 26608 35634 26660 35640
rect 27160 35692 27212 35698
rect 27160 35634 27212 35640
rect 27436 35692 27488 35698
rect 27436 35634 27488 35640
rect 26332 35080 26384 35086
rect 26332 35022 26384 35028
rect 26516 35080 26568 35086
rect 26516 35022 26568 35028
rect 26240 34604 26292 34610
rect 26240 34546 26292 34552
rect 26148 33312 26200 33318
rect 26148 33254 26200 33260
rect 25780 33108 25832 33114
rect 25780 33050 25832 33056
rect 26056 32904 26108 32910
rect 26056 32846 26108 32852
rect 25872 32224 25924 32230
rect 25872 32166 25924 32172
rect 25688 31952 25740 31958
rect 25688 31894 25740 31900
rect 25700 29714 25728 31894
rect 25884 31804 25912 32166
rect 25964 31816 26016 31822
rect 25884 31776 25964 31804
rect 25884 31278 25912 31776
rect 25964 31758 26016 31764
rect 25964 31340 26016 31346
rect 25964 31282 26016 31288
rect 25872 31272 25924 31278
rect 25872 31214 25924 31220
rect 25780 30048 25832 30054
rect 25780 29990 25832 29996
rect 25688 29708 25740 29714
rect 25688 29650 25740 29656
rect 25700 28966 25728 29650
rect 25792 29646 25820 29990
rect 25780 29640 25832 29646
rect 25780 29582 25832 29588
rect 25688 28960 25740 28966
rect 25688 28902 25740 28908
rect 25688 28688 25740 28694
rect 25688 28630 25740 28636
rect 25792 28642 25820 29582
rect 25884 29238 25912 31214
rect 25976 30938 26004 31282
rect 26068 31210 26096 32846
rect 26332 32836 26384 32842
rect 26332 32778 26384 32784
rect 26240 32224 26292 32230
rect 26240 32166 26292 32172
rect 26252 32026 26280 32166
rect 26240 32020 26292 32026
rect 26240 31962 26292 31968
rect 26344 31890 26372 32778
rect 26516 32496 26568 32502
rect 26516 32438 26568 32444
rect 26528 31890 26556 32438
rect 26332 31884 26384 31890
rect 26332 31826 26384 31832
rect 26516 31884 26568 31890
rect 26516 31826 26568 31832
rect 26148 31340 26200 31346
rect 26148 31282 26200 31288
rect 26056 31204 26108 31210
rect 26056 31146 26108 31152
rect 25964 30932 26016 30938
rect 25964 30874 26016 30880
rect 25964 29640 26016 29646
rect 25964 29582 26016 29588
rect 25872 29232 25924 29238
rect 25872 29174 25924 29180
rect 25976 28966 26004 29582
rect 26056 29572 26108 29578
rect 26160 29560 26188 31282
rect 26344 30802 26372 31826
rect 26424 31748 26476 31754
rect 26424 31690 26476 31696
rect 26332 30796 26384 30802
rect 26332 30738 26384 30744
rect 26240 30728 26292 30734
rect 26240 30670 26292 30676
rect 26252 30138 26280 30670
rect 26344 30258 26372 30738
rect 26436 30734 26464 31690
rect 26424 30728 26476 30734
rect 26424 30670 26476 30676
rect 26436 30394 26464 30670
rect 26424 30388 26476 30394
rect 26424 30330 26476 30336
rect 26332 30252 26384 30258
rect 26332 30194 26384 30200
rect 26424 30252 26476 30258
rect 26424 30194 26476 30200
rect 26252 30110 26372 30138
rect 26108 29532 26188 29560
rect 26056 29514 26108 29520
rect 25964 28960 26016 28966
rect 25964 28902 26016 28908
rect 25596 28552 25648 28558
rect 25596 28494 25648 28500
rect 25700 28082 25728 28630
rect 25792 28614 25912 28642
rect 25780 28552 25832 28558
rect 25780 28494 25832 28500
rect 25688 28076 25740 28082
rect 25688 28018 25740 28024
rect 25792 28014 25820 28494
rect 25884 28082 25912 28614
rect 25964 28484 26016 28490
rect 25964 28426 26016 28432
rect 25872 28076 25924 28082
rect 25872 28018 25924 28024
rect 25780 28008 25832 28014
rect 25780 27950 25832 27956
rect 25596 27940 25648 27946
rect 25596 27882 25648 27888
rect 25608 27606 25636 27882
rect 25884 27674 25912 28018
rect 25872 27668 25924 27674
rect 25872 27610 25924 27616
rect 25596 27600 25648 27606
rect 25596 27542 25648 27548
rect 25688 27532 25740 27538
rect 25688 27474 25740 27480
rect 25504 27464 25556 27470
rect 25504 27406 25556 27412
rect 25504 24812 25556 24818
rect 25504 24754 25556 24760
rect 25516 23730 25544 24754
rect 25504 23724 25556 23730
rect 25504 23666 25556 23672
rect 25596 23724 25648 23730
rect 25596 23666 25648 23672
rect 25608 22438 25636 23666
rect 25700 23032 25728 27474
rect 25872 27056 25924 27062
rect 25976 27044 26004 28426
rect 25924 27016 26004 27044
rect 25872 26998 25924 27004
rect 25872 24676 25924 24682
rect 25872 24618 25924 24624
rect 25884 24410 25912 24618
rect 25872 24404 25924 24410
rect 25872 24346 25924 24352
rect 25872 23588 25924 23594
rect 25872 23530 25924 23536
rect 25780 23044 25832 23050
rect 25700 23004 25780 23032
rect 25780 22986 25832 22992
rect 25792 22642 25820 22986
rect 25780 22636 25832 22642
rect 25780 22578 25832 22584
rect 25596 22432 25648 22438
rect 25596 22374 25648 22380
rect 25608 21486 25636 22374
rect 25688 22024 25740 22030
rect 25740 21972 25820 21978
rect 25688 21966 25820 21972
rect 25700 21950 25820 21966
rect 25596 21480 25648 21486
rect 25596 21422 25648 21428
rect 25412 20392 25464 20398
rect 25412 20334 25464 20340
rect 25596 20392 25648 20398
rect 25596 20334 25648 20340
rect 25424 19394 25452 20334
rect 25608 19514 25636 20334
rect 25792 19854 25820 21950
rect 25780 19848 25832 19854
rect 25780 19790 25832 19796
rect 25596 19508 25648 19514
rect 25596 19450 25648 19456
rect 25688 19508 25740 19514
rect 25688 19450 25740 19456
rect 25700 19394 25728 19450
rect 25792 19446 25820 19790
rect 25424 19366 25728 19394
rect 25780 19440 25832 19446
rect 25780 19382 25832 19388
rect 25424 12434 25452 19366
rect 25688 18964 25740 18970
rect 25688 18906 25740 18912
rect 25504 18080 25556 18086
rect 25504 18022 25556 18028
rect 25516 17746 25544 18022
rect 25596 17876 25648 17882
rect 25596 17818 25648 17824
rect 25504 17740 25556 17746
rect 25504 17682 25556 17688
rect 25516 13938 25544 17682
rect 25608 15706 25636 17818
rect 25596 15700 25648 15706
rect 25596 15642 25648 15648
rect 25596 15496 25648 15502
rect 25596 15438 25648 15444
rect 25608 15094 25636 15438
rect 25596 15088 25648 15094
rect 25596 15030 25648 15036
rect 25504 13932 25556 13938
rect 25504 13874 25556 13880
rect 25516 13530 25544 13874
rect 25504 13524 25556 13530
rect 25504 13466 25556 13472
rect 25516 12918 25544 13466
rect 25700 13258 25728 18906
rect 25792 18766 25820 19382
rect 25884 19310 25912 23530
rect 25964 21956 26016 21962
rect 25964 21898 26016 21904
rect 25976 21690 26004 21898
rect 25964 21684 26016 21690
rect 25964 21626 26016 21632
rect 26068 20346 26096 29514
rect 26148 28552 26200 28558
rect 26148 28494 26200 28500
rect 26160 27402 26188 28494
rect 26240 28008 26292 28014
rect 26240 27950 26292 27956
rect 26252 27674 26280 27950
rect 26240 27668 26292 27674
rect 26240 27610 26292 27616
rect 26344 27554 26372 30110
rect 26436 29510 26464 30194
rect 26528 29714 26556 31826
rect 26620 31142 26648 35634
rect 27252 35556 27304 35562
rect 27252 35498 27304 35504
rect 27264 35222 27292 35498
rect 27252 35216 27304 35222
rect 27252 35158 27304 35164
rect 26792 35080 26844 35086
rect 26792 35022 26844 35028
rect 26700 32904 26752 32910
rect 26700 32846 26752 32852
rect 26712 31754 26740 32846
rect 26804 32434 26832 35022
rect 27448 35018 27476 35634
rect 27436 35012 27488 35018
rect 27436 34954 27488 34960
rect 27160 34944 27212 34950
rect 27160 34886 27212 34892
rect 27172 33522 27200 34886
rect 27448 34626 27476 34954
rect 27356 34610 27476 34626
rect 27344 34604 27476 34610
rect 27396 34598 27476 34604
rect 27344 34546 27396 34552
rect 27160 33516 27212 33522
rect 27160 33458 27212 33464
rect 27620 33516 27672 33522
rect 27620 33458 27672 33464
rect 27068 33448 27120 33454
rect 27068 33390 27120 33396
rect 27080 32910 27108 33390
rect 27172 32978 27200 33458
rect 27632 33046 27660 33458
rect 27620 33040 27672 33046
rect 27620 32982 27672 32988
rect 27160 32972 27212 32978
rect 27160 32914 27212 32920
rect 27528 32972 27580 32978
rect 27528 32914 27580 32920
rect 27068 32904 27120 32910
rect 27068 32846 27120 32852
rect 27540 32774 27568 32914
rect 27528 32768 27580 32774
rect 27528 32710 27580 32716
rect 27540 32434 27568 32710
rect 26792 32428 26844 32434
rect 26792 32370 26844 32376
rect 27528 32428 27580 32434
rect 27528 32370 27580 32376
rect 26700 31748 26752 31754
rect 26700 31690 26752 31696
rect 26804 31210 26832 32370
rect 27632 32298 27660 32982
rect 27724 32570 27752 35866
rect 27894 34842 27950 35878
rect 28172 35692 28224 35698
rect 28172 35634 28224 35640
rect 28080 35488 28132 35494
rect 28080 35430 28132 35436
rect 28092 35018 28120 35430
rect 28080 35012 28132 35018
rect 28080 34954 28132 34960
rect 27894 34790 27896 34842
rect 27948 34790 27950 34842
rect 27804 33856 27856 33862
rect 27804 33798 27856 33804
rect 27816 32910 27844 33798
rect 27894 33754 27950 34790
rect 27894 33702 27896 33754
rect 27948 33702 27950 33754
rect 27804 32904 27856 32910
rect 27804 32846 27856 32852
rect 27894 32666 27950 33702
rect 28092 32842 28120 34954
rect 28184 34746 28212 35634
rect 28276 35494 28304 35974
rect 28540 35760 28592 35766
rect 28540 35702 28592 35708
rect 28448 35624 28500 35630
rect 28448 35566 28500 35572
rect 28264 35488 28316 35494
rect 28264 35430 28316 35436
rect 28172 34740 28224 34746
rect 28172 34682 28224 34688
rect 28460 34610 28488 35566
rect 28448 34604 28500 34610
rect 28448 34546 28500 34552
rect 28172 33312 28224 33318
rect 28172 33254 28224 33260
rect 28080 32836 28132 32842
rect 27894 32614 27896 32666
rect 27948 32614 27950 32666
rect 27712 32564 27764 32570
rect 27712 32506 27764 32512
rect 27528 32292 27580 32298
rect 27528 32234 27580 32240
rect 27620 32292 27672 32298
rect 27620 32234 27672 32240
rect 27540 31890 27568 32234
rect 27632 32026 27660 32234
rect 27620 32020 27672 32026
rect 27620 31962 27672 31968
rect 27528 31884 27580 31890
rect 27528 31826 27580 31832
rect 26792 31204 26844 31210
rect 26792 31146 26844 31152
rect 26608 31136 26660 31142
rect 26608 31078 26660 31084
rect 26620 30852 26648 31078
rect 26620 30824 26740 30852
rect 26608 30116 26660 30122
rect 26608 30058 26660 30064
rect 26516 29708 26568 29714
rect 26516 29650 26568 29656
rect 26620 29578 26648 30058
rect 26712 29850 26740 30824
rect 26700 29844 26752 29850
rect 26700 29786 26752 29792
rect 26608 29572 26660 29578
rect 26608 29514 26660 29520
rect 26424 29504 26476 29510
rect 26424 29446 26476 29452
rect 26436 28422 26464 29446
rect 26516 29028 26568 29034
rect 26516 28970 26568 28976
rect 26424 28416 26476 28422
rect 26424 28358 26476 28364
rect 26252 27526 26372 27554
rect 26148 27396 26200 27402
rect 26148 27338 26200 27344
rect 26252 23730 26280 27526
rect 26332 27056 26384 27062
rect 26332 26998 26384 27004
rect 26344 26246 26372 26998
rect 26436 26926 26464 28358
rect 26424 26920 26476 26926
rect 26424 26862 26476 26868
rect 26528 26246 26556 28970
rect 26804 28370 26832 31146
rect 27724 30326 27752 32506
rect 27894 31578 27950 32614
rect 27894 31526 27896 31578
rect 27948 31526 27950 31578
rect 27894 30490 27950 31526
rect 28000 32796 28080 32824
rect 28000 31346 28028 32796
rect 28080 32778 28132 32784
rect 28080 32564 28132 32570
rect 28080 32506 28132 32512
rect 27988 31340 28040 31346
rect 27988 31282 28040 31288
rect 28000 30734 28028 31282
rect 27988 30728 28040 30734
rect 27988 30670 28040 30676
rect 27894 30438 27896 30490
rect 27948 30438 27950 30490
rect 27712 30320 27764 30326
rect 27712 30262 27764 30268
rect 27344 30184 27396 30190
rect 27344 30126 27396 30132
rect 27356 29102 27384 30126
rect 27528 30048 27580 30054
rect 27528 29990 27580 29996
rect 27540 29646 27568 29990
rect 27528 29640 27580 29646
rect 27528 29582 27580 29588
rect 27160 29096 27212 29102
rect 27160 29038 27212 29044
rect 27344 29096 27396 29102
rect 27344 29038 27396 29044
rect 27540 29050 27568 29582
rect 27894 29402 27950 30438
rect 27894 29350 27896 29402
rect 27948 29350 27950 29402
rect 26884 28960 26936 28966
rect 26884 28902 26936 28908
rect 26896 28762 26924 28902
rect 26884 28756 26936 28762
rect 26884 28698 26936 28704
rect 26620 28342 26832 28370
rect 26332 26240 26384 26246
rect 26332 26182 26384 26188
rect 26516 26240 26568 26246
rect 26516 26182 26568 26188
rect 26344 25294 26372 26182
rect 26528 25294 26556 26182
rect 26332 25288 26384 25294
rect 26516 25288 26568 25294
rect 26384 25236 26464 25242
rect 26332 25230 26464 25236
rect 26516 25230 26568 25236
rect 26344 25214 26464 25230
rect 26240 23724 26292 23730
rect 26240 23666 26292 23672
rect 26436 23662 26464 25214
rect 26528 24886 26556 25230
rect 26516 24880 26568 24886
rect 26516 24822 26568 24828
rect 26424 23656 26476 23662
rect 26424 23598 26476 23604
rect 26240 23520 26292 23526
rect 26240 23462 26292 23468
rect 26148 22976 26200 22982
rect 26148 22918 26200 22924
rect 26160 21554 26188 22918
rect 26148 21548 26200 21554
rect 26148 21490 26200 21496
rect 26148 20800 26200 20806
rect 26148 20742 26200 20748
rect 25976 20318 26096 20346
rect 25872 19304 25924 19310
rect 25872 19246 25924 19252
rect 25780 18760 25832 18766
rect 25780 18702 25832 18708
rect 25792 17542 25820 18702
rect 25872 18284 25924 18290
rect 25872 18226 25924 18232
rect 25780 17536 25832 17542
rect 25780 17478 25832 17484
rect 25780 16584 25832 16590
rect 25780 16526 25832 16532
rect 25792 15366 25820 16526
rect 25780 15360 25832 15366
rect 25780 15302 25832 15308
rect 25792 13938 25820 15302
rect 25780 13932 25832 13938
rect 25780 13874 25832 13880
rect 25792 13530 25820 13874
rect 25780 13524 25832 13530
rect 25780 13466 25832 13472
rect 25688 13252 25740 13258
rect 25688 13194 25740 13200
rect 25504 12912 25556 12918
rect 25504 12854 25556 12860
rect 25700 12850 25728 13194
rect 25884 12850 25912 18226
rect 25976 17882 26004 20318
rect 26056 20256 26108 20262
rect 26056 20198 26108 20204
rect 26068 18766 26096 20198
rect 26160 19854 26188 20742
rect 26252 20058 26280 23462
rect 26436 22778 26464 23598
rect 26424 22772 26476 22778
rect 26424 22714 26476 22720
rect 26424 21684 26476 21690
rect 26424 21626 26476 21632
rect 26436 21010 26464 21626
rect 26516 21344 26568 21350
rect 26516 21286 26568 21292
rect 26424 21004 26476 21010
rect 26424 20946 26476 20952
rect 26528 20942 26556 21286
rect 26516 20936 26568 20942
rect 26516 20878 26568 20884
rect 26332 20256 26384 20262
rect 26332 20198 26384 20204
rect 26240 20052 26292 20058
rect 26240 19994 26292 20000
rect 26148 19848 26200 19854
rect 26148 19790 26200 19796
rect 26344 19334 26372 20198
rect 26344 19306 26556 19334
rect 26148 19168 26200 19174
rect 26148 19110 26200 19116
rect 26056 18760 26108 18766
rect 26056 18702 26108 18708
rect 26160 18426 26188 19110
rect 26148 18420 26200 18426
rect 26148 18362 26200 18368
rect 26148 18080 26200 18086
rect 26148 18022 26200 18028
rect 26160 17882 26188 18022
rect 25964 17876 26016 17882
rect 25964 17818 26016 17824
rect 26148 17876 26200 17882
rect 26148 17818 26200 17824
rect 26056 17672 26108 17678
rect 26056 17614 26108 17620
rect 26068 16998 26096 17614
rect 26148 17604 26200 17610
rect 26148 17546 26200 17552
rect 26056 16992 26108 16998
rect 26056 16934 26108 16940
rect 26068 16794 26096 16934
rect 26056 16788 26108 16794
rect 26056 16730 26108 16736
rect 26160 16658 26188 17546
rect 26148 16652 26200 16658
rect 26148 16594 26200 16600
rect 26056 16448 26108 16454
rect 26056 16390 26108 16396
rect 26068 16114 26096 16390
rect 25964 16108 26016 16114
rect 25964 16050 26016 16056
rect 26056 16108 26108 16114
rect 26056 16050 26108 16056
rect 25976 14618 26004 16050
rect 26160 15994 26188 16594
rect 26068 15966 26188 15994
rect 25964 14612 26016 14618
rect 25964 14554 26016 14560
rect 25964 14476 26016 14482
rect 25964 14418 26016 14424
rect 25976 14074 26004 14418
rect 25964 14068 26016 14074
rect 25964 14010 26016 14016
rect 25964 13456 26016 13462
rect 25964 13398 26016 13404
rect 25976 12986 26004 13398
rect 25964 12980 26016 12986
rect 25964 12922 26016 12928
rect 25688 12844 25740 12850
rect 25688 12786 25740 12792
rect 25872 12844 25924 12850
rect 25872 12786 25924 12792
rect 25964 12640 26016 12646
rect 25964 12582 26016 12588
rect 25424 12406 25636 12434
rect 25412 12164 25464 12170
rect 25412 12106 25464 12112
rect 25424 11830 25452 12106
rect 25412 11824 25464 11830
rect 25412 11766 25464 11772
rect 25504 11076 25556 11082
rect 25504 11018 25556 11024
rect 25516 9654 25544 11018
rect 25504 9648 25556 9654
rect 25504 9590 25556 9596
rect 25608 9586 25636 12406
rect 25976 12238 26004 12582
rect 25964 12232 26016 12238
rect 25964 12174 26016 12180
rect 26068 11558 26096 15966
rect 26240 15904 26292 15910
rect 26240 15846 26292 15852
rect 26252 15076 26280 15846
rect 26332 15088 26384 15094
rect 26252 15048 26332 15076
rect 26148 15020 26200 15026
rect 26148 14962 26200 14968
rect 26160 14006 26188 14962
rect 26252 14550 26280 15048
rect 26332 15030 26384 15036
rect 26240 14544 26292 14550
rect 26240 14486 26292 14492
rect 26332 14544 26384 14550
rect 26332 14486 26384 14492
rect 26240 14408 26292 14414
rect 26240 14350 26292 14356
rect 26148 14000 26200 14006
rect 26148 13942 26200 13948
rect 26148 12776 26200 12782
rect 26148 12718 26200 12724
rect 26056 11552 26108 11558
rect 26056 11494 26108 11500
rect 25688 11144 25740 11150
rect 25688 11086 25740 11092
rect 25872 11144 25924 11150
rect 25872 11086 25924 11092
rect 25700 10810 25728 11086
rect 25688 10804 25740 10810
rect 25688 10746 25740 10752
rect 25884 10470 25912 11086
rect 25964 11008 26016 11014
rect 25964 10950 26016 10956
rect 25976 10674 26004 10950
rect 25964 10668 26016 10674
rect 25964 10610 26016 10616
rect 25872 10464 25924 10470
rect 25872 10406 25924 10412
rect 25596 9580 25648 9586
rect 25596 9522 25648 9528
rect 25780 9580 25832 9586
rect 25780 9522 25832 9528
rect 25792 8430 25820 9522
rect 25884 9110 25912 10406
rect 25964 10260 26016 10266
rect 25964 10202 26016 10208
rect 25976 9382 26004 10202
rect 25964 9376 26016 9382
rect 25964 9318 26016 9324
rect 25872 9104 25924 9110
rect 25872 9046 25924 9052
rect 25964 8832 26016 8838
rect 25964 8774 26016 8780
rect 25780 8424 25832 8430
rect 25780 8366 25832 8372
rect 25596 8288 25648 8294
rect 25596 8230 25648 8236
rect 25608 7886 25636 8230
rect 25596 7880 25648 7886
rect 25596 7822 25648 7828
rect 25780 7744 25832 7750
rect 25780 7686 25832 7692
rect 25148 7410 25360 7426
rect 25136 7404 25360 7410
rect 25188 7398 25360 7404
rect 25136 7346 25188 7352
rect 25504 7200 25556 7206
rect 25504 7142 25556 7148
rect 25516 6866 25544 7142
rect 25504 6860 25556 6866
rect 25504 6802 25556 6808
rect 25044 6656 25096 6662
rect 25044 6598 25096 6604
rect 25792 6322 25820 7686
rect 25976 7002 26004 8774
rect 26068 8566 26096 11494
rect 26160 10810 26188 12718
rect 26148 10804 26200 10810
rect 26148 10746 26200 10752
rect 26252 10674 26280 14350
rect 26344 13190 26372 14486
rect 26528 13530 26556 19306
rect 26620 17814 26648 28342
rect 26896 27946 26924 28698
rect 27068 28416 27120 28422
rect 27068 28358 27120 28364
rect 27080 28082 27108 28358
rect 27068 28076 27120 28082
rect 27068 28018 27120 28024
rect 26884 27940 26936 27946
rect 26884 27882 26936 27888
rect 26700 27464 26752 27470
rect 26700 27406 26752 27412
rect 26712 26738 26740 27406
rect 26792 27396 26844 27402
rect 26792 27338 26844 27344
rect 26804 27130 26832 27338
rect 26792 27124 26844 27130
rect 26792 27066 26844 27072
rect 26712 26710 26832 26738
rect 26700 26580 26752 26586
rect 26700 26522 26752 26528
rect 26712 21706 26740 26522
rect 26804 26382 26832 26710
rect 26792 26376 26844 26382
rect 26792 26318 26844 26324
rect 26976 26308 27028 26314
rect 26976 26250 27028 26256
rect 26988 24818 27016 26250
rect 27172 25430 27200 29038
rect 27356 28150 27384 29038
rect 27540 29022 27660 29050
rect 27632 28626 27660 29022
rect 27804 29028 27856 29034
rect 27804 28970 27856 28976
rect 27620 28620 27672 28626
rect 27620 28562 27672 28568
rect 27816 28218 27844 28970
rect 27894 28314 27950 29350
rect 28092 29170 28120 32506
rect 28184 31346 28212 33254
rect 28264 32904 28316 32910
rect 28264 32846 28316 32852
rect 28276 32434 28304 32846
rect 28460 32722 28488 34546
rect 28552 34134 28580 35702
rect 28540 34128 28592 34134
rect 28540 34070 28592 34076
rect 28540 33516 28592 33522
rect 28540 33458 28592 33464
rect 28368 32694 28488 32722
rect 28368 32570 28396 32694
rect 28356 32564 28408 32570
rect 28356 32506 28408 32512
rect 28448 32564 28500 32570
rect 28448 32506 28500 32512
rect 28264 32428 28316 32434
rect 28264 32370 28316 32376
rect 28356 31816 28408 31822
rect 28356 31758 28408 31764
rect 28368 31482 28396 31758
rect 28356 31476 28408 31482
rect 28356 31418 28408 31424
rect 28172 31340 28224 31346
rect 28172 31282 28224 31288
rect 28264 30320 28316 30326
rect 28264 30262 28316 30268
rect 28080 29164 28132 29170
rect 28080 29106 28132 29112
rect 27894 28262 27896 28314
rect 27948 28262 27950 28314
rect 27804 28212 27856 28218
rect 27804 28154 27856 28160
rect 27344 28144 27396 28150
rect 27344 28086 27396 28092
rect 27344 27872 27396 27878
rect 27344 27814 27396 27820
rect 27356 27130 27384 27814
rect 27436 27668 27488 27674
rect 27436 27610 27488 27616
rect 27344 27124 27396 27130
rect 27344 27066 27396 27072
rect 27448 26976 27476 27610
rect 27894 27226 27950 28262
rect 28172 28144 28224 28150
rect 28172 28086 28224 28092
rect 27894 27174 27896 27226
rect 27948 27174 27950 27226
rect 27528 26988 27580 26994
rect 27448 26948 27528 26976
rect 27160 25424 27212 25430
rect 27160 25366 27212 25372
rect 27160 25152 27212 25158
rect 27160 25094 27212 25100
rect 27172 24818 27200 25094
rect 27448 24818 27476 26948
rect 27528 26930 27580 26936
rect 27712 26376 27764 26382
rect 27712 26318 27764 26324
rect 27724 25906 27752 26318
rect 27894 26138 27950 27174
rect 27988 26988 28040 26994
rect 27988 26930 28040 26936
rect 27894 26086 27896 26138
rect 27948 26086 27950 26138
rect 27712 25900 27764 25906
rect 27764 25860 27844 25888
rect 27712 25842 27764 25848
rect 27816 25158 27844 25860
rect 27804 25152 27856 25158
rect 27804 25094 27856 25100
rect 26792 24812 26844 24818
rect 26792 24754 26844 24760
rect 26976 24812 27028 24818
rect 26976 24754 27028 24760
rect 27160 24812 27212 24818
rect 27160 24754 27212 24760
rect 27436 24812 27488 24818
rect 27436 24754 27488 24760
rect 26804 22030 26832 24754
rect 27712 24744 27764 24750
rect 27712 24686 27764 24692
rect 27436 24608 27488 24614
rect 27436 24550 27488 24556
rect 27344 24268 27396 24274
rect 27344 24210 27396 24216
rect 27356 24018 27384 24210
rect 27448 24138 27476 24550
rect 27620 24336 27672 24342
rect 27620 24278 27672 24284
rect 27436 24132 27488 24138
rect 27436 24074 27488 24080
rect 27528 24132 27580 24138
rect 27528 24074 27580 24080
rect 27540 24018 27568 24074
rect 27172 23990 27384 24018
rect 27448 23990 27568 24018
rect 27172 23730 27200 23990
rect 27448 23730 27476 23990
rect 27632 23730 27660 24278
rect 27160 23724 27212 23730
rect 27160 23666 27212 23672
rect 27436 23724 27488 23730
rect 27436 23666 27488 23672
rect 27620 23724 27672 23730
rect 27620 23666 27672 23672
rect 27172 23186 27200 23666
rect 27448 23594 27476 23666
rect 27436 23588 27488 23594
rect 27436 23530 27488 23536
rect 27160 23180 27212 23186
rect 27160 23122 27212 23128
rect 27172 22982 27200 23122
rect 27252 23112 27304 23118
rect 27252 23054 27304 23060
rect 27160 22976 27212 22982
rect 27160 22918 27212 22924
rect 26792 22024 26844 22030
rect 26792 21966 26844 21972
rect 26712 21678 26832 21706
rect 26700 21616 26752 21622
rect 26700 21558 26752 21564
rect 26712 21146 26740 21558
rect 26700 21140 26752 21146
rect 26700 21082 26752 21088
rect 26608 17808 26660 17814
rect 26608 17750 26660 17756
rect 26620 17202 26648 17750
rect 26700 17740 26752 17746
rect 26700 17682 26752 17688
rect 26608 17196 26660 17202
rect 26608 17138 26660 17144
rect 26712 16590 26740 17682
rect 26804 16590 26832 21678
rect 27172 21554 27200 22918
rect 27264 22166 27292 23054
rect 27448 23050 27476 23530
rect 27436 23044 27488 23050
rect 27436 22986 27488 22992
rect 27252 22160 27304 22166
rect 27252 22102 27304 22108
rect 27160 21548 27212 21554
rect 27160 21490 27212 21496
rect 26976 20460 27028 20466
rect 26976 20402 27028 20408
rect 26988 18426 27016 20402
rect 27068 18624 27120 18630
rect 27068 18566 27120 18572
rect 26976 18420 27028 18426
rect 26976 18362 27028 18368
rect 27080 18358 27108 18566
rect 27068 18352 27120 18358
rect 27068 18294 27120 18300
rect 27172 17338 27200 21490
rect 27264 21010 27292 22102
rect 27344 21684 27396 21690
rect 27344 21626 27396 21632
rect 27356 21078 27384 21626
rect 27448 21554 27476 22986
rect 27436 21548 27488 21554
rect 27436 21490 27488 21496
rect 27528 21412 27580 21418
rect 27528 21354 27580 21360
rect 27344 21072 27396 21078
rect 27344 21014 27396 21020
rect 27252 21004 27304 21010
rect 27252 20946 27304 20952
rect 27540 20942 27568 21354
rect 27528 20936 27580 20942
rect 27528 20878 27580 20884
rect 27436 20868 27488 20874
rect 27436 20810 27488 20816
rect 27252 20800 27304 20806
rect 27252 20742 27304 20748
rect 27264 20602 27292 20742
rect 27252 20596 27304 20602
rect 27252 20538 27304 20544
rect 27448 20074 27476 20810
rect 27632 20602 27660 23666
rect 27724 22522 27752 24686
rect 27816 24070 27844 25094
rect 27894 25050 27950 26086
rect 27894 24998 27896 25050
rect 27948 24998 27950 25050
rect 27804 24064 27856 24070
rect 27804 24006 27856 24012
rect 27816 23186 27844 24006
rect 27894 23962 27950 24998
rect 27894 23910 27896 23962
rect 27948 23910 27950 23962
rect 27804 23180 27856 23186
rect 27804 23122 27856 23128
rect 27816 22642 27844 23122
rect 27894 22874 27950 23910
rect 28000 23322 28028 26930
rect 28080 26784 28132 26790
rect 28080 26726 28132 26732
rect 27988 23316 28040 23322
rect 27988 23258 28040 23264
rect 27894 22822 27896 22874
rect 27948 22822 27950 22874
rect 27804 22636 27856 22642
rect 27804 22578 27856 22584
rect 27724 22494 27844 22522
rect 27712 22092 27764 22098
rect 27712 22034 27764 22040
rect 27724 21622 27752 22034
rect 27712 21616 27764 21622
rect 27712 21558 27764 21564
rect 27816 21554 27844 22494
rect 27894 21786 27950 22822
rect 28092 22710 28120 26726
rect 28184 24936 28212 28086
rect 28276 25294 28304 30262
rect 28356 29164 28408 29170
rect 28356 29106 28408 29112
rect 28264 25288 28316 25294
rect 28264 25230 28316 25236
rect 28184 24908 28304 24936
rect 28172 24812 28224 24818
rect 28172 24754 28224 24760
rect 28184 23662 28212 24754
rect 28276 23730 28304 24908
rect 28368 23866 28396 29106
rect 28460 28218 28488 32506
rect 28552 32026 28580 33458
rect 28644 33114 28672 36110
rect 29012 35562 29040 36790
rect 29288 36786 29316 37080
rect 29276 36780 29328 36786
rect 29276 36722 29328 36728
rect 29276 35692 29328 35698
rect 29276 35634 29328 35640
rect 29000 35556 29052 35562
rect 29000 35498 29052 35504
rect 28724 35148 28776 35154
rect 28724 35090 28776 35096
rect 28736 33998 28764 35090
rect 29012 35086 29040 35498
rect 29184 35284 29236 35290
rect 29184 35226 29236 35232
rect 29000 35080 29052 35086
rect 29000 35022 29052 35028
rect 28908 34672 28960 34678
rect 28908 34614 28960 34620
rect 28920 34134 28948 34614
rect 29012 34202 29040 35022
rect 29000 34196 29052 34202
rect 29000 34138 29052 34144
rect 28908 34128 28960 34134
rect 28908 34070 28960 34076
rect 28724 33992 28776 33998
rect 28724 33934 28776 33940
rect 28724 33856 28776 33862
rect 28724 33798 28776 33804
rect 28632 33108 28684 33114
rect 28632 33050 28684 33056
rect 28632 32904 28684 32910
rect 28632 32846 28684 32852
rect 28540 32020 28592 32026
rect 28540 31962 28592 31968
rect 28644 31346 28672 32846
rect 28736 31822 28764 33798
rect 28920 33046 28948 34070
rect 29012 33590 29040 34138
rect 29092 33652 29144 33658
rect 29092 33594 29144 33600
rect 29000 33584 29052 33590
rect 29000 33526 29052 33532
rect 29104 33114 29132 33594
rect 29092 33108 29144 33114
rect 29092 33050 29144 33056
rect 28908 33040 28960 33046
rect 28908 32982 28960 32988
rect 28920 32774 28948 32982
rect 28908 32768 28960 32774
rect 28908 32710 28960 32716
rect 28920 32042 28948 32710
rect 29092 32224 29144 32230
rect 29092 32166 29144 32172
rect 28828 32014 28948 32042
rect 28828 31822 28856 32014
rect 28908 31952 28960 31958
rect 28908 31894 28960 31900
rect 28724 31816 28776 31822
rect 28724 31758 28776 31764
rect 28816 31816 28868 31822
rect 28816 31758 28868 31764
rect 28632 31340 28684 31346
rect 28632 31282 28684 31288
rect 28920 30734 28948 31894
rect 28908 30728 28960 30734
rect 28908 30670 28960 30676
rect 29000 30728 29052 30734
rect 29000 30670 29052 30676
rect 28724 30116 28776 30122
rect 28724 30058 28776 30064
rect 28736 29646 28764 30058
rect 28920 29646 28948 30670
rect 28724 29640 28776 29646
rect 28724 29582 28776 29588
rect 28908 29640 28960 29646
rect 28908 29582 28960 29588
rect 28540 28484 28592 28490
rect 28540 28426 28592 28432
rect 28448 28212 28500 28218
rect 28448 28154 28500 28160
rect 28448 28008 28500 28014
rect 28448 27950 28500 27956
rect 28460 27334 28488 27950
rect 28552 27674 28580 28426
rect 28632 27872 28684 27878
rect 28632 27814 28684 27820
rect 28724 27872 28776 27878
rect 28724 27814 28776 27820
rect 28644 27674 28672 27814
rect 28540 27668 28592 27674
rect 28540 27610 28592 27616
rect 28632 27668 28684 27674
rect 28632 27610 28684 27616
rect 28736 27470 28764 27814
rect 28920 27470 28948 29582
rect 29012 28762 29040 30670
rect 29000 28756 29052 28762
rect 29000 28698 29052 28704
rect 29104 28694 29132 32166
rect 29196 31890 29224 35226
rect 29288 35222 29316 35634
rect 29276 35216 29328 35222
rect 29276 35158 29328 35164
rect 29288 34610 29316 35158
rect 29276 34604 29328 34610
rect 29276 34546 29328 34552
rect 29288 34066 29316 34546
rect 29276 34060 29328 34066
rect 29276 34002 29328 34008
rect 29276 33584 29328 33590
rect 29276 33526 29328 33532
rect 29288 32978 29316 33526
rect 29276 32972 29328 32978
rect 29276 32914 29328 32920
rect 29184 31884 29236 31890
rect 29184 31826 29236 31832
rect 29276 29640 29328 29646
rect 29276 29582 29328 29588
rect 29288 29170 29316 29582
rect 29276 29164 29328 29170
rect 29276 29106 29328 29112
rect 29184 29096 29236 29102
rect 29184 29038 29236 29044
rect 29092 28688 29144 28694
rect 29092 28630 29144 28636
rect 29196 28422 29224 29038
rect 29184 28416 29236 28422
rect 29184 28358 29236 28364
rect 29196 27538 29224 28358
rect 29276 27940 29328 27946
rect 29276 27882 29328 27888
rect 29184 27532 29236 27538
rect 29184 27474 29236 27480
rect 28724 27464 28776 27470
rect 28724 27406 28776 27412
rect 28908 27464 28960 27470
rect 28908 27406 28960 27412
rect 28448 27328 28500 27334
rect 28448 27270 28500 27276
rect 28540 26920 28592 26926
rect 28540 26862 28592 26868
rect 28448 26784 28500 26790
rect 28448 26726 28500 26732
rect 28460 24614 28488 26726
rect 28448 24608 28500 24614
rect 28448 24550 28500 24556
rect 28356 23860 28408 23866
rect 28356 23802 28408 23808
rect 28264 23724 28316 23730
rect 28264 23666 28316 23672
rect 28172 23656 28224 23662
rect 28172 23598 28224 23604
rect 28080 22704 28132 22710
rect 28080 22646 28132 22652
rect 28460 22098 28488 24550
rect 28552 24342 28580 26862
rect 28920 26858 28948 27406
rect 29184 26988 29236 26994
rect 29184 26930 29236 26936
rect 28908 26852 28960 26858
rect 28908 26794 28960 26800
rect 28632 26784 28684 26790
rect 28632 26726 28684 26732
rect 28644 25906 28672 26726
rect 29000 26444 29052 26450
rect 29000 26386 29052 26392
rect 28632 25900 28684 25906
rect 28632 25842 28684 25848
rect 29012 25702 29040 26386
rect 29092 26376 29144 26382
rect 29092 26318 29144 26324
rect 29000 25696 29052 25702
rect 29000 25638 29052 25644
rect 28540 24336 28592 24342
rect 28540 24278 28592 24284
rect 29012 24206 29040 25638
rect 29104 24818 29132 26318
rect 29092 24812 29144 24818
rect 29092 24754 29144 24760
rect 29196 24410 29224 26930
rect 29184 24404 29236 24410
rect 29184 24346 29236 24352
rect 28724 24200 28776 24206
rect 28724 24142 28776 24148
rect 29000 24200 29052 24206
rect 29000 24142 29052 24148
rect 28448 22092 28500 22098
rect 28448 22034 28500 22040
rect 27894 21734 27896 21786
rect 27948 21734 27950 21786
rect 27804 21548 27856 21554
rect 27804 21490 27856 21496
rect 27712 21480 27764 21486
rect 27712 21422 27764 21428
rect 27724 20942 27752 21422
rect 27712 20936 27764 20942
rect 27712 20878 27764 20884
rect 27816 20602 27844 21490
rect 27894 20698 27950 21734
rect 28264 21548 28316 21554
rect 28264 21490 28316 21496
rect 27988 21344 28040 21350
rect 27988 21286 28040 21292
rect 28172 21344 28224 21350
rect 28172 21286 28224 21292
rect 27894 20646 27896 20698
rect 27948 20646 27950 20698
rect 27620 20596 27672 20602
rect 27620 20538 27672 20544
rect 27804 20596 27856 20602
rect 27804 20538 27856 20544
rect 27712 20392 27764 20398
rect 27712 20334 27764 20340
rect 27620 20324 27672 20330
rect 27620 20266 27672 20272
rect 27448 20046 27568 20074
rect 27540 19990 27568 20046
rect 27436 19984 27488 19990
rect 27436 19926 27488 19932
rect 27528 19984 27580 19990
rect 27528 19926 27580 19932
rect 27344 19304 27396 19310
rect 27344 19246 27396 19252
rect 27252 19168 27304 19174
rect 27252 19110 27304 19116
rect 27160 17332 27212 17338
rect 27160 17274 27212 17280
rect 27264 17270 27292 19110
rect 27356 18902 27384 19246
rect 27344 18896 27396 18902
rect 27344 18838 27396 18844
rect 27344 18284 27396 18290
rect 27344 18226 27396 18232
rect 27356 17882 27384 18226
rect 27448 17882 27476 19926
rect 27632 19922 27660 20266
rect 27724 19938 27752 20334
rect 27816 20058 27844 20538
rect 27804 20052 27856 20058
rect 27804 19994 27856 20000
rect 27620 19916 27672 19922
rect 27724 19910 27844 19938
rect 27620 19858 27672 19864
rect 27632 19768 27660 19858
rect 27816 19786 27844 19910
rect 27804 19780 27856 19786
rect 27632 19740 27752 19768
rect 27528 18624 27580 18630
rect 27528 18566 27580 18572
rect 27540 18290 27568 18566
rect 27724 18426 27752 19740
rect 27804 19722 27856 19728
rect 27712 18420 27764 18426
rect 27712 18362 27764 18368
rect 27528 18284 27580 18290
rect 27528 18226 27580 18232
rect 27344 17876 27396 17882
rect 27344 17818 27396 17824
rect 27436 17876 27488 17882
rect 27436 17818 27488 17824
rect 27252 17264 27304 17270
rect 27252 17206 27304 17212
rect 26700 16584 26752 16590
rect 26700 16526 26752 16532
rect 26792 16584 26844 16590
rect 26792 16526 26844 16532
rect 27252 16584 27304 16590
rect 27252 16526 27304 16532
rect 26804 14958 26832 16526
rect 26976 16108 27028 16114
rect 26976 16050 27028 16056
rect 26884 15428 26936 15434
rect 26884 15370 26936 15376
rect 26792 14952 26844 14958
rect 26792 14894 26844 14900
rect 26896 13802 26924 15370
rect 26988 15366 27016 16050
rect 27264 16046 27292 16526
rect 27252 16040 27304 16046
rect 27252 15982 27304 15988
rect 27264 15434 27292 15982
rect 27448 15910 27476 17818
rect 27540 16046 27568 18226
rect 27816 18086 27844 19722
rect 27894 19610 27950 20646
rect 27894 19558 27896 19610
rect 27948 19558 27950 19610
rect 27894 18522 27950 19558
rect 28000 18698 28028 21286
rect 28184 21078 28212 21286
rect 28080 21072 28132 21078
rect 28080 21014 28132 21020
rect 28172 21072 28224 21078
rect 28172 21014 28224 21020
rect 28092 20856 28120 21014
rect 28172 20868 28224 20874
rect 28092 20828 28172 20856
rect 28172 20810 28224 20816
rect 28276 20058 28304 21490
rect 28540 21480 28592 21486
rect 28540 21422 28592 21428
rect 28552 21146 28580 21422
rect 28632 21412 28684 21418
rect 28632 21354 28684 21360
rect 28540 21140 28592 21146
rect 28540 21082 28592 21088
rect 28540 21004 28592 21010
rect 28540 20946 28592 20952
rect 28448 20936 28500 20942
rect 28448 20878 28500 20884
rect 28460 20330 28488 20878
rect 28448 20324 28500 20330
rect 28448 20266 28500 20272
rect 28264 20052 28316 20058
rect 28264 19994 28316 20000
rect 28356 19780 28408 19786
rect 28356 19722 28408 19728
rect 28172 19712 28224 19718
rect 28172 19654 28224 19660
rect 28080 19168 28132 19174
rect 28080 19110 28132 19116
rect 28092 18766 28120 19110
rect 28080 18760 28132 18766
rect 28080 18702 28132 18708
rect 27988 18692 28040 18698
rect 27988 18634 28040 18640
rect 27894 18470 27896 18522
rect 27948 18470 27950 18522
rect 27804 18080 27856 18086
rect 27804 18022 27856 18028
rect 27804 17604 27856 17610
rect 27804 17546 27856 17552
rect 27620 17536 27672 17542
rect 27620 17478 27672 17484
rect 27632 17202 27660 17478
rect 27620 17196 27672 17202
rect 27620 17138 27672 17144
rect 27528 16040 27580 16046
rect 27528 15982 27580 15988
rect 27436 15904 27488 15910
rect 27436 15846 27488 15852
rect 27252 15428 27304 15434
rect 27252 15370 27304 15376
rect 26976 15360 27028 15366
rect 26976 15302 27028 15308
rect 26988 15026 27016 15302
rect 27448 15162 27476 15846
rect 27436 15156 27488 15162
rect 27436 15098 27488 15104
rect 26976 15020 27028 15026
rect 26976 14962 27028 14968
rect 27252 15020 27304 15026
rect 27252 14962 27304 14968
rect 26988 13818 27016 14962
rect 27068 14816 27120 14822
rect 27068 14758 27120 14764
rect 27160 14816 27212 14822
rect 27160 14758 27212 14764
rect 27080 13938 27108 14758
rect 27172 14414 27200 14758
rect 27264 14414 27292 14962
rect 27344 14952 27396 14958
rect 27344 14894 27396 14900
rect 27160 14408 27212 14414
rect 27160 14350 27212 14356
rect 27252 14408 27304 14414
rect 27252 14350 27304 14356
rect 27068 13932 27120 13938
rect 27068 13874 27120 13880
rect 26884 13796 26936 13802
rect 26988 13790 27108 13818
rect 26884 13738 26936 13744
rect 26516 13524 26568 13530
rect 26516 13466 26568 13472
rect 26332 13184 26384 13190
rect 26332 13126 26384 13132
rect 26528 12442 26556 13466
rect 27080 13394 27108 13790
rect 27160 13796 27212 13802
rect 27160 13738 27212 13744
rect 27172 13530 27200 13738
rect 27160 13524 27212 13530
rect 27160 13466 27212 13472
rect 27068 13388 27120 13394
rect 27068 13330 27120 13336
rect 26792 13320 26844 13326
rect 26792 13262 26844 13268
rect 26804 12986 26832 13262
rect 26976 13184 27028 13190
rect 26976 13126 27028 13132
rect 26792 12980 26844 12986
rect 26792 12922 26844 12928
rect 26516 12436 26568 12442
rect 26516 12378 26568 12384
rect 26988 12238 27016 13126
rect 26700 12232 26752 12238
rect 26700 12174 26752 12180
rect 26976 12232 27028 12238
rect 26976 12174 27028 12180
rect 26712 11150 26740 12174
rect 26792 12096 26844 12102
rect 26792 12038 26844 12044
rect 26804 11150 26832 12038
rect 26700 11144 26752 11150
rect 26700 11086 26752 11092
rect 26792 11144 26844 11150
rect 26792 11086 26844 11092
rect 26240 10668 26292 10674
rect 26292 10628 26464 10656
rect 26240 10610 26292 10616
rect 26252 10538 26280 10610
rect 26240 10532 26292 10538
rect 26240 10474 26292 10480
rect 26332 10464 26384 10470
rect 26332 10406 26384 10412
rect 26148 9988 26200 9994
rect 26148 9930 26200 9936
rect 26160 9178 26188 9930
rect 26240 9920 26292 9926
rect 26240 9862 26292 9868
rect 26252 9722 26280 9862
rect 26240 9716 26292 9722
rect 26240 9658 26292 9664
rect 26148 9172 26200 9178
rect 26148 9114 26200 9120
rect 26344 8974 26372 10406
rect 26436 9722 26464 10628
rect 26712 10010 26740 11086
rect 27264 11082 27292 14350
rect 27356 13530 27384 14894
rect 27448 14618 27476 15098
rect 27436 14612 27488 14618
rect 27436 14554 27488 14560
rect 27540 13938 27568 15982
rect 27620 15564 27672 15570
rect 27620 15506 27672 15512
rect 27632 14618 27660 15506
rect 27712 15496 27764 15502
rect 27712 15438 27764 15444
rect 27724 15162 27752 15438
rect 27712 15156 27764 15162
rect 27712 15098 27764 15104
rect 27620 14612 27672 14618
rect 27620 14554 27672 14560
rect 27528 13932 27580 13938
rect 27528 13874 27580 13880
rect 27816 13870 27844 17546
rect 27894 17434 27950 18470
rect 28184 18222 28212 19654
rect 28368 19514 28396 19722
rect 28552 19514 28580 20946
rect 28356 19508 28408 19514
rect 28356 19450 28408 19456
rect 28540 19508 28592 19514
rect 28540 19450 28592 19456
rect 28448 19372 28500 19378
rect 28448 19314 28500 19320
rect 28460 18426 28488 19314
rect 28644 19310 28672 21354
rect 28736 19854 28764 24142
rect 28908 23724 28960 23730
rect 28908 23666 28960 23672
rect 28920 22710 28948 23666
rect 29184 23248 29236 23254
rect 29184 23190 29236 23196
rect 28908 22704 28960 22710
rect 28908 22646 28960 22652
rect 29196 21622 29224 23190
rect 29288 23050 29316 27882
rect 29380 27334 29408 42026
rect 29736 41608 29788 41614
rect 29736 41550 29788 41556
rect 29828 41608 29880 41614
rect 29828 41550 29880 41556
rect 29644 41472 29696 41478
rect 29644 41414 29696 41420
rect 29552 40588 29604 40594
rect 29552 40530 29604 40536
rect 29460 39976 29512 39982
rect 29460 39918 29512 39924
rect 29472 38350 29500 39918
rect 29564 39506 29592 40530
rect 29656 40526 29684 41414
rect 29644 40520 29696 40526
rect 29644 40462 29696 40468
rect 29644 40044 29696 40050
rect 29644 39986 29696 39992
rect 29656 39914 29684 39986
rect 29644 39908 29696 39914
rect 29644 39850 29696 39856
rect 29552 39500 29604 39506
rect 29552 39442 29604 39448
rect 29460 38344 29512 38350
rect 29460 38286 29512 38292
rect 29564 37942 29592 39442
rect 29656 38894 29684 39850
rect 29644 38888 29696 38894
rect 29644 38830 29696 38836
rect 29748 38554 29776 41550
rect 29840 40050 29868 41550
rect 29920 41064 29972 41070
rect 29920 41006 29972 41012
rect 29932 40730 29960 41006
rect 29920 40724 29972 40730
rect 29920 40666 29972 40672
rect 29828 40044 29880 40050
rect 29828 39986 29880 39992
rect 29736 38548 29788 38554
rect 29736 38490 29788 38496
rect 29736 38344 29788 38350
rect 29736 38286 29788 38292
rect 29552 37936 29604 37942
rect 29552 37878 29604 37884
rect 29552 37800 29604 37806
rect 29552 37742 29604 37748
rect 29644 37800 29696 37806
rect 29644 37742 29696 37748
rect 29564 36582 29592 37742
rect 29656 37126 29684 37742
rect 29748 37398 29776 38286
rect 29840 38282 29868 39986
rect 30012 38888 30064 38894
rect 30012 38830 30064 38836
rect 30024 38350 30052 38830
rect 30012 38344 30064 38350
rect 30012 38286 30064 38292
rect 29828 38276 29880 38282
rect 29828 38218 29880 38224
rect 29828 37460 29880 37466
rect 29828 37402 29880 37408
rect 29736 37392 29788 37398
rect 29736 37334 29788 37340
rect 29644 37120 29696 37126
rect 29644 37062 29696 37068
rect 29552 36576 29604 36582
rect 29552 36518 29604 36524
rect 29552 36236 29604 36242
rect 29656 36224 29684 37062
rect 29748 36786 29776 37334
rect 29736 36780 29788 36786
rect 29736 36722 29788 36728
rect 29604 36196 29684 36224
rect 29552 36178 29604 36184
rect 29460 35692 29512 35698
rect 29460 35634 29512 35640
rect 29472 35290 29500 35634
rect 29564 35562 29592 36178
rect 29736 35624 29788 35630
rect 29736 35566 29788 35572
rect 29552 35556 29604 35562
rect 29552 35498 29604 35504
rect 29460 35284 29512 35290
rect 29460 35226 29512 35232
rect 29748 34610 29776 35566
rect 29736 34604 29788 34610
rect 29736 34546 29788 34552
rect 29552 34536 29604 34542
rect 29552 34478 29604 34484
rect 29460 33992 29512 33998
rect 29460 33934 29512 33940
rect 29472 33454 29500 33934
rect 29460 33448 29512 33454
rect 29460 33390 29512 33396
rect 29472 32434 29500 33390
rect 29564 32842 29592 34478
rect 29748 33998 29776 34546
rect 29840 34474 29868 37402
rect 30024 36854 30052 38286
rect 30116 37194 30144 42502
rect 31392 42220 31444 42226
rect 31392 42162 31444 42168
rect 31024 41676 31076 41682
rect 31024 41618 31076 41624
rect 30288 41472 30340 41478
rect 30288 41414 30340 41420
rect 30300 40730 30328 41414
rect 30472 40928 30524 40934
rect 30472 40870 30524 40876
rect 30288 40724 30340 40730
rect 30288 40666 30340 40672
rect 30484 40050 30512 40870
rect 30932 40384 30984 40390
rect 30932 40326 30984 40332
rect 30656 40112 30708 40118
rect 30656 40054 30708 40060
rect 30472 40044 30524 40050
rect 30472 39986 30524 39992
rect 30472 39364 30524 39370
rect 30472 39306 30524 39312
rect 30484 39098 30512 39306
rect 30472 39092 30524 39098
rect 30472 39034 30524 39040
rect 30668 38962 30696 40054
rect 30656 38956 30708 38962
rect 30656 38898 30708 38904
rect 30944 38894 30972 40326
rect 31036 38962 31064 41618
rect 31300 41608 31352 41614
rect 31300 41550 31352 41556
rect 31116 41472 31168 41478
rect 31116 41414 31168 41420
rect 31024 38956 31076 38962
rect 31024 38898 31076 38904
rect 30932 38888 30984 38894
rect 30932 38830 30984 38836
rect 30944 38418 30972 38830
rect 31036 38554 31064 38898
rect 31024 38548 31076 38554
rect 31024 38490 31076 38496
rect 30932 38412 30984 38418
rect 30932 38354 30984 38360
rect 30288 38344 30340 38350
rect 30288 38286 30340 38292
rect 30104 37188 30156 37194
rect 30104 37130 30156 37136
rect 30300 36922 30328 38286
rect 30656 38208 30708 38214
rect 30656 38150 30708 38156
rect 30668 37942 30696 38150
rect 30656 37936 30708 37942
rect 30656 37878 30708 37884
rect 30288 36916 30340 36922
rect 30288 36858 30340 36864
rect 30012 36848 30064 36854
rect 30012 36790 30064 36796
rect 31036 36650 31064 38490
rect 31128 38010 31156 41414
rect 31312 41206 31340 41550
rect 31404 41546 31432 42162
rect 31484 42152 31536 42158
rect 31484 42094 31536 42100
rect 31392 41540 31444 41546
rect 31392 41482 31444 41488
rect 31300 41200 31352 41206
rect 31300 41142 31352 41148
rect 31300 40044 31352 40050
rect 31300 39986 31352 39992
rect 31312 39302 31340 39986
rect 31300 39296 31352 39302
rect 31300 39238 31352 39244
rect 31312 39030 31340 39238
rect 31300 39024 31352 39030
rect 31300 38966 31352 38972
rect 31312 38418 31340 38966
rect 31300 38412 31352 38418
rect 31300 38354 31352 38360
rect 31116 38004 31168 38010
rect 31116 37946 31168 37952
rect 31300 37664 31352 37670
rect 31300 37606 31352 37612
rect 31312 36786 31340 37606
rect 31300 36780 31352 36786
rect 31300 36722 31352 36728
rect 31024 36644 31076 36650
rect 31024 36586 31076 36592
rect 30840 36032 30892 36038
rect 30840 35974 30892 35980
rect 30196 35080 30248 35086
rect 30196 35022 30248 35028
rect 30208 34610 30236 35022
rect 30852 34746 30880 35974
rect 31300 35488 31352 35494
rect 31300 35430 31352 35436
rect 31312 35086 31340 35430
rect 30932 35080 30984 35086
rect 30932 35022 30984 35028
rect 31300 35080 31352 35086
rect 31300 35022 31352 35028
rect 30380 34740 30432 34746
rect 30380 34682 30432 34688
rect 30840 34740 30892 34746
rect 30840 34682 30892 34688
rect 30196 34604 30248 34610
rect 30196 34546 30248 34552
rect 29828 34468 29880 34474
rect 29828 34410 29880 34416
rect 30024 34054 30236 34082
rect 29736 33992 29788 33998
rect 29736 33934 29788 33940
rect 29748 33522 29776 33934
rect 30024 33658 30052 34054
rect 30208 33998 30236 34054
rect 30104 33992 30156 33998
rect 30104 33934 30156 33940
rect 30196 33992 30248 33998
rect 30196 33934 30248 33940
rect 30012 33652 30064 33658
rect 30012 33594 30064 33600
rect 30116 33590 30144 33934
rect 30196 33856 30248 33862
rect 30196 33798 30248 33804
rect 30104 33584 30156 33590
rect 30104 33526 30156 33532
rect 29736 33516 29788 33522
rect 29736 33458 29788 33464
rect 29552 32836 29604 32842
rect 29552 32778 29604 32784
rect 29644 32768 29696 32774
rect 29644 32710 29696 32716
rect 29460 32428 29512 32434
rect 29460 32370 29512 32376
rect 29656 32366 29684 32710
rect 29644 32360 29696 32366
rect 29644 32302 29696 32308
rect 29748 32026 29776 33458
rect 30208 32910 30236 33798
rect 30196 32904 30248 32910
rect 30196 32846 30248 32852
rect 30392 32366 30420 34682
rect 30748 34468 30800 34474
rect 30748 34410 30800 34416
rect 30472 32836 30524 32842
rect 30472 32778 30524 32784
rect 30484 32366 30512 32778
rect 30380 32360 30432 32366
rect 30380 32302 30432 32308
rect 30472 32360 30524 32366
rect 30472 32302 30524 32308
rect 30656 32360 30708 32366
rect 30656 32302 30708 32308
rect 29828 32292 29880 32298
rect 29828 32234 29880 32240
rect 29736 32020 29788 32026
rect 29736 31962 29788 31968
rect 29840 30190 29868 32234
rect 30668 32230 30696 32302
rect 30380 32224 30432 32230
rect 30380 32166 30432 32172
rect 30656 32224 30708 32230
rect 30656 32166 30708 32172
rect 30104 31884 30156 31890
rect 30104 31826 30156 31832
rect 29920 31272 29972 31278
rect 29920 31214 29972 31220
rect 29828 30184 29880 30190
rect 29828 30126 29880 30132
rect 29736 29572 29788 29578
rect 29736 29514 29788 29520
rect 29748 28966 29776 29514
rect 29840 29034 29868 30126
rect 29932 30054 29960 31214
rect 30116 30734 30144 31826
rect 30288 31816 30340 31822
rect 30288 31758 30340 31764
rect 30196 31680 30248 31686
rect 30196 31622 30248 31628
rect 30208 31346 30236 31622
rect 30196 31340 30248 31346
rect 30196 31282 30248 31288
rect 30300 30938 30328 31758
rect 30288 30932 30340 30938
rect 30288 30874 30340 30880
rect 30104 30728 30156 30734
rect 30104 30670 30156 30676
rect 30012 30592 30064 30598
rect 30012 30534 30064 30540
rect 29920 30048 29972 30054
rect 29920 29990 29972 29996
rect 29932 29714 29960 29990
rect 29920 29708 29972 29714
rect 29920 29650 29972 29656
rect 30024 29646 30052 30534
rect 30116 29850 30144 30670
rect 30104 29844 30156 29850
rect 30104 29786 30156 29792
rect 30012 29640 30064 29646
rect 30012 29582 30064 29588
rect 30012 29504 30064 29510
rect 30012 29446 30064 29452
rect 29828 29028 29880 29034
rect 29828 28970 29880 28976
rect 29736 28960 29788 28966
rect 29736 28902 29788 28908
rect 29736 28756 29788 28762
rect 29736 28698 29788 28704
rect 29748 28082 29776 28698
rect 30024 28558 30052 29446
rect 30116 29170 30144 29786
rect 30392 29578 30420 32166
rect 30760 31822 30788 34410
rect 30840 33992 30892 33998
rect 30840 33934 30892 33940
rect 30852 33658 30880 33934
rect 30840 33652 30892 33658
rect 30840 33594 30892 33600
rect 30944 32842 30972 35022
rect 31116 33992 31168 33998
rect 31116 33934 31168 33940
rect 30932 32836 30984 32842
rect 30932 32778 30984 32784
rect 31128 32774 31156 33934
rect 31300 33448 31352 33454
rect 31300 33390 31352 33396
rect 31312 33114 31340 33390
rect 31300 33108 31352 33114
rect 31300 33050 31352 33056
rect 31116 32768 31168 32774
rect 31116 32710 31168 32716
rect 30748 31816 30800 31822
rect 30748 31758 30800 31764
rect 31128 31482 31156 32710
rect 31208 31680 31260 31686
rect 31208 31622 31260 31628
rect 31116 31476 31168 31482
rect 31116 31418 31168 31424
rect 30656 31136 30708 31142
rect 30656 31078 30708 31084
rect 30668 30666 30696 31078
rect 31220 30802 31248 31622
rect 31300 31476 31352 31482
rect 31300 31418 31352 31424
rect 30748 30796 30800 30802
rect 30748 30738 30800 30744
rect 31208 30796 31260 30802
rect 31208 30738 31260 30744
rect 30656 30660 30708 30666
rect 30656 30602 30708 30608
rect 30668 30258 30696 30602
rect 30760 30258 30788 30738
rect 31312 30734 31340 31418
rect 31300 30728 31352 30734
rect 31300 30670 31352 30676
rect 30656 30252 30708 30258
rect 30656 30194 30708 30200
rect 30748 30252 30800 30258
rect 30748 30194 30800 30200
rect 31116 30252 31168 30258
rect 31116 30194 31168 30200
rect 30380 29572 30432 29578
rect 30380 29514 30432 29520
rect 30392 29170 30420 29514
rect 30104 29164 30156 29170
rect 30104 29106 30156 29112
rect 30380 29164 30432 29170
rect 30380 29106 30432 29112
rect 30196 29096 30248 29102
rect 30196 29038 30248 29044
rect 30208 28762 30236 29038
rect 30196 28756 30248 28762
rect 30196 28698 30248 28704
rect 29920 28552 29972 28558
rect 29920 28494 29972 28500
rect 30012 28552 30064 28558
rect 30012 28494 30064 28500
rect 29736 28076 29788 28082
rect 29736 28018 29788 28024
rect 29828 27668 29880 27674
rect 29828 27610 29880 27616
rect 29368 27328 29420 27334
rect 29368 27270 29420 27276
rect 29460 26920 29512 26926
rect 29460 26862 29512 26868
rect 29472 23118 29500 26862
rect 29736 26512 29788 26518
rect 29736 26454 29788 26460
rect 29748 26246 29776 26454
rect 29736 26240 29788 26246
rect 29736 26182 29788 26188
rect 29748 24818 29776 26182
rect 29736 24812 29788 24818
rect 29736 24754 29788 24760
rect 29460 23112 29512 23118
rect 29460 23054 29512 23060
rect 29276 23044 29328 23050
rect 29276 22986 29328 22992
rect 29472 22778 29500 23054
rect 29460 22772 29512 22778
rect 29460 22714 29512 22720
rect 29276 22024 29328 22030
rect 29276 21966 29328 21972
rect 29184 21616 29236 21622
rect 29184 21558 29236 21564
rect 28908 21344 28960 21350
rect 28908 21286 28960 21292
rect 28816 20256 28868 20262
rect 28816 20198 28868 20204
rect 28724 19848 28776 19854
rect 28724 19790 28776 19796
rect 28828 19802 28856 20198
rect 28920 19990 28948 21286
rect 29196 20602 29224 21558
rect 29092 20596 29144 20602
rect 29092 20538 29144 20544
rect 29184 20596 29236 20602
rect 29184 20538 29236 20544
rect 29104 20330 29132 20538
rect 29092 20324 29144 20330
rect 29092 20266 29144 20272
rect 28908 19984 28960 19990
rect 28908 19926 28960 19932
rect 28908 19848 28960 19854
rect 28828 19796 28908 19802
rect 28828 19790 28960 19796
rect 28828 19774 28948 19790
rect 29196 19446 29224 20538
rect 29184 19440 29236 19446
rect 29184 19382 29236 19388
rect 28632 19304 28684 19310
rect 28632 19246 28684 19252
rect 28908 19236 28960 19242
rect 28908 19178 28960 19184
rect 28920 18902 28948 19178
rect 28908 18896 28960 18902
rect 28908 18838 28960 18844
rect 28540 18760 28592 18766
rect 28540 18702 28592 18708
rect 28448 18420 28500 18426
rect 28448 18362 28500 18368
rect 28552 18222 28580 18702
rect 28632 18692 28684 18698
rect 28632 18634 28684 18640
rect 28172 18216 28224 18222
rect 28172 18158 28224 18164
rect 28540 18216 28592 18222
rect 28540 18158 28592 18164
rect 28644 17814 28672 18634
rect 28816 18624 28868 18630
rect 28816 18566 28868 18572
rect 29000 18624 29052 18630
rect 29000 18566 29052 18572
rect 28632 17808 28684 17814
rect 28632 17750 28684 17756
rect 28264 17536 28316 17542
rect 28264 17478 28316 17484
rect 27894 17382 27896 17434
rect 27948 17382 27950 17434
rect 27894 16346 27950 17382
rect 27894 16294 27896 16346
rect 27948 16294 27950 16346
rect 27894 15258 27950 16294
rect 28276 16250 28304 17478
rect 28356 16584 28408 16590
rect 28356 16526 28408 16532
rect 28264 16244 28316 16250
rect 28264 16186 28316 16192
rect 28264 15428 28316 15434
rect 28264 15370 28316 15376
rect 27894 15206 27896 15258
rect 27948 15206 27950 15258
rect 27894 14170 27950 15206
rect 28276 15094 28304 15370
rect 28264 15088 28316 15094
rect 28264 15030 28316 15036
rect 27894 14118 27896 14170
rect 27948 14118 27950 14170
rect 27804 13864 27856 13870
rect 27804 13806 27856 13812
rect 27344 13524 27396 13530
rect 27344 13466 27396 13472
rect 27356 12714 27384 13466
rect 27712 13388 27764 13394
rect 27712 13330 27764 13336
rect 27620 13184 27672 13190
rect 27620 13126 27672 13132
rect 27632 12850 27660 13126
rect 27724 12918 27752 13330
rect 27712 12912 27764 12918
rect 27712 12854 27764 12860
rect 27436 12844 27488 12850
rect 27436 12786 27488 12792
rect 27620 12844 27672 12850
rect 27620 12786 27672 12792
rect 27344 12708 27396 12714
rect 27344 12650 27396 12656
rect 27252 11076 27304 11082
rect 27252 11018 27304 11024
rect 27264 10742 27292 11018
rect 27252 10736 27304 10742
rect 27252 10678 27304 10684
rect 27264 10266 27292 10678
rect 27448 10674 27476 12786
rect 27632 12170 27660 12786
rect 27724 12442 27752 12854
rect 27712 12436 27764 12442
rect 27712 12378 27764 12384
rect 27816 12322 27844 13806
rect 27724 12294 27844 12322
rect 27894 13082 27950 14118
rect 27894 13030 27896 13082
rect 27948 13030 27950 13082
rect 27620 12164 27672 12170
rect 27620 12106 27672 12112
rect 27724 12050 27752 12294
rect 27632 12022 27752 12050
rect 27436 10668 27488 10674
rect 27436 10610 27488 10616
rect 27528 10600 27580 10606
rect 27528 10542 27580 10548
rect 27252 10260 27304 10266
rect 27252 10202 27304 10208
rect 27540 10062 27568 10542
rect 26792 10056 26844 10062
rect 26712 10004 26792 10010
rect 26712 9998 26844 10004
rect 27528 10056 27580 10062
rect 27528 9998 27580 10004
rect 26712 9982 26832 9998
rect 26712 9722 26740 9982
rect 26424 9716 26476 9722
rect 26424 9658 26476 9664
rect 26700 9716 26752 9722
rect 26700 9658 26752 9664
rect 26332 8968 26384 8974
rect 26332 8910 26384 8916
rect 27344 8832 27396 8838
rect 27344 8774 27396 8780
rect 26056 8560 26108 8566
rect 26056 8502 26108 8508
rect 27356 8430 27384 8774
rect 27344 8424 27396 8430
rect 27344 8366 27396 8372
rect 26608 8356 26660 8362
rect 26608 8298 26660 8304
rect 26148 7812 26200 7818
rect 26148 7754 26200 7760
rect 26160 7546 26188 7754
rect 26148 7540 26200 7546
rect 26148 7482 26200 7488
rect 26056 7404 26108 7410
rect 26056 7346 26108 7352
rect 26424 7404 26476 7410
rect 26424 7346 26476 7352
rect 25964 6996 26016 7002
rect 25964 6938 26016 6944
rect 25976 6322 26004 6938
rect 24860 6316 24912 6322
rect 24860 6258 24912 6264
rect 24952 6316 25004 6322
rect 24952 6258 25004 6264
rect 25596 6316 25648 6322
rect 25596 6258 25648 6264
rect 25780 6316 25832 6322
rect 25964 6316 26016 6322
rect 25832 6276 25912 6304
rect 25780 6258 25832 6264
rect 24872 4690 24900 6258
rect 24964 5030 24992 6258
rect 25412 5704 25464 5710
rect 25412 5646 25464 5652
rect 25424 5030 25452 5646
rect 24952 5024 25004 5030
rect 24952 4966 25004 4972
rect 25412 5024 25464 5030
rect 25412 4966 25464 4972
rect 24860 4684 24912 4690
rect 24860 4626 24912 4632
rect 24872 4214 24900 4626
rect 24860 4208 24912 4214
rect 24860 4150 24912 4156
rect 24860 3392 24912 3398
rect 24860 3334 24912 3340
rect 24688 2746 24808 2774
rect 24584 2372 24636 2378
rect 24584 2314 24636 2320
rect 24676 1964 24728 1970
rect 24676 1906 24728 1912
rect 24688 1562 24716 1906
rect 24676 1556 24728 1562
rect 24676 1498 24728 1504
rect 24780 882 24808 2746
rect 24872 1358 24900 3334
rect 24964 1426 24992 4966
rect 25228 4208 25280 4214
rect 25228 4150 25280 4156
rect 25044 4072 25096 4078
rect 25044 4014 25096 4020
rect 25056 3534 25084 4014
rect 25240 3534 25268 4150
rect 25608 3534 25636 6258
rect 25688 6248 25740 6254
rect 25688 6190 25740 6196
rect 25700 5914 25728 6190
rect 25780 6112 25832 6118
rect 25780 6054 25832 6060
rect 25688 5908 25740 5914
rect 25688 5850 25740 5856
rect 25700 5302 25728 5850
rect 25688 5296 25740 5302
rect 25688 5238 25740 5244
rect 25700 4146 25728 5238
rect 25792 5234 25820 6054
rect 25884 5642 25912 6276
rect 25964 6258 26016 6264
rect 25872 5636 25924 5642
rect 25872 5578 25924 5584
rect 25780 5228 25832 5234
rect 25780 5170 25832 5176
rect 25688 4140 25740 4146
rect 25688 4082 25740 4088
rect 26068 3942 26096 7346
rect 26332 5840 26384 5846
rect 26332 5782 26384 5788
rect 26148 5636 26200 5642
rect 26148 5578 26200 5584
rect 26056 3936 26108 3942
rect 26056 3878 26108 3884
rect 26160 3534 26188 5578
rect 26240 4752 26292 4758
rect 26240 4694 26292 4700
rect 26252 3738 26280 4694
rect 26344 4078 26372 5782
rect 26436 5098 26464 7346
rect 26516 6316 26568 6322
rect 26516 6258 26568 6264
rect 26424 5092 26476 5098
rect 26424 5034 26476 5040
rect 26424 4140 26476 4146
rect 26424 4082 26476 4088
rect 26332 4072 26384 4078
rect 26332 4014 26384 4020
rect 26240 3732 26292 3738
rect 26240 3674 26292 3680
rect 25044 3528 25096 3534
rect 25044 3470 25096 3476
rect 25228 3528 25280 3534
rect 25228 3470 25280 3476
rect 25596 3528 25648 3534
rect 25596 3470 25648 3476
rect 26148 3528 26200 3534
rect 26148 3470 26200 3476
rect 25056 3058 25084 3470
rect 25240 3126 25268 3470
rect 25228 3120 25280 3126
rect 25228 3062 25280 3068
rect 25044 3052 25096 3058
rect 25044 2994 25096 3000
rect 25240 2650 25268 3062
rect 25320 2848 25372 2854
rect 25320 2790 25372 2796
rect 25228 2644 25280 2650
rect 25228 2586 25280 2592
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 25148 1426 25176 2246
rect 24952 1420 25004 1426
rect 24952 1362 25004 1368
rect 25136 1420 25188 1426
rect 25136 1362 25188 1368
rect 25332 1358 25360 2790
rect 25608 2106 25636 3470
rect 25872 3392 25924 3398
rect 25872 3334 25924 3340
rect 25884 3058 25912 3334
rect 25872 3052 25924 3058
rect 25872 2994 25924 3000
rect 25780 2372 25832 2378
rect 25780 2314 25832 2320
rect 25596 2100 25648 2106
rect 25596 2042 25648 2048
rect 25792 1562 25820 2314
rect 25884 2310 25912 2994
rect 26148 2848 26200 2854
rect 26148 2790 26200 2796
rect 25964 2372 26016 2378
rect 25964 2314 26016 2320
rect 25872 2304 25924 2310
rect 25872 2246 25924 2252
rect 25976 2106 26004 2314
rect 25964 2100 26016 2106
rect 25964 2042 26016 2048
rect 26160 1970 26188 2790
rect 26252 2774 26280 3674
rect 26436 3670 26464 4082
rect 26424 3664 26476 3670
rect 26424 3606 26476 3612
rect 26528 3534 26556 6258
rect 26620 5710 26648 8298
rect 27252 8288 27304 8294
rect 27252 8230 27304 8236
rect 26976 7948 27028 7954
rect 26976 7890 27028 7896
rect 26700 7744 26752 7750
rect 26700 7686 26752 7692
rect 26712 6390 26740 7686
rect 26988 7478 27016 7890
rect 26976 7472 27028 7478
rect 26976 7414 27028 7420
rect 27068 7336 27120 7342
rect 27068 7278 27120 7284
rect 27080 6866 27108 7278
rect 27068 6860 27120 6866
rect 27068 6802 27120 6808
rect 27264 6798 27292 8230
rect 27356 7886 27384 8366
rect 27540 8362 27568 9998
rect 27632 8498 27660 12022
rect 27894 11994 27950 13030
rect 28080 12436 28132 12442
rect 28368 12434 28396 16526
rect 28540 16516 28592 16522
rect 28540 16458 28592 16464
rect 28448 15972 28500 15978
rect 28448 15914 28500 15920
rect 28080 12378 28132 12384
rect 28276 12406 28396 12434
rect 27988 12164 28040 12170
rect 27988 12106 28040 12112
rect 27894 11942 27896 11994
rect 27948 11942 27950 11994
rect 27894 10906 27950 11942
rect 28000 11830 28028 12106
rect 27988 11824 28040 11830
rect 27988 11766 28040 11772
rect 28092 11694 28120 12378
rect 28172 12096 28224 12102
rect 28172 12038 28224 12044
rect 28184 11898 28212 12038
rect 28172 11892 28224 11898
rect 28172 11834 28224 11840
rect 28080 11688 28132 11694
rect 28080 11630 28132 11636
rect 28092 11286 28120 11630
rect 28080 11280 28132 11286
rect 28080 11222 28132 11228
rect 27894 10854 27896 10906
rect 27948 10854 27950 10906
rect 27894 9818 27950 10854
rect 27894 9766 27896 9818
rect 27948 9766 27950 9818
rect 27712 9580 27764 9586
rect 27712 9522 27764 9528
rect 27724 9178 27752 9522
rect 27712 9172 27764 9178
rect 27712 9114 27764 9120
rect 27894 8730 27950 9766
rect 28092 9110 28120 11222
rect 28276 9330 28304 12406
rect 28184 9302 28304 9330
rect 28356 9376 28408 9382
rect 28356 9318 28408 9324
rect 28080 9104 28132 9110
rect 28080 9046 28132 9052
rect 27894 8678 27896 8730
rect 27948 8678 27950 8730
rect 27804 8560 27856 8566
rect 27804 8502 27856 8508
rect 27620 8492 27672 8498
rect 27620 8434 27672 8440
rect 27528 8356 27580 8362
rect 27528 8298 27580 8304
rect 27344 7880 27396 7886
rect 27344 7822 27396 7828
rect 27436 7336 27488 7342
rect 27488 7296 27660 7324
rect 27436 7278 27488 7284
rect 27632 7206 27660 7296
rect 27528 7200 27580 7206
rect 27528 7142 27580 7148
rect 27620 7200 27672 7206
rect 27620 7142 27672 7148
rect 27344 6996 27396 7002
rect 27344 6938 27396 6944
rect 27252 6792 27304 6798
rect 27252 6734 27304 6740
rect 27068 6452 27120 6458
rect 27120 6412 27292 6440
rect 27068 6394 27120 6400
rect 26700 6384 26752 6390
rect 26700 6326 26752 6332
rect 26608 5704 26660 5710
rect 26608 5646 26660 5652
rect 26712 5234 26740 6326
rect 27264 6202 27292 6412
rect 27356 6322 27384 6938
rect 27436 6452 27488 6458
rect 27436 6394 27488 6400
rect 27344 6316 27396 6322
rect 27344 6258 27396 6264
rect 27448 6202 27476 6394
rect 27264 6174 27476 6202
rect 27068 6112 27120 6118
rect 27068 6054 27120 6060
rect 27080 5710 27108 6054
rect 27540 5710 27568 7142
rect 27712 6656 27764 6662
rect 27712 6598 27764 6604
rect 27620 6248 27672 6254
rect 27620 6190 27672 6196
rect 27068 5704 27120 5710
rect 27528 5704 27580 5710
rect 27068 5646 27120 5652
rect 27264 5664 27528 5692
rect 26700 5228 26752 5234
rect 26700 5170 26752 5176
rect 26608 4140 26660 4146
rect 26608 4082 26660 4088
rect 26620 3738 26648 4082
rect 26712 4078 26740 5170
rect 27264 5098 27292 5664
rect 27528 5646 27580 5652
rect 27632 5250 27660 6190
rect 27724 5914 27752 6598
rect 27712 5908 27764 5914
rect 27712 5850 27764 5856
rect 27632 5222 27752 5250
rect 27620 5160 27672 5166
rect 27620 5102 27672 5108
rect 27252 5092 27304 5098
rect 27252 5034 27304 5040
rect 26976 4548 27028 4554
rect 26976 4490 27028 4496
rect 26700 4072 26752 4078
rect 26700 4014 26752 4020
rect 26608 3732 26660 3738
rect 26608 3674 26660 3680
rect 26988 3534 27016 4490
rect 27264 4146 27292 5034
rect 27344 4208 27396 4214
rect 27344 4150 27396 4156
rect 27068 4140 27120 4146
rect 27068 4082 27120 4088
rect 27252 4140 27304 4146
rect 27252 4082 27304 4088
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 26976 3528 27028 3534
rect 26976 3470 27028 3476
rect 26252 2746 26372 2774
rect 26240 2304 26292 2310
rect 26240 2246 26292 2252
rect 26148 1964 26200 1970
rect 26148 1906 26200 1912
rect 25780 1556 25832 1562
rect 25780 1498 25832 1504
rect 26252 1426 26280 2246
rect 26344 1970 26372 2746
rect 27080 2310 27108 4082
rect 27356 2650 27384 4150
rect 27344 2644 27396 2650
rect 27344 2586 27396 2592
rect 27068 2304 27120 2310
rect 27068 2246 27120 2252
rect 27356 1970 27384 2586
rect 27632 2446 27660 5102
rect 27724 3534 27752 5222
rect 27816 4554 27844 8502
rect 27894 7642 27950 8678
rect 27988 8288 28040 8294
rect 27988 8230 28040 8236
rect 27894 7590 27896 7642
rect 27948 7590 27950 7642
rect 27894 6554 27950 7590
rect 28000 7410 28028 8230
rect 28080 7880 28132 7886
rect 28080 7822 28132 7828
rect 28092 7750 28120 7822
rect 28080 7744 28132 7750
rect 28080 7686 28132 7692
rect 27988 7404 28040 7410
rect 27988 7346 28040 7352
rect 28184 7206 28212 9302
rect 28368 9178 28396 9318
rect 28264 9172 28316 9178
rect 28264 9114 28316 9120
rect 28356 9172 28408 9178
rect 28356 9114 28408 9120
rect 28276 8362 28304 9114
rect 28264 8356 28316 8362
rect 28264 8298 28316 8304
rect 28172 7200 28224 7206
rect 28172 7142 28224 7148
rect 28276 6866 28304 8298
rect 28356 7880 28408 7886
rect 28356 7822 28408 7828
rect 28368 7546 28396 7822
rect 28356 7540 28408 7546
rect 28356 7482 28408 7488
rect 28264 6860 28316 6866
rect 28264 6802 28316 6808
rect 27988 6792 28040 6798
rect 27988 6734 28040 6740
rect 27894 6502 27896 6554
rect 27948 6502 27950 6554
rect 27894 5466 27950 6502
rect 28000 6322 28028 6734
rect 27988 6316 28040 6322
rect 27988 6258 28040 6264
rect 27894 5414 27896 5466
rect 27948 5414 27950 5466
rect 27804 4548 27856 4554
rect 27804 4490 27856 4496
rect 27894 4378 27950 5414
rect 28000 4690 28028 6258
rect 28080 5908 28132 5914
rect 28080 5850 28132 5856
rect 28092 5574 28120 5850
rect 28080 5568 28132 5574
rect 28080 5510 28132 5516
rect 27988 4684 28040 4690
rect 27988 4626 28040 4632
rect 28092 4622 28120 5510
rect 28080 4616 28132 4622
rect 28080 4558 28132 4564
rect 27894 4326 27896 4378
rect 27948 4326 27950 4378
rect 27712 3528 27764 3534
rect 27712 3470 27764 3476
rect 27894 3290 27950 4326
rect 27894 3238 27896 3290
rect 27948 3238 27950 3290
rect 27620 2440 27672 2446
rect 27620 2382 27672 2388
rect 27632 2038 27660 2382
rect 27894 2202 27950 3238
rect 28184 4542 28396 4570
rect 27988 3052 28040 3058
rect 27988 2994 28040 3000
rect 28000 2310 28028 2994
rect 27988 2304 28040 2310
rect 27988 2246 28040 2252
rect 28080 2304 28132 2310
rect 28080 2246 28132 2252
rect 27894 2150 27896 2202
rect 27948 2150 27950 2202
rect 27620 2032 27672 2038
rect 27620 1974 27672 1980
rect 26332 1964 26384 1970
rect 26332 1906 26384 1912
rect 27344 1964 27396 1970
rect 27344 1906 27396 1912
rect 27712 1964 27764 1970
rect 27712 1906 27764 1912
rect 26344 1562 26372 1906
rect 27724 1562 27752 1906
rect 26332 1556 26384 1562
rect 26332 1498 26384 1504
rect 27712 1556 27764 1562
rect 27712 1498 27764 1504
rect 26240 1420 26292 1426
rect 26240 1362 26292 1368
rect 24860 1352 24912 1358
rect 24860 1294 24912 1300
rect 25320 1352 25372 1358
rect 25320 1294 25372 1300
rect 26344 1222 26372 1498
rect 27436 1352 27488 1358
rect 27436 1294 27488 1300
rect 26332 1216 26384 1222
rect 26332 1158 26384 1164
rect 24860 944 24912 950
rect 24860 886 24912 892
rect 24768 876 24820 882
rect 24768 818 24820 824
rect 24308 808 24360 814
rect 11980 740 12032 746
rect 11980 682 12032 688
rect 13818 0 13874 800
rect 19338 0 19394 800
rect 24872 800 24900 886
rect 27448 814 27476 1294
rect 27894 1114 27950 2150
rect 28092 1358 28120 2246
rect 28080 1352 28132 1358
rect 28080 1294 28132 1300
rect 28184 1290 28212 4542
rect 28368 4486 28396 4542
rect 28264 4480 28316 4486
rect 28264 4422 28316 4428
rect 28356 4480 28408 4486
rect 28356 4422 28408 4428
rect 28276 4146 28304 4422
rect 28264 4140 28316 4146
rect 28264 4082 28316 4088
rect 28276 3126 28304 4082
rect 28356 3596 28408 3602
rect 28356 3538 28408 3544
rect 28264 3120 28316 3126
rect 28264 3062 28316 3068
rect 28276 2446 28304 3062
rect 28368 2582 28396 3538
rect 28356 2576 28408 2582
rect 28356 2518 28408 2524
rect 28264 2440 28316 2446
rect 28264 2382 28316 2388
rect 28368 1358 28396 2518
rect 28356 1352 28408 1358
rect 28356 1294 28408 1300
rect 28172 1284 28224 1290
rect 28172 1226 28224 1232
rect 27894 1062 27896 1114
rect 27948 1062 27950 1114
rect 27894 1040 27950 1062
rect 27436 808 27488 814
rect 24308 750 24360 756
rect 24858 0 24914 800
rect 27436 750 27488 756
rect 28460 678 28488 15914
rect 28552 12434 28580 16458
rect 28724 15360 28776 15366
rect 28724 15302 28776 15308
rect 28632 15020 28684 15026
rect 28632 14962 28684 14968
rect 28644 14618 28672 14962
rect 28632 14612 28684 14618
rect 28632 14554 28684 14560
rect 28736 14414 28764 15302
rect 28724 14408 28776 14414
rect 28724 14350 28776 14356
rect 28724 14000 28776 14006
rect 28724 13942 28776 13948
rect 28632 13728 28684 13734
rect 28632 13670 28684 13676
rect 28644 13530 28672 13670
rect 28632 13524 28684 13530
rect 28632 13466 28684 13472
rect 28736 13394 28764 13942
rect 28724 13388 28776 13394
rect 28724 13330 28776 13336
rect 28828 13190 28856 18566
rect 29012 18290 29040 18566
rect 29184 18420 29236 18426
rect 29184 18362 29236 18368
rect 29000 18284 29052 18290
rect 29000 18226 29052 18232
rect 29092 18284 29144 18290
rect 29092 18226 29144 18232
rect 29104 17338 29132 18226
rect 29196 18222 29224 18362
rect 29184 18216 29236 18222
rect 29184 18158 29236 18164
rect 29092 17332 29144 17338
rect 29092 17274 29144 17280
rect 29092 17196 29144 17202
rect 29092 17138 29144 17144
rect 29000 16108 29052 16114
rect 29000 16050 29052 16056
rect 28908 15904 28960 15910
rect 28908 15846 28960 15852
rect 28920 15502 28948 15846
rect 29012 15706 29040 16050
rect 29000 15700 29052 15706
rect 29000 15642 29052 15648
rect 28908 15496 28960 15502
rect 28908 15438 28960 15444
rect 29000 15088 29052 15094
rect 29000 15030 29052 15036
rect 28908 13320 28960 13326
rect 28908 13262 28960 13268
rect 28724 13184 28776 13190
rect 28724 13126 28776 13132
rect 28816 13184 28868 13190
rect 28816 13126 28868 13132
rect 28736 12442 28764 13126
rect 28724 12436 28776 12442
rect 28552 12406 28672 12434
rect 28540 9920 28592 9926
rect 28540 9862 28592 9868
rect 28552 8974 28580 9862
rect 28644 9450 28672 12406
rect 28724 12378 28776 12384
rect 28920 11898 28948 13262
rect 29012 12918 29040 15030
rect 29104 14074 29132 17138
rect 29196 16998 29224 18158
rect 29288 17610 29316 21966
rect 29472 21622 29500 22714
rect 29460 21616 29512 21622
rect 29460 21558 29512 21564
rect 29644 20936 29696 20942
rect 29644 20878 29696 20884
rect 29460 20868 29512 20874
rect 29460 20810 29512 20816
rect 29368 20392 29420 20398
rect 29368 20334 29420 20340
rect 29380 19718 29408 20334
rect 29472 20262 29500 20810
rect 29656 20602 29684 20878
rect 29644 20596 29696 20602
rect 29644 20538 29696 20544
rect 29748 20466 29776 24754
rect 29840 22778 29868 27610
rect 29932 27538 29960 28494
rect 30668 28082 30696 30194
rect 30760 28082 30788 30194
rect 30840 28960 30892 28966
rect 31024 28960 31076 28966
rect 30892 28908 30972 28914
rect 30840 28902 30972 28908
rect 31024 28902 31076 28908
rect 30852 28886 30972 28902
rect 30944 28082 30972 28886
rect 31036 28150 31064 28902
rect 31128 28422 31156 30194
rect 31116 28416 31168 28422
rect 31116 28358 31168 28364
rect 31208 28212 31260 28218
rect 31208 28154 31260 28160
rect 31024 28144 31076 28150
rect 31024 28086 31076 28092
rect 30656 28076 30708 28082
rect 30656 28018 30708 28024
rect 30748 28076 30800 28082
rect 30748 28018 30800 28024
rect 30932 28076 30984 28082
rect 30932 28018 30984 28024
rect 30564 27872 30616 27878
rect 30564 27814 30616 27820
rect 29920 27532 29972 27538
rect 29920 27474 29972 27480
rect 30380 27396 30432 27402
rect 30380 27338 30432 27344
rect 30104 27328 30156 27334
rect 30104 27270 30156 27276
rect 29920 26988 29972 26994
rect 29920 26930 29972 26936
rect 29932 26586 29960 26930
rect 29920 26580 29972 26586
rect 29920 26522 29972 26528
rect 30116 26450 30144 27270
rect 30392 27130 30420 27338
rect 30380 27124 30432 27130
rect 30380 27066 30432 27072
rect 30576 26994 30604 27814
rect 30564 26988 30616 26994
rect 30564 26930 30616 26936
rect 31024 26920 31076 26926
rect 31024 26862 31076 26868
rect 30932 26580 30984 26586
rect 30932 26522 30984 26528
rect 30104 26444 30156 26450
rect 30104 26386 30156 26392
rect 30564 26376 30616 26382
rect 30564 26318 30616 26324
rect 30104 26308 30156 26314
rect 30104 26250 30156 26256
rect 30116 25974 30144 26250
rect 30104 25968 30156 25974
rect 30104 25910 30156 25916
rect 30288 25220 30340 25226
rect 30288 25162 30340 25168
rect 30012 24812 30064 24818
rect 30012 24754 30064 24760
rect 30024 24206 30052 24754
rect 30012 24200 30064 24206
rect 30012 24142 30064 24148
rect 29828 22772 29880 22778
rect 29828 22714 29880 22720
rect 30024 22642 30052 24142
rect 30300 23866 30328 25162
rect 30576 24750 30604 26318
rect 30656 24812 30708 24818
rect 30656 24754 30708 24760
rect 30564 24744 30616 24750
rect 30564 24686 30616 24692
rect 30668 24206 30696 24754
rect 30380 24200 30432 24206
rect 30380 24142 30432 24148
rect 30656 24200 30708 24206
rect 30656 24142 30708 24148
rect 30288 23860 30340 23866
rect 30288 23802 30340 23808
rect 30392 23662 30420 24142
rect 30472 24132 30524 24138
rect 30472 24074 30524 24080
rect 30380 23656 30432 23662
rect 30380 23598 30432 23604
rect 30392 22642 30420 23598
rect 30012 22636 30064 22642
rect 30012 22578 30064 22584
rect 30380 22636 30432 22642
rect 30380 22578 30432 22584
rect 29920 22024 29972 22030
rect 29920 21966 29972 21972
rect 29736 20460 29788 20466
rect 29736 20402 29788 20408
rect 29460 20256 29512 20262
rect 29460 20198 29512 20204
rect 29472 20058 29500 20198
rect 29460 20052 29512 20058
rect 29460 19994 29512 20000
rect 29552 20052 29604 20058
rect 29552 19994 29604 20000
rect 29368 19712 29420 19718
rect 29368 19654 29420 19660
rect 29564 19514 29592 19994
rect 29932 19922 29960 21966
rect 30024 21554 30052 22578
rect 30392 21554 30420 22578
rect 30012 21548 30064 21554
rect 30012 21490 30064 21496
rect 30380 21548 30432 21554
rect 30380 21490 30432 21496
rect 29920 19916 29972 19922
rect 29920 19858 29972 19864
rect 29828 19712 29880 19718
rect 29828 19654 29880 19660
rect 29552 19508 29604 19514
rect 29552 19450 29604 19456
rect 29368 19372 29420 19378
rect 29840 19352 29868 19654
rect 29368 19314 29420 19320
rect 29828 19346 29880 19352
rect 29276 17604 29328 17610
rect 29276 17546 29328 17552
rect 29184 16992 29236 16998
rect 29184 16934 29236 16940
rect 29196 14414 29224 16934
rect 29288 16114 29316 17546
rect 29276 16108 29328 16114
rect 29276 16050 29328 16056
rect 29184 14408 29236 14414
rect 29184 14350 29236 14356
rect 29288 14278 29316 16050
rect 29380 15162 29408 19314
rect 29828 19288 29880 19294
rect 29932 17746 29960 19858
rect 30024 18426 30052 21490
rect 30104 21480 30156 21486
rect 30104 21422 30156 21428
rect 30116 20942 30144 21422
rect 30104 20936 30156 20942
rect 30104 20878 30156 20884
rect 30116 19378 30144 20878
rect 30484 20874 30512 24074
rect 30840 24064 30892 24070
rect 30840 24006 30892 24012
rect 30852 23730 30880 24006
rect 30944 23730 30972 26522
rect 30840 23724 30892 23730
rect 30840 23666 30892 23672
rect 30932 23724 30984 23730
rect 30932 23666 30984 23672
rect 30564 22976 30616 22982
rect 30564 22918 30616 22924
rect 30576 22642 30604 22918
rect 30564 22636 30616 22642
rect 30564 22578 30616 22584
rect 30656 22432 30708 22438
rect 30656 22374 30708 22380
rect 30564 21888 30616 21894
rect 30564 21830 30616 21836
rect 30576 21554 30604 21830
rect 30564 21548 30616 21554
rect 30564 21490 30616 21496
rect 30472 20868 30524 20874
rect 30472 20810 30524 20816
rect 30576 20534 30604 21490
rect 30564 20528 30616 20534
rect 30564 20470 30616 20476
rect 30196 20324 30248 20330
rect 30196 20266 30248 20272
rect 30104 19372 30156 19378
rect 30104 19314 30156 19320
rect 30208 18902 30236 20266
rect 30288 20256 30340 20262
rect 30288 20198 30340 20204
rect 30300 19378 30328 20198
rect 30484 20058 30604 20074
rect 30484 20052 30616 20058
rect 30484 20046 30564 20052
rect 30380 19780 30432 19786
rect 30380 19722 30432 19728
rect 30288 19372 30340 19378
rect 30288 19314 30340 19320
rect 30196 18896 30248 18902
rect 30196 18838 30248 18844
rect 30196 18692 30248 18698
rect 30196 18634 30248 18640
rect 30012 18420 30064 18426
rect 30012 18362 30064 18368
rect 30208 18306 30236 18634
rect 30199 18290 30236 18306
rect 30187 18284 30239 18290
rect 30187 18226 30239 18232
rect 29920 17740 29972 17746
rect 29920 17682 29972 17688
rect 29828 17196 29880 17202
rect 29828 17138 29880 17144
rect 29460 16992 29512 16998
rect 29460 16934 29512 16940
rect 29368 15156 29420 15162
rect 29368 15098 29420 15104
rect 29472 14414 29500 16934
rect 29840 15502 29868 17138
rect 29932 16726 29960 17682
rect 30012 17128 30064 17134
rect 30012 17070 30064 17076
rect 29920 16720 29972 16726
rect 29920 16662 29972 16668
rect 29932 16114 29960 16662
rect 29920 16108 29972 16114
rect 29920 16050 29972 16056
rect 29828 15496 29880 15502
rect 29828 15438 29880 15444
rect 29736 14544 29788 14550
rect 29736 14486 29788 14492
rect 29460 14408 29512 14414
rect 29460 14350 29512 14356
rect 29276 14272 29328 14278
rect 29276 14214 29328 14220
rect 29644 14272 29696 14278
rect 29644 14214 29696 14220
rect 29092 14068 29144 14074
rect 29092 14010 29144 14016
rect 29184 13932 29236 13938
rect 29184 13874 29236 13880
rect 29092 13864 29144 13870
rect 29092 13806 29144 13812
rect 29104 13530 29132 13806
rect 29092 13524 29144 13530
rect 29092 13466 29144 13472
rect 29000 12912 29052 12918
rect 29000 12854 29052 12860
rect 29012 12306 29040 12854
rect 29000 12300 29052 12306
rect 29000 12242 29052 12248
rect 28908 11892 28960 11898
rect 28908 11834 28960 11840
rect 29092 11756 29144 11762
rect 29092 11698 29144 11704
rect 29104 11558 29132 11698
rect 29092 11552 29144 11558
rect 29092 11494 29144 11500
rect 29000 11008 29052 11014
rect 29000 10950 29052 10956
rect 29012 10742 29040 10950
rect 29000 10736 29052 10742
rect 29000 10678 29052 10684
rect 29104 9926 29132 11494
rect 29196 11286 29224 13874
rect 29656 13734 29684 14214
rect 29748 13870 29776 14486
rect 29736 13864 29788 13870
rect 29736 13806 29788 13812
rect 29644 13728 29696 13734
rect 29644 13670 29696 13676
rect 29644 13252 29696 13258
rect 29644 13194 29696 13200
rect 29552 13184 29604 13190
rect 29552 13126 29604 13132
rect 29564 12850 29592 13126
rect 29656 12986 29684 13194
rect 29644 12980 29696 12986
rect 29644 12922 29696 12928
rect 29552 12844 29604 12850
rect 29552 12786 29604 12792
rect 29552 11892 29604 11898
rect 29552 11834 29604 11840
rect 29368 11756 29420 11762
rect 29368 11698 29420 11704
rect 29184 11280 29236 11286
rect 29184 11222 29236 11228
rect 29380 11082 29408 11698
rect 29276 11076 29328 11082
rect 29276 11018 29328 11024
rect 29368 11076 29420 11082
rect 29368 11018 29420 11024
rect 29184 10736 29236 10742
rect 29184 10678 29236 10684
rect 29196 10062 29224 10678
rect 29184 10056 29236 10062
rect 29184 9998 29236 10004
rect 29092 9920 29144 9926
rect 29092 9862 29144 9868
rect 29196 9738 29224 9998
rect 29104 9710 29224 9738
rect 29104 9654 29132 9710
rect 29092 9648 29144 9654
rect 29092 9590 29144 9596
rect 28632 9444 28684 9450
rect 28632 9386 28684 9392
rect 29000 9376 29052 9382
rect 29000 9318 29052 9324
rect 29012 8974 29040 9318
rect 28540 8968 28592 8974
rect 28540 8910 28592 8916
rect 29000 8968 29052 8974
rect 29000 8910 29052 8916
rect 29104 8294 29132 9590
rect 29288 9586 29316 11018
rect 29276 9580 29328 9586
rect 29196 9540 29276 9568
rect 29092 8288 29144 8294
rect 29092 8230 29144 8236
rect 29000 7744 29052 7750
rect 29000 7686 29052 7692
rect 29012 6730 29040 7686
rect 29000 6724 29052 6730
rect 29000 6666 29052 6672
rect 29196 6322 29224 9540
rect 29276 9522 29328 9528
rect 29276 9104 29328 9110
rect 29276 9046 29328 9052
rect 29288 8090 29316 9046
rect 29276 8084 29328 8090
rect 29276 8026 29328 8032
rect 29288 7546 29316 8026
rect 29276 7540 29328 7546
rect 29276 7482 29328 7488
rect 29564 7154 29592 11834
rect 29656 11762 29684 12922
rect 29644 11756 29696 11762
rect 29644 11698 29696 11704
rect 29736 11756 29788 11762
rect 29736 11698 29788 11704
rect 29656 11150 29684 11698
rect 29748 11558 29776 11698
rect 29736 11552 29788 11558
rect 29736 11494 29788 11500
rect 29748 11150 29776 11494
rect 29644 11144 29696 11150
rect 29644 11086 29696 11092
rect 29736 11144 29788 11150
rect 29736 11086 29788 11092
rect 29644 11008 29696 11014
rect 29644 10950 29696 10956
rect 29656 10742 29684 10950
rect 29644 10736 29696 10742
rect 29644 10678 29696 10684
rect 29656 9518 29684 10678
rect 29748 10674 29776 11086
rect 29840 10810 29868 15438
rect 29932 15094 29960 16050
rect 30024 15502 30052 17070
rect 30392 16182 30420 19722
rect 30484 19446 30512 20046
rect 30564 19994 30616 20000
rect 30564 19712 30616 19718
rect 30564 19654 30616 19660
rect 30472 19440 30524 19446
rect 30472 19382 30524 19388
rect 30472 18760 30524 18766
rect 30472 18702 30524 18708
rect 30484 18222 30512 18702
rect 30472 18216 30524 18222
rect 30472 18158 30524 18164
rect 30484 17134 30512 18158
rect 30576 17882 30604 19654
rect 30668 18766 30696 22374
rect 30944 22030 30972 23666
rect 30932 22024 30984 22030
rect 30932 21966 30984 21972
rect 30748 21956 30800 21962
rect 30748 21898 30800 21904
rect 30760 21146 30788 21898
rect 30840 21548 30892 21554
rect 30840 21490 30892 21496
rect 30748 21140 30800 21146
rect 30748 21082 30800 21088
rect 30852 20398 30880 21490
rect 30932 21344 30984 21350
rect 30932 21286 30984 21292
rect 30944 20942 30972 21286
rect 30932 20936 30984 20942
rect 30932 20878 30984 20884
rect 30840 20392 30892 20398
rect 30840 20334 30892 20340
rect 30748 20256 30800 20262
rect 30748 20198 30800 20204
rect 30840 20256 30892 20262
rect 30840 20198 30892 20204
rect 30760 19854 30788 20198
rect 30748 19848 30800 19854
rect 30748 19790 30800 19796
rect 30656 18760 30708 18766
rect 30656 18702 30708 18708
rect 30748 18692 30800 18698
rect 30748 18634 30800 18640
rect 30760 18272 30788 18634
rect 30852 18630 30880 20198
rect 31036 19496 31064 26862
rect 31116 25696 31168 25702
rect 31116 25638 31168 25644
rect 31128 24818 31156 25638
rect 31220 25498 31248 28154
rect 31300 28076 31352 28082
rect 31300 28018 31352 28024
rect 31312 27674 31340 28018
rect 31300 27668 31352 27674
rect 31300 27610 31352 27616
rect 31208 25492 31260 25498
rect 31208 25434 31260 25440
rect 31116 24812 31168 24818
rect 31116 24754 31168 24760
rect 31128 23662 31156 24754
rect 31220 24206 31248 25434
rect 31208 24200 31260 24206
rect 31208 24142 31260 24148
rect 31116 23656 31168 23662
rect 31116 23598 31168 23604
rect 31128 21690 31156 23598
rect 31300 22976 31352 22982
rect 31300 22918 31352 22924
rect 31116 21684 31168 21690
rect 31116 21626 31168 21632
rect 31312 21010 31340 22918
rect 31300 21004 31352 21010
rect 31300 20946 31352 20952
rect 31208 20868 31260 20874
rect 31208 20810 31260 20816
rect 31116 20596 31168 20602
rect 31116 20538 31168 20544
rect 31128 19718 31156 20538
rect 31220 20262 31248 20810
rect 31208 20256 31260 20262
rect 31208 20198 31260 20204
rect 31220 19786 31248 20198
rect 31208 19780 31260 19786
rect 31208 19722 31260 19728
rect 31116 19712 31168 19718
rect 31116 19654 31168 19660
rect 30944 19468 31064 19496
rect 30840 18624 30892 18630
rect 30840 18566 30892 18572
rect 30840 18284 30892 18290
rect 30760 18244 30840 18272
rect 30840 18226 30892 18232
rect 30748 18080 30800 18086
rect 30748 18022 30800 18028
rect 30564 17876 30616 17882
rect 30616 17836 30696 17864
rect 30564 17818 30616 17824
rect 30564 17604 30616 17610
rect 30564 17546 30616 17552
rect 30472 17128 30524 17134
rect 30472 17070 30524 17076
rect 30380 16176 30432 16182
rect 30380 16118 30432 16124
rect 30392 15638 30420 16118
rect 30576 15706 30604 17546
rect 30668 17202 30696 17836
rect 30656 17196 30708 17202
rect 30656 17138 30708 17144
rect 30656 16108 30708 16114
rect 30656 16050 30708 16056
rect 30564 15700 30616 15706
rect 30564 15642 30616 15648
rect 30380 15632 30432 15638
rect 30380 15574 30432 15580
rect 30012 15496 30064 15502
rect 30012 15438 30064 15444
rect 30196 15496 30248 15502
rect 30196 15438 30248 15444
rect 30208 15162 30236 15438
rect 30196 15156 30248 15162
rect 30196 15098 30248 15104
rect 29920 15088 29972 15094
rect 29920 15030 29972 15036
rect 29920 14340 29972 14346
rect 29920 14282 29972 14288
rect 29932 13530 29960 14282
rect 29920 13524 29972 13530
rect 29920 13466 29972 13472
rect 29932 12782 29960 13466
rect 30208 13326 30236 15098
rect 30392 14890 30420 15574
rect 30668 15162 30696 16050
rect 30656 15156 30708 15162
rect 30656 15098 30708 15104
rect 30760 15026 30788 18022
rect 30852 17270 30880 18226
rect 30840 17264 30892 17270
rect 30840 17206 30892 17212
rect 30840 16992 30892 16998
rect 30840 16934 30892 16940
rect 30852 15502 30880 16934
rect 30840 15496 30892 15502
rect 30840 15438 30892 15444
rect 30748 15020 30800 15026
rect 30748 14962 30800 14968
rect 30380 14884 30432 14890
rect 30380 14826 30432 14832
rect 30944 14074 30972 19468
rect 31024 19372 31076 19378
rect 31024 19314 31076 19320
rect 31036 18154 31064 19314
rect 31128 18766 31156 19654
rect 31300 19236 31352 19242
rect 31300 19178 31352 19184
rect 31116 18760 31168 18766
rect 31116 18702 31168 18708
rect 31024 18148 31076 18154
rect 31024 18090 31076 18096
rect 31024 17196 31076 17202
rect 31024 17138 31076 17144
rect 31036 15026 31064 17138
rect 31128 15502 31156 18702
rect 31312 18290 31340 19178
rect 31300 18284 31352 18290
rect 31300 18226 31352 18232
rect 31312 16250 31340 18226
rect 31404 16522 31432 41482
rect 31392 16516 31444 16522
rect 31392 16458 31444 16464
rect 31300 16244 31352 16250
rect 31300 16186 31352 16192
rect 31496 16182 31524 42094
rect 31484 16176 31536 16182
rect 31484 16118 31536 16124
rect 31116 15496 31168 15502
rect 31116 15438 31168 15444
rect 31024 15020 31076 15026
rect 31024 14962 31076 14968
rect 30932 14068 30984 14074
rect 30984 14028 31064 14056
rect 30932 14010 30984 14016
rect 30932 13932 30984 13938
rect 30932 13874 30984 13880
rect 30840 13864 30892 13870
rect 30840 13806 30892 13812
rect 30196 13320 30248 13326
rect 30196 13262 30248 13268
rect 30288 12844 30340 12850
rect 30288 12786 30340 12792
rect 29920 12776 29972 12782
rect 29920 12718 29972 12724
rect 29932 11354 29960 12718
rect 30196 12640 30248 12646
rect 30196 12582 30248 12588
rect 30208 12238 30236 12582
rect 30196 12232 30248 12238
rect 30196 12174 30248 12180
rect 30012 12096 30064 12102
rect 30012 12038 30064 12044
rect 29920 11348 29972 11354
rect 29920 11290 29972 11296
rect 29828 10804 29880 10810
rect 29828 10746 29880 10752
rect 29736 10668 29788 10674
rect 29736 10610 29788 10616
rect 30024 9586 30052 12038
rect 30300 11898 30328 12786
rect 30852 12170 30880 13806
rect 30944 13530 30972 13874
rect 30932 13524 30984 13530
rect 30932 13466 30984 13472
rect 30944 12850 30972 13466
rect 31036 13190 31064 14028
rect 31116 13932 31168 13938
rect 31116 13874 31168 13880
rect 31128 13530 31156 13874
rect 31116 13524 31168 13530
rect 31116 13466 31168 13472
rect 31024 13184 31076 13190
rect 31024 13126 31076 13132
rect 30932 12844 30984 12850
rect 30932 12786 30984 12792
rect 31036 12442 31064 13126
rect 31208 12844 31260 12850
rect 31208 12786 31260 12792
rect 31024 12436 31076 12442
rect 31024 12378 31076 12384
rect 30840 12164 30892 12170
rect 30840 12106 30892 12112
rect 30288 11892 30340 11898
rect 30288 11834 30340 11840
rect 31036 11762 31064 12378
rect 31024 11756 31076 11762
rect 31024 11698 31076 11704
rect 30196 11144 30248 11150
rect 30196 11086 30248 11092
rect 30840 11144 30892 11150
rect 30840 11086 30892 11092
rect 30104 11076 30156 11082
rect 30104 11018 30156 11024
rect 30116 10062 30144 11018
rect 30208 10810 30236 11086
rect 30852 10810 30880 11086
rect 30196 10804 30248 10810
rect 30196 10746 30248 10752
rect 30840 10804 30892 10810
rect 30840 10746 30892 10752
rect 31220 10674 31248 12786
rect 31300 11620 31352 11626
rect 31300 11562 31352 11568
rect 31208 10668 31260 10674
rect 31208 10610 31260 10616
rect 31220 10266 31248 10610
rect 31208 10260 31260 10266
rect 31208 10202 31260 10208
rect 30104 10056 30156 10062
rect 30104 9998 30156 10004
rect 30012 9580 30064 9586
rect 30012 9522 30064 9528
rect 29644 9512 29696 9518
rect 29644 9454 29696 9460
rect 29656 9042 29684 9454
rect 30932 9444 30984 9450
rect 30932 9386 30984 9392
rect 29644 9036 29696 9042
rect 29644 8978 29696 8984
rect 30944 8974 30972 9386
rect 31116 9376 31168 9382
rect 31116 9318 31168 9324
rect 30932 8968 30984 8974
rect 30932 8910 30984 8916
rect 30380 8900 30432 8906
rect 30380 8842 30432 8848
rect 29828 8832 29880 8838
rect 29828 8774 29880 8780
rect 29736 8492 29788 8498
rect 29736 8434 29788 8440
rect 29644 8288 29696 8294
rect 29644 8230 29696 8236
rect 29656 7886 29684 8230
rect 29644 7880 29696 7886
rect 29644 7822 29696 7828
rect 29656 7478 29684 7822
rect 29644 7472 29696 7478
rect 29644 7414 29696 7420
rect 29656 7342 29684 7414
rect 29644 7336 29696 7342
rect 29644 7278 29696 7284
rect 29564 7126 29684 7154
rect 29276 6452 29328 6458
rect 29276 6394 29328 6400
rect 29184 6316 29236 6322
rect 29184 6258 29236 6264
rect 28632 6112 28684 6118
rect 28632 6054 28684 6060
rect 28644 5030 28672 6054
rect 28736 5778 29132 5794
rect 28724 5772 29132 5778
rect 28776 5766 29132 5772
rect 28724 5714 28776 5720
rect 29104 5030 29132 5766
rect 28632 5024 28684 5030
rect 28632 4966 28684 4972
rect 29092 5024 29144 5030
rect 29092 4966 29144 4972
rect 28540 4616 28592 4622
rect 28540 4558 28592 4564
rect 28552 4146 28580 4558
rect 28540 4140 28592 4146
rect 28540 4082 28592 4088
rect 28552 2990 28580 4082
rect 29104 4078 29132 4966
rect 29196 4690 29224 6258
rect 29288 5710 29316 6394
rect 29276 5704 29328 5710
rect 29276 5646 29328 5652
rect 29460 5568 29512 5574
rect 29460 5510 29512 5516
rect 29184 4684 29236 4690
rect 29184 4626 29236 4632
rect 29368 4548 29420 4554
rect 29368 4490 29420 4496
rect 29380 4282 29408 4490
rect 29368 4276 29420 4282
rect 29368 4218 29420 4224
rect 29472 4146 29500 5510
rect 29552 5160 29604 5166
rect 29552 5102 29604 5108
rect 29564 4690 29592 5102
rect 29552 4684 29604 4690
rect 29552 4626 29604 4632
rect 29460 4140 29512 4146
rect 29460 4082 29512 4088
rect 29092 4072 29144 4078
rect 29092 4014 29144 4020
rect 28632 3936 28684 3942
rect 28632 3878 28684 3884
rect 28644 3602 28672 3878
rect 28632 3596 28684 3602
rect 28632 3538 28684 3544
rect 28724 3460 28776 3466
rect 28724 3402 28776 3408
rect 28736 2990 28764 3402
rect 28540 2984 28592 2990
rect 28540 2926 28592 2932
rect 28724 2984 28776 2990
rect 28724 2926 28776 2932
rect 28552 2446 28580 2926
rect 28908 2916 28960 2922
rect 28908 2858 28960 2864
rect 28540 2440 28592 2446
rect 28540 2382 28592 2388
rect 28816 2440 28868 2446
rect 28816 2382 28868 2388
rect 28828 1834 28856 2382
rect 28920 2038 28948 2858
rect 29092 2644 29144 2650
rect 29092 2586 29144 2592
rect 28908 2032 28960 2038
rect 28908 1974 28960 1980
rect 28816 1828 28868 1834
rect 28816 1770 28868 1776
rect 28816 1556 28868 1562
rect 28816 1498 28868 1504
rect 28828 1290 28856 1498
rect 29000 1352 29052 1358
rect 29000 1294 29052 1300
rect 28816 1284 28868 1290
rect 28816 1226 28868 1232
rect 29012 882 29040 1294
rect 29000 876 29052 882
rect 29000 818 29052 824
rect 29104 746 29132 2586
rect 29656 1494 29684 7126
rect 29748 6866 29776 8434
rect 29840 7886 29868 8774
rect 30196 8356 30248 8362
rect 30196 8298 30248 8304
rect 29828 7880 29880 7886
rect 29828 7822 29880 7828
rect 30208 7478 30236 8298
rect 30288 7540 30340 7546
rect 30288 7482 30340 7488
rect 30196 7472 30248 7478
rect 30196 7414 30248 7420
rect 29920 7336 29972 7342
rect 29920 7278 29972 7284
rect 29736 6860 29788 6866
rect 29736 6802 29788 6808
rect 29736 6180 29788 6186
rect 29736 6122 29788 6128
rect 29748 4010 29776 6122
rect 29828 5840 29880 5846
rect 29828 5782 29880 5788
rect 29840 4146 29868 5782
rect 29932 5166 29960 7278
rect 30300 6798 30328 7482
rect 30288 6792 30340 6798
rect 30288 6734 30340 6740
rect 30196 6656 30248 6662
rect 30196 6598 30248 6604
rect 30012 5636 30064 5642
rect 30012 5578 30064 5584
rect 29920 5160 29972 5166
rect 29920 5102 29972 5108
rect 30024 4486 30052 5578
rect 30208 5234 30236 6598
rect 30392 6458 30420 8842
rect 30656 8832 30708 8838
rect 30656 8774 30708 8780
rect 30564 6792 30616 6798
rect 30564 6734 30616 6740
rect 30472 6724 30524 6730
rect 30472 6666 30524 6672
rect 30380 6452 30432 6458
rect 30380 6394 30432 6400
rect 30484 6322 30512 6666
rect 30472 6316 30524 6322
rect 30472 6258 30524 6264
rect 30484 5710 30512 6258
rect 30472 5704 30524 5710
rect 30472 5646 30524 5652
rect 30484 5574 30512 5646
rect 30472 5568 30524 5574
rect 30472 5510 30524 5516
rect 30380 5296 30432 5302
rect 30380 5238 30432 5244
rect 30196 5228 30248 5234
rect 30196 5170 30248 5176
rect 30012 4480 30064 4486
rect 30012 4422 30064 4428
rect 29828 4140 29880 4146
rect 29828 4082 29880 4088
rect 30104 4072 30156 4078
rect 30104 4014 30156 4020
rect 29736 4004 29788 4010
rect 29736 3946 29788 3952
rect 29748 3670 29776 3946
rect 29736 3664 29788 3670
rect 29736 3606 29788 3612
rect 29736 3528 29788 3534
rect 29736 3470 29788 3476
rect 30012 3528 30064 3534
rect 30012 3470 30064 3476
rect 29748 2446 29776 3470
rect 30024 2446 30052 3470
rect 30116 2514 30144 4014
rect 30104 2508 30156 2514
rect 30104 2450 30156 2456
rect 29736 2440 29788 2446
rect 29736 2382 29788 2388
rect 30012 2440 30064 2446
rect 30012 2382 30064 2388
rect 30288 2440 30340 2446
rect 30288 2382 30340 2388
rect 30300 1834 30328 2382
rect 30288 1828 30340 1834
rect 30288 1770 30340 1776
rect 29644 1488 29696 1494
rect 29644 1430 29696 1436
rect 29736 1352 29788 1358
rect 29736 1294 29788 1300
rect 29748 1018 29776 1294
rect 29736 1012 29788 1018
rect 29736 954 29788 960
rect 30392 800 30420 5238
rect 30484 4146 30512 5510
rect 30472 4140 30524 4146
rect 30472 4082 30524 4088
rect 30576 4078 30604 6734
rect 30668 6118 30696 8774
rect 30748 6860 30800 6866
rect 30748 6802 30800 6808
rect 30760 6322 30788 6802
rect 30748 6316 30800 6322
rect 30748 6258 30800 6264
rect 30656 6112 30708 6118
rect 30656 6054 30708 6060
rect 30760 5710 30788 6258
rect 30748 5704 30800 5710
rect 30748 5646 30800 5652
rect 30656 5024 30708 5030
rect 30656 4966 30708 4972
rect 30564 4072 30616 4078
rect 30564 4014 30616 4020
rect 30668 3738 30696 4966
rect 30760 4146 30788 5646
rect 30944 5522 30972 8910
rect 31128 8634 31156 9318
rect 31312 8974 31340 11562
rect 31300 8968 31352 8974
rect 31300 8910 31352 8916
rect 31392 8900 31444 8906
rect 31392 8842 31444 8848
rect 31116 8628 31168 8634
rect 31116 8570 31168 8576
rect 31024 8492 31076 8498
rect 31024 8434 31076 8440
rect 31036 5914 31064 8434
rect 31300 8424 31352 8430
rect 31300 8366 31352 8372
rect 31312 8090 31340 8366
rect 31404 8362 31432 8842
rect 31392 8356 31444 8362
rect 31392 8298 31444 8304
rect 31300 8084 31352 8090
rect 31300 8026 31352 8032
rect 31208 7744 31260 7750
rect 31208 7686 31260 7692
rect 31220 7546 31248 7686
rect 31208 7540 31260 7546
rect 31128 7500 31208 7528
rect 31128 6866 31156 7500
rect 31208 7482 31260 7488
rect 31116 6860 31168 6866
rect 31116 6802 31168 6808
rect 31024 5908 31076 5914
rect 31024 5850 31076 5856
rect 31128 5710 31156 6802
rect 31312 6322 31340 8026
rect 31404 6798 31432 8298
rect 31392 6792 31444 6798
rect 31392 6734 31444 6740
rect 31300 6316 31352 6322
rect 31300 6258 31352 6264
rect 31116 5704 31168 5710
rect 31116 5646 31168 5652
rect 30944 5494 31248 5522
rect 31116 4480 31168 4486
rect 31116 4422 31168 4428
rect 30748 4140 30800 4146
rect 30748 4082 30800 4088
rect 30656 3732 30708 3738
rect 30656 3674 30708 3680
rect 31024 3664 31076 3670
rect 31024 3606 31076 3612
rect 30748 3460 30800 3466
rect 30748 3402 30800 3408
rect 30564 3392 30616 3398
rect 30564 3334 30616 3340
rect 30576 2446 30604 3334
rect 30760 3194 30788 3402
rect 30748 3188 30800 3194
rect 30748 3130 30800 3136
rect 30656 3052 30708 3058
rect 30656 2994 30708 3000
rect 30668 2650 30696 2994
rect 30656 2644 30708 2650
rect 30656 2586 30708 2592
rect 31036 2446 31064 3606
rect 31128 3602 31156 4422
rect 31116 3596 31168 3602
rect 31116 3538 31168 3544
rect 31116 3188 31168 3194
rect 31116 3130 31168 3136
rect 30564 2440 30616 2446
rect 30564 2382 30616 2388
rect 31024 2440 31076 2446
rect 31024 2382 31076 2388
rect 30840 2304 30892 2310
rect 30840 2246 30892 2252
rect 30656 1964 30708 1970
rect 30656 1906 30708 1912
rect 30668 1562 30696 1906
rect 30656 1556 30708 1562
rect 30656 1498 30708 1504
rect 30852 1358 30880 2246
rect 31036 1426 31064 2382
rect 31024 1420 31076 1426
rect 31024 1362 31076 1368
rect 31128 1358 31156 3130
rect 31220 3126 31248 5494
rect 31300 5024 31352 5030
rect 31300 4966 31352 4972
rect 31312 4214 31340 4966
rect 31300 4208 31352 4214
rect 31300 4150 31352 4156
rect 31208 3120 31260 3126
rect 31208 3062 31260 3068
rect 31300 1964 31352 1970
rect 31300 1906 31352 1912
rect 30840 1352 30892 1358
rect 30840 1294 30892 1300
rect 31116 1352 31168 1358
rect 31116 1294 31168 1300
rect 31312 814 31340 1906
rect 31300 808 31352 814
rect 29092 740 29144 746
rect 29092 682 29144 688
rect 28448 672 28500 678
rect 28448 614 28500 620
rect 30378 0 30434 800
rect 31300 750 31352 756
use sky130_fd_sc_hd__diode_2  ANTENNA_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21988 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform -1 0 2024 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_0_3 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1380 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_11
timestamp 1644511149
transform 1 0 2116 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_0_19 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2852 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_0_33
timestamp 1644511149
transform 1 0 4140 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_0_41
timestamp 1644511149
transform 1 0 4876 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_0_52
timestamp 1644511149
transform 1 0 5888 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_63
timestamp 1644511149
transform 1 0 6900 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_73
timestamp 1644511149
transform 1 0 7820 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_80
timestamp 1644511149
transform 1 0 8464 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_95
timestamp 1644511149
transform 1 0 9844 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_105
timestamp 1644511149
transform 1 0 10764 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_109 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11132 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1644511149
transform 1 0 11316 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_0_118
timestamp 1644511149
transform 1 0 11960 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_129
timestamp 1644511149
transform 1 0 12972 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_0_136
timestamp 1644511149
transform 1 0 13616 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_144
timestamp 1644511149
transform 1 0 14352 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_154
timestamp 1644511149
transform 1 0 15272 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_164
timestamp 1644511149
transform 1 0 16192 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_175
timestamp 1644511149
transform 1 0 17204 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_182
timestamp 1644511149
transform 1 0 17848 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_192
timestamp 1644511149
transform 1 0 18768 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_0_202
timestamp 1644511149
transform 1 0 19688 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_209
timestamp 1644511149
transform 1 0 20332 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_213
timestamp 1644511149
transform 1 0 20700 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_0_220
timestamp 1644511149
transform 1 0 21344 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_228
timestamp 1644511149
transform 1 0 22080 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_238
timestamp 1644511149
transform 1 0 23000 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_248
timestamp 1644511149
transform 1 0 23920 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_255
timestamp 1644511149
transform 1 0 24564 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_0_262
timestamp 1644511149
transform 1 0 25208 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_266
timestamp 1644511149
transform 1 0 25576 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_0_274
timestamp 1644511149
transform 1 0 26312 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1644511149
transform 1 0 26680 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_283
timestamp 1644511149
transform 1 0 27140 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_0_287
timestamp 1644511149
transform 1 0 27508 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_297
timestamp 1644511149
transform 1 0 28428 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_0_304
timestamp 1644511149
transform 1 0 29072 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_0_312
timestamp 1644511149
transform 1 0 29808 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_320
timestamp 1644511149
transform 1 0 30544 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_0_327
timestamp 1644511149
transform 1 0 31188 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_331
timestamp 1644511149
transform 1 0 31556 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_1_7
timestamp 1644511149
transform 1 0 1748 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_17
timestamp 1644511149
transform 1 0 2668 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_21
timestamp 1644511149
transform 1 0 3036 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_1_28
timestamp 1644511149
transform 1 0 3680 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_1_52
timestamp 1644511149
transform 1 0 5888 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_1_62
timestamp 1644511149
transform 1 0 6808 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_1_82
timestamp 1644511149
transform 1 0 8648 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_90
timestamp 1644511149
transform 1 0 9384 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_1_108
timestamp 1644511149
transform 1 0 11040 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_129
timestamp 1644511149
transform 1 0 12972 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_139
timestamp 1644511149
transform 1 0 13892 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_143
timestamp 1644511149
transform 1 0 14260 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_145
timestamp 1644511149
transform 1 0 14444 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_1_162
timestamp 1644511149
transform 1 0 16008 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1644511149
transform 1 0 16376 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_1_179
timestamp 1644511149
transform 1 0 17572 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_183
timestamp 1644511149
transform 1 0 17940 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_1_200
timestamp 1644511149
transform 1 0 19504 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_220
timestamp 1644511149
transform 1 0 21344 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_1_242
timestamp 1644511149
transform 1 0 23368 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_246
timestamp 1644511149
transform 1 0 23736 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_248
timestamp 1644511149
transform 1 0 23920 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_1_265
timestamp 1644511149
transform 1 0 25484 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_269
timestamp 1644511149
transform 1 0 25852 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_1_276
timestamp 1644511149
transform 1 0 26496 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_285
timestamp 1644511149
transform 1 0 27324 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_1_302
timestamp 1644511149
transform 1 0 28888 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_322
timestamp 1644511149
transform 1 0 30728 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_1_329
timestamp 1644511149
transform 1 0 31372 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_2_21
timestamp 1644511149
transform 1 0 3036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_25
timestamp 1644511149
transform 1 0 3404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_2_45
timestamp 1644511149
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_53
timestamp 1644511149
transform 1 0 5980 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_2_66
timestamp 1644511149
transform 1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_80
timestamp 1644511149
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_101
timestamp 1644511149
transform 1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_109
timestamp 1644511149
transform 1 0 11132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_129
timestamp 1644511149
transform 1 0 12972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_136
timestamp 1644511149
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_145
timestamp 1644511149
transform 1 0 14444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_2_162
timestamp 1644511149
transform 1 0 16008 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_182
timestamp 1644511149
transform 1 0 17848 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_192
timestamp 1644511149
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_213
timestamp 1644511149
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_217
timestamp 1644511149
transform 1 0 21068 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1644511149
transform 1 0 21252 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_2_236
timestamp 1644511149
transform 1 0 22816 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_248
timestamp 1644511149
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_2_270
timestamp 1644511149
transform 1 0 25944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_290
timestamp 1644511149
transform 1 0 27784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_302
timestamp 1644511149
transform 1 0 28888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_306
timestamp 1644511149
transform 1 0 29256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_2_317
timestamp 1644511149
transform 1 0 30268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_2_327
timestamp 1644511149
transform 1 0 31188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_331
timestamp 1644511149
transform 1 0 31556 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_7
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_3_17
timestamp 1644511149
transform 1 0 2668 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_3_29
timestamp 1644511149
transform 1 0 3772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_33
timestamp 1644511149
transform 1 0 4140 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_35
timestamp 1644511149
transform 1 0 4324 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_3_52
timestamp 1644511149
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_3_65
timestamp 1644511149
transform 1 0 7084 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_3_79
timestamp 1644511149
transform 1 0 8372 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_3_88
timestamp 1644511149
transform 1 0 9200 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_3_108
timestamp 1644511149
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_3_119
timestamp 1644511149
transform 1 0 12052 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_3_143
timestamp 1644511149
transform 1 0 14260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_3_155
timestamp 1644511149
transform 1 0 15364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_3_162
timestamp 1644511149
transform 1 0 16008 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1644511149
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_3_177
timestamp 1644511149
transform 1 0 17388 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_3_193
timestamp 1644511149
transform 1 0 18860 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_197
timestamp 1644511149
transform 1 0 19228 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_199
timestamp 1644511149
transform 1 0 19412 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_3_206
timestamp 1644511149
transform 1 0 20056 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_3_218
timestamp 1644511149
transform 1 0 21160 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1644511149
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_227
timestamp 1644511149
transform 1 0 21988 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_3_236
timestamp 1644511149
transform 1 0 22816 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_3_256
timestamp 1644511149
transform 1 0 24656 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_260
timestamp 1644511149
transform 1 0 25024 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_262
timestamp 1644511149
transform 1 0 25208 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_3_271
timestamp 1644511149
transform 1 0 26036 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_285
timestamp 1644511149
transform 1 0 27324 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_3_294
timestamp 1644511149
transform 1 0 28152 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_298
timestamp 1644511149
transform 1 0 28520 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_3_303
timestamp 1644511149
transform 1 0 28980 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_3_323
timestamp 1644511149
transform 1 0 30820 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_331
timestamp 1644511149
transform 1 0 31556 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_7
timestamp 1644511149
transform 1 0 1748 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_4_14
timestamp 1644511149
transform 1 0 2392 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_4_24
timestamp 1644511149
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_4_43
timestamp 1644511149
transform 1 0 5060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_57
timestamp 1644511149
transform 1 0 6348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_4_76
timestamp 1644511149
transform 1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_4_94
timestamp 1644511149
transform 1 0 9752 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_4_106
timestamp 1644511149
transform 1 0 10856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_110
timestamp 1644511149
transform 1 0 11224 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_112
timestamp 1644511149
transform 1 0 11408 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_4_129
timestamp 1644511149
transform 1 0 12972 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_4_136
timestamp 1644511149
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_4_149
timestamp 1644511149
transform 1 0 14812 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_181
timestamp 1644511149
transform 1 0 17756 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_183
timestamp 1644511149
transform 1 0 17940 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_4_192
timestamp 1644511149
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_4_200
timestamp 1644511149
transform 1 0 19504 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_4_212
timestamp 1644511149
transform 1 0 20608 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_4_224
timestamp 1644511149
transform 1 0 21712 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_4_236
timestamp 1644511149
transform 1 0 22816 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_240
timestamp 1644511149
transform 1 0 23184 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_4_248
timestamp 1644511149
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_269
timestamp 1644511149
transform 1 0 25852 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_305
timestamp 1644511149
transform 1 0 29164 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_4_317
timestamp 1644511149
transform 1 0 30268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_4_327
timestamp 1644511149
transform 1 0 31188 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_331
timestamp 1644511149
transform 1 0 31556 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_7
timestamp 1644511149
transform 1 0 1748 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_5_17
timestamp 1644511149
transform 1 0 2668 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_5_30
timestamp 1644511149
transform 1 0 3864 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_5_50
timestamp 1644511149
transform 1 0 5704 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1644511149
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_5_66
timestamp 1644511149
transform 1 0 7176 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_5_76
timestamp 1644511149
transform 1 0 8096 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_5_84
timestamp 1644511149
transform 1 0 8832 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_5_96
timestamp 1644511149
transform 1 0 9936 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_5_106
timestamp 1644511149
transform 1 0 10856 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1644511149
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_165
timestamp 1644511149
transform 1 0 16284 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_171
timestamp 1644511149
transform 1 0 16836 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_5_180
timestamp 1644511149
transform 1 0 17664 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_184
timestamp 1644511149
transform 1 0 18032 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_5_200
timestamp 1644511149
transform 1 0 19504 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_5_220
timestamp 1644511149
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_5_228
timestamp 1644511149
transform 1 0 22080 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_232
timestamp 1644511149
transform 1 0 22448 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_5_243
timestamp 1644511149
transform 1 0 23460 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_5_257
timestamp 1644511149
transform 1 0 24748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_5_269
timestamp 1644511149
transform 1 0 25852 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_5_276
timestamp 1644511149
transform 1 0 26496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_5_289
timestamp 1644511149
transform 1 0 27692 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_5_301
timestamp 1644511149
transform 1 0 28796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_5_313
timestamp 1644511149
transform 1 0 29900 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_5_325
timestamp 1644511149
transform 1 0 31004 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_19
timestamp 1644511149
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_6_47
timestamp 1644511149
transform 1 0 5428 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_51
timestamp 1644511149
transform 1 0 5796 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_6_61
timestamp 1644511149
transform 1 0 6716 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_6_75
timestamp 1644511149
transform 1 0 8004 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_89
timestamp 1644511149
transform 1 0 9292 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_6_107
timestamp 1644511149
transform 1 0 10948 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_111
timestamp 1644511149
transform 1 0 11316 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_6_129
timestamp 1644511149
transform 1 0 12972 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_6_136
timestamp 1644511149
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_6_151
timestamp 1644511149
transform 1 0 14996 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_6_162
timestamp 1644511149
transform 1 0 16008 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_170
timestamp 1644511149
transform 1 0 16744 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_6_182
timestamp 1644511149
transform 1 0 17848 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_6_192
timestamp 1644511149
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_6_200
timestamp 1644511149
transform 1 0 19504 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_6_210
timestamp 1644511149
transform 1 0 20424 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_6_220
timestamp 1644511149
transform 1 0 21344 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_6_244
timestamp 1644511149
transform 1 0 23552 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_6_283
timestamp 1644511149
transform 1 0 27140 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_6_290
timestamp 1644511149
transform 1 0 27784 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_6_304
timestamp 1644511149
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_6_325
timestamp 1644511149
transform 1 0 31004 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7
timestamp 1644511149
transform 1 0 1748 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_7_14
timestamp 1644511149
transform 1 0 2392 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_7_34
timestamp 1644511149
transform 1 0 4232 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_7_42
timestamp 1644511149
transform 1 0 4968 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_7_52
timestamp 1644511149
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_7_65
timestamp 1644511149
transform 1 0 7084 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_7_88
timestamp 1644511149
transform 1 0 9200 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_7_102
timestamp 1644511149
transform 1 0 10488 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1644511149
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_115
timestamp 1644511149
transform 1 0 11684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_7_122
timestamp 1644511149
transform 1 0 12328 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_7_136
timestamp 1644511149
transform 1 0 13616 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_7_148
timestamp 1644511149
transform 1 0 14720 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_7_159
timestamp 1644511149
transform 1 0 15732 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_7_177
timestamp 1644511149
transform 1 0 17388 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_7_201
timestamp 1644511149
transform 1 0 19596 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_7_211
timestamp 1644511149
transform 1 0 20516 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_7_220
timestamp 1644511149
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_7_244
timestamp 1644511149
transform 1 0 23552 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_7_264
timestamp 1644511149
transform 1 0 25392 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_7_276
timestamp 1644511149
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_7_285
timestamp 1644511149
transform 1 0 27324 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_6
timestamp 1644511149
transform 1 0 1656 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_8_14
timestamp 1644511149
transform 1 0 2392 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_8_24
timestamp 1644511149
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_8_38
timestamp 1644511149
transform 1 0 4600 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_42
timestamp 1644511149
transform 1 0 4968 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_8_59
timestamp 1644511149
transform 1 0 6532 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_8_72
timestamp 1644511149
transform 1 0 7728 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_8_80
timestamp 1644511149
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_8_94
timestamp 1644511149
transform 1 0 9752 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_8_114
timestamp 1644511149
transform 1 0 11592 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_8_131
timestamp 1644511149
transform 1 0 13156 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_145
timestamp 1644511149
transform 1 0 14444 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_8_154
timestamp 1644511149
transform 1 0 15272 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_8_163
timestamp 1644511149
transform 1 0 16100 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_167
timestamp 1644511149
transform 1 0 16468 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_8_176
timestamp 1644511149
transform 1 0 17296 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_180
timestamp 1644511149
transform 1 0 17664 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_8_188
timestamp 1644511149
transform 1 0 18400 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_8_213
timestamp 1644511149
transform 1 0 20700 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_8_242
timestamp 1644511149
transform 1 0 23368 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1644511149
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_8_271
timestamp 1644511149
transform 1 0 26036 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_8_278
timestamp 1644511149
transform 1 0 26680 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_8_290
timestamp 1644511149
transform 1 0 27784 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_294
timestamp 1644511149
transform 1 0 28152 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_8_304
timestamp 1644511149
transform 1 0 29072 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_8_312
timestamp 1644511149
transform 1 0 29808 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_316
timestamp 1644511149
transform 1 0 30176 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_318
timestamp 1644511149
transform 1 0 30360 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_8_327
timestamp 1644511149
transform 1 0 31188 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_331
timestamp 1644511149
transform 1 0 31556 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_9_13
timestamp 1644511149
transform 1 0 2300 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_21
timestamp 1644511149
transform 1 0 3036 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_9_43
timestamp 1644511149
transform 1 0 5060 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_59
timestamp 1644511149
transform 1 0 6532 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_9_70
timestamp 1644511149
transform 1 0 7544 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_9_84
timestamp 1644511149
transform 1 0 8832 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_9_96
timestamp 1644511149
transform 1 0 9936 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_9_106
timestamp 1644511149
transform 1 0 10856 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1644511149
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_9_117
timestamp 1644511149
transform 1 0 11868 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_9_127
timestamp 1644511149
transform 1 0 12788 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_135
timestamp 1644511149
transform 1 0 13524 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_9_144
timestamp 1644511149
transform 1 0 14352 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_9_152
timestamp 1644511149
transform 1 0 15088 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_156
timestamp 1644511149
transform 1 0 15456 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_9_164
timestamp 1644511149
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_9_177
timestamp 1644511149
transform 1 0 17388 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_9_184
timestamp 1644511149
transform 1 0 18032 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_9_208
timestamp 1644511149
transform 1 0 20240 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_9_218
timestamp 1644511149
transform 1 0 21160 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1644511149
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_229
timestamp 1644511149
transform 1 0 22172 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_9_236
timestamp 1644511149
transform 1 0 22816 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_240
timestamp 1644511149
transform 1 0 23184 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_242
timestamp 1644511149
transform 1 0 23368 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_265
timestamp 1644511149
transform 1 0 25484 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_277
timestamp 1644511149
transform 1 0 26588 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_9_288
timestamp 1644511149
transform 1 0 27600 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_292
timestamp 1644511149
transform 1 0 27968 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_9_297
timestamp 1644511149
transform 1 0 28428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_9_315
timestamp 1644511149
transform 1 0 30084 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_9_327
timestamp 1644511149
transform 1 0 31188 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_331
timestamp 1644511149
transform 1 0 31556 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_10_19
timestamp 1644511149
transform 1 0 2852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_10_35
timestamp 1644511149
transform 1 0 4324 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_57
timestamp 1644511149
transform 1 0 6348 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_59
timestamp 1644511149
transform 1 0 6532 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_10_80
timestamp 1644511149
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_10_95
timestamp 1644511149
transform 1 0 9844 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_10_105
timestamp 1644511149
transform 1 0 10764 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_10_127
timestamp 1644511149
transform 1 0 12788 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_10_135
timestamp 1644511149
transform 1 0 13524 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_143
timestamp 1644511149
transform 1 0 14260 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_169
timestamp 1644511149
transform 1 0 16652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_10_176
timestamp 1644511149
transform 1 0 17296 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_10_186
timestamp 1644511149
transform 1 0 18216 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1644511149
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_10_204
timestamp 1644511149
transform 1 0 19872 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_10_224
timestamp 1644511149
transform 1 0 21712 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_228
timestamp 1644511149
transform 1 0 22080 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_230
timestamp 1644511149
transform 1 0 22264 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_10_236
timestamp 1644511149
transform 1 0 22816 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_10_248
timestamp 1644511149
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_10_256
timestamp 1644511149
transform 1 0 24656 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_10_269
timestamp 1644511149
transform 1 0 25852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_10_286
timestamp 1644511149
transform 1 0 27416 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_290
timestamp 1644511149
transform 1 0 27784 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_292
timestamp 1644511149
transform 1 0 27968 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_10_303
timestamp 1644511149
transform 1 0 28980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_10_319
timestamp 1644511149
transform 1 0 30452 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_10_329
timestamp 1644511149
transform 1 0 31372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_11_6
timestamp 1644511149
transform 1 0 1656 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_11_18
timestamp 1644511149
transform 1 0 2760 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_11_34
timestamp 1644511149
transform 1 0 4232 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_42
timestamp 1644511149
transform 1 0 4968 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_11_52
timestamp 1644511149
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_11_63
timestamp 1644511149
transform 1 0 6900 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_67
timestamp 1644511149
transform 1 0 7268 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_11_84
timestamp 1644511149
transform 1 0 8832 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_11_108
timestamp 1644511149
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_11_130
timestamp 1644511149
transform 1 0 13064 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_11_142
timestamp 1644511149
transform 1 0 14168 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_11_154
timestamp 1644511149
transform 1 0 15272 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_11_164
timestamp 1644511149
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_11_177
timestamp 1644511149
transform 1 0 17388 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_183
timestamp 1644511149
transform 1 0 17940 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_11_200
timestamp 1644511149
transform 1 0 19504 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_11_213
timestamp 1644511149
transform 1 0 20700 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_11_220
timestamp 1644511149
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_11_232
timestamp 1644511149
transform 1 0 22448 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_240
timestamp 1644511149
transform 1 0 23184 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_11_259
timestamp 1644511149
transform 1 0 24932 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_11_276
timestamp 1644511149
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_11_287
timestamp 1644511149
transform 1 0 27508 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_11_307
timestamp 1644511149
transform 1 0 29348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_311
timestamp 1644511149
transform 1 0 29716 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_12_6
timestamp 1644511149
transform 1 0 1656 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_12_18
timestamp 1644511149
transform 1 0 2760 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1644511149
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_12_35
timestamp 1644511149
transform 1 0 4324 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_12_47
timestamp 1644511149
transform 1 0 5428 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_51
timestamp 1644511149
transform 1 0 5796 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_12_61
timestamp 1644511149
transform 1 0 6716 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_12_68
timestamp 1644511149
transform 1 0 7360 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_12_78
timestamp 1644511149
transform 1 0 8280 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1644511149
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_12_91
timestamp 1644511149
transform 1 0 9476 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_95
timestamp 1644511149
transform 1 0 9844 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_12_105
timestamp 1644511149
transform 1 0 10764 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_12_117
timestamp 1644511149
transform 1 0 11868 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_12_128
timestamp 1644511149
transform 1 0 12880 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_12_136
timestamp 1644511149
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_12_151
timestamp 1644511149
transform 1 0 14996 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_12_163
timestamp 1644511149
transform 1 0 16100 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_171
timestamp 1644511149
transform 1 0 16836 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_193
timestamp 1644511149
transform 1 0 18860 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_12_215
timestamp 1644511149
transform 1 0 20884 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_12_227
timestamp 1644511149
transform 1 0 21988 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_12_247
timestamp 1644511149
transform 1 0 23828 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_12_262
timestamp 1644511149
transform 1 0 25208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_12_269
timestamp 1644511149
transform 1 0 25852 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_12_279
timestamp 1644511149
transform 1 0 26772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_12_304
timestamp 1644511149
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_12_325
timestamp 1644511149
transform 1 0 31004 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1644511149
transform 1 0 1748 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_13_12
timestamp 1644511149
transform 1 0 2208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_13_25
timestamp 1644511149
transform 1 0 3404 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_13_49
timestamp 1644511149
transform 1 0 5612 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_53
timestamp 1644511149
transform 1 0 5980 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_13_73
timestamp 1644511149
transform 1 0 7820 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_13_86
timestamp 1644511149
transform 1 0 9016 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_13_97
timestamp 1644511149
transform 1 0 10028 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_13_107
timestamp 1644511149
transform 1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_13_117
timestamp 1644511149
transform 1 0 11868 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_13_145
timestamp 1644511149
transform 1 0 14444 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_153
timestamp 1644511149
transform 1 0 15180 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_13_164
timestamp 1644511149
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_13_185
timestamp 1644511149
transform 1 0 18124 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_13_202
timestamp 1644511149
transform 1 0 19688 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_13_214
timestamp 1644511149
transform 1 0 20792 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1644511149
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_13_244
timestamp 1644511149
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_13_253
timestamp 1644511149
transform 1 0 24380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_13_267
timestamp 1644511149
transform 1 0 25668 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_13_275
timestamp 1644511149
transform 1 0 26404 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_13_285
timestamp 1644511149
transform 1 0 27324 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_13_295
timestamp 1644511149
transform 1 0 28244 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_13_319
timestamp 1644511149
transform 1 0 30452 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_7
timestamp 1644511149
transform 1 0 1748 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_14_18
timestamp 1644511149
transform 1 0 2760 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1644511149
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_14_36
timestamp 1644511149
transform 1 0 4416 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_14_48
timestamp 1644511149
transform 1 0 5520 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_14_58
timestamp 1644511149
transform 1 0 6440 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_62
timestamp 1644511149
transform 1 0 6808 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_14_73
timestamp 1644511149
transform 1 0 7820 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_14_80
timestamp 1644511149
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_101
timestamp 1644511149
transform 1 0 10396 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_14_119
timestamp 1644511149
transform 1 0 12052 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_123
timestamp 1644511149
transform 1 0 12420 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_14_131
timestamp 1644511149
transform 1 0 13156 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_145
timestamp 1644511149
transform 1 0 14444 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_14_163
timestamp 1644511149
transform 1 0 16100 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_14_173
timestamp 1644511149
transform 1 0 17020 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_14_180
timestamp 1644511149
transform 1 0 17664 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_14_190
timestamp 1644511149
transform 1 0 18584 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1644511149
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_14_204
timestamp 1644511149
transform 1 0 19872 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_14_224
timestamp 1644511149
transform 1 0 21712 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_228
timestamp 1644511149
transform 1 0 22080 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_14_235
timestamp 1644511149
transform 1 0 22724 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_14_243
timestamp 1644511149
transform 1 0 23460 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_257
timestamp 1644511149
transform 1 0 24748 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_14_264
timestamp 1644511149
transform 1 0 25392 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_14_278
timestamp 1644511149
transform 1 0 26680 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_14_292
timestamp 1644511149
transform 1 0 27968 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_14_304
timestamp 1644511149
transform 1 0 29072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_14_315
timestamp 1644511149
transform 1 0 30084 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_14_322
timestamp 1644511149
transform 1 0 30728 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_14_329
timestamp 1644511149
transform 1 0 31372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_15_6
timestamp 1644511149
transform 1 0 1656 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_15_20
timestamp 1644511149
transform 1 0 2944 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_15_37
timestamp 1644511149
transform 1 0 4508 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_15_47
timestamp 1644511149
transform 1 0 5428 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_15_70
timestamp 1644511149
transform 1 0 7544 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_15_83
timestamp 1644511149
transform 1 0 8740 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_15_94
timestamp 1644511149
transform 1 0 9752 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_15_108
timestamp 1644511149
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_15_121
timestamp 1644511149
transform 1 0 12236 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_129
timestamp 1644511149
transform 1 0 12972 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_15_157
timestamp 1644511149
transform 1 0 15548 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_15_164
timestamp 1644511149
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_15_175
timestamp 1644511149
transform 1 0 17204 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_15_190
timestamp 1644511149
transform 1 0 18584 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_15_200
timestamp 1644511149
transform 1 0 19504 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_204
timestamp 1644511149
transform 1 0 19872 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_206
timestamp 1644511149
transform 1 0 20056 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_15_215
timestamp 1644511149
transform 1 0 20884 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_15_231
timestamp 1644511149
transform 1 0 22356 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_15_241
timestamp 1644511149
transform 1 0 23276 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_15_255
timestamp 1644511149
transform 1 0 24564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_15_275
timestamp 1644511149
transform 1 0 26404 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_15_284
timestamp 1644511149
transform 1 0 27232 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_15_304
timestamp 1644511149
transform 1 0 29072 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_15_318
timestamp 1644511149
transform 1 0 30360 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_16_19
timestamp 1644511149
transform 1 0 2852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_16_49
timestamp 1644511149
transform 1 0 5612 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_55
timestamp 1644511149
transform 1 0 6164 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_16_62
timestamp 1644511149
transform 1 0 6808 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_16_69
timestamp 1644511149
transform 1 0 7452 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_16_80
timestamp 1644511149
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_16_90
timestamp 1644511149
transform 1 0 9384 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_16_110
timestamp 1644511149
transform 1 0 11224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_114
timestamp 1644511149
transform 1 0 11592 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_137
timestamp 1644511149
transform 1 0 13708 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_16_185
timestamp 1644511149
transform 1 0 18124 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_16_192
timestamp 1644511149
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_16_201
timestamp 1644511149
transform 1 0 19596 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_217
timestamp 1644511149
transform 1 0 21068 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_16_223
timestamp 1644511149
transform 1 0 21620 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_16_243
timestamp 1644511149
transform 1 0 23460 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_16_269
timestamp 1644511149
transform 1 0 25852 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_297
timestamp 1644511149
transform 1 0 28428 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_16_302
timestamp 1644511149
transform 1 0 28888 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1644511149
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_311
timestamp 1644511149
transform 1 0 29716 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_16_329
timestamp 1644511149
transform 1 0 31372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_17_13
timestamp 1644511149
transform 1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_17
timestamp 1644511149
transform 1 0 2668 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_19
timestamp 1644511149
transform 1 0 2852 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_35
timestamp 1644511149
transform 1 0 4324 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_17_45
timestamp 1644511149
transform 1 0 5244 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_17_52
timestamp 1644511149
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_17_70
timestamp 1644511149
transform 1 0 7544 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_17_78
timestamp 1644511149
transform 1 0 8280 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_17_95
timestamp 1644511149
transform 1 0 9844 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_17_107
timestamp 1644511149
transform 1 0 10948 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_17_119
timestamp 1644511149
transform 1 0 12052 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_127
timestamp 1644511149
transform 1 0 12788 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_17_133
timestamp 1644511149
transform 1 0 13340 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_17_143
timestamp 1644511149
transform 1 0 14260 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_17_156
timestamp 1644511149
transform 1 0 15456 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_17_164
timestamp 1644511149
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_17_175
timestamp 1644511149
transform 1 0 17204 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_179
timestamp 1644511149
transform 1 0 17572 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_17_198
timestamp 1644511149
transform 1 0 19320 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_17_209
timestamp 1644511149
transform 1 0 20332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_17_219
timestamp 1644511149
transform 1 0 21252 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_17_233
timestamp 1644511149
transform 1 0 22540 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_17_247
timestamp 1644511149
transform 1 0 23828 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_17_257
timestamp 1644511149
transform 1 0 24748 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_277
timestamp 1644511149
transform 1 0 26588 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_17_289
timestamp 1644511149
transform 1 0 27692 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_17_296
timestamp 1644511149
transform 1 0 28336 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_17_316
timestamp 1644511149
transform 1 0 30176 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_17_328
timestamp 1644511149
transform 1 0 31280 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_332
timestamp 1644511149
transform 1 0 31648 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_18_9
timestamp 1644511149
transform 1 0 1932 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_18_21
timestamp 1644511149
transform 1 0 3036 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_25
timestamp 1644511149
transform 1 0 3404 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_18_39
timestamp 1644511149
transform 1 0 4692 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_18_49
timestamp 1644511149
transform 1 0 5612 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_18_71
timestamp 1644511149
transform 1 0 7636 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_18_80
timestamp 1644511149
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_18_89
timestamp 1644511149
transform 1 0 9292 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_18_101
timestamp 1644511149
transform 1 0 10396 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_18_115
timestamp 1644511149
transform 1 0 11684 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_123
timestamp 1644511149
transform 1 0 12420 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_18_130
timestamp 1644511149
transform 1 0 13064 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1644511149
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_18_161
timestamp 1644511149
transform 1 0 15916 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_169
timestamp 1644511149
transform 1 0 16652 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_193
timestamp 1644511149
transform 1 0 18860 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_199
timestamp 1644511149
transform 1 0 19412 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1644511149
transform 1 0 20700 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_18_230
timestamp 1644511149
transform 1 0 22264 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_18_242
timestamp 1644511149
transform 1 0 23368 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1644511149
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_18_261
timestamp 1644511149
transform 1 0 25116 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_18_271
timestamp 1644511149
transform 1 0 26036 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_275
timestamp 1644511149
transform 1 0 26404 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_18_294
timestamp 1644511149
transform 1 0 28152 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_18_304
timestamp 1644511149
transform 1 0 29072 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_18_317
timestamp 1644511149
transform 1 0 30268 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_18_327
timestamp 1644511149
transform 1 0 31188 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_331
timestamp 1644511149
transform 1 0 31556 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_19_13
timestamp 1644511149
transform 1 0 2300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_19_33
timestamp 1644511149
transform 1 0 4140 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_37
timestamp 1644511149
transform 1 0 4508 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_19_46
timestamp 1644511149
transform 1 0 5336 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1644511149
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_19_66
timestamp 1644511149
transform 1 0 7176 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_19_79
timestamp 1644511149
transform 1 0 8372 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_19_86
timestamp 1644511149
transform 1 0 9016 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_19_100
timestamp 1644511149
transform 1 0 10304 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_19_108
timestamp 1644511149
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_115
timestamp 1644511149
transform 1 0 11684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_19_132
timestamp 1644511149
transform 1 0 13248 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_19_145
timestamp 1644511149
transform 1 0 14444 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_153
timestamp 1644511149
transform 1 0 15180 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_19_158
timestamp 1644511149
transform 1 0 15640 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1644511149
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_19_177
timestamp 1644511149
transform 1 0 17388 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_185
timestamp 1644511149
transform 1 0 18124 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_19_194
timestamp 1644511149
transform 1 0 18952 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_19_214
timestamp 1644511149
transform 1 0 20792 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1644511149
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_19_229
timestamp 1644511149
transform 1 0 22172 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_233
timestamp 1644511149
transform 1 0 22540 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_19_238
timestamp 1644511149
transform 1 0 23000 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_19_256
timestamp 1644511149
transform 1 0 24656 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_19_265
timestamp 1644511149
transform 1 0 25484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_19_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_277
timestamp 1644511149
transform 1 0 26588 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_285
timestamp 1644511149
transform 1 0 27324 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_19_292
timestamp 1644511149
transform 1 0 27968 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_300
timestamp 1644511149
transform 1 0 28704 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_19_310
timestamp 1644511149
transform 1 0 29624 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_314
timestamp 1644511149
transform 1 0 29992 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_316
timestamp 1644511149
transform 1 0 30176 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_19_325
timestamp 1644511149
transform 1 0 31004 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_20_19
timestamp 1644511149
transform 1 0 2852 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_20_33
timestamp 1644511149
transform 1 0 4140 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_20_62
timestamp 1644511149
transform 1 0 6808 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_70
timestamp 1644511149
transform 1 0 7544 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_20_80
timestamp 1644511149
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_20_101
timestamp 1644511149
transform 1 0 10396 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_20_115
timestamp 1644511149
transform 1 0 11684 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_123
timestamp 1644511149
transform 1 0 12420 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_20_129
timestamp 1644511149
transform 1 0 12972 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_20_136
timestamp 1644511149
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_20_157
timestamp 1644511149
transform 1 0 15548 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_20_181
timestamp 1644511149
transform 1 0 17756 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_185
timestamp 1644511149
transform 1 0 18124 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_187
timestamp 1644511149
transform 1 0 18308 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_20_192
timestamp 1644511149
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_20_217
timestamp 1644511149
transform 1 0 21068 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_20_225
timestamp 1644511149
transform 1 0 21804 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_229
timestamp 1644511149
transform 1 0 22172 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_231
timestamp 1644511149
transform 1 0 22356 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_20_236
timestamp 1644511149
transform 1 0 22816 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_240
timestamp 1644511149
transform 1 0 23184 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_20_248
timestamp 1644511149
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_20_263
timestamp 1644511149
transform 1 0 25300 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_267
timestamp 1644511149
transform 1 0 25668 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_20_274
timestamp 1644511149
transform 1 0 26312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_20_294
timestamp 1644511149
transform 1 0 28152 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_20_303
timestamp 1644511149
transform 1 0 28980 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_20_329
timestamp 1644511149
transform 1 0 31372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_21_7
timestamp 1644511149
transform 1 0 1748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_21_19
timestamp 1644511149
transform 1 0 2852 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_21_29
timestamp 1644511149
transform 1 0 3772 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_21_36
timestamp 1644511149
transform 1 0 4416 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_21_49
timestamp 1644511149
transform 1 0 5612 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_53
timestamp 1644511149
transform 1 0 5980 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_21_67
timestamp 1644511149
transform 1 0 7268 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_21_76
timestamp 1644511149
transform 1 0 8096 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_21_84
timestamp 1644511149
transform 1 0 8832 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_88
timestamp 1644511149
transform 1 0 9200 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_21_95
timestamp 1644511149
transform 1 0 9844 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_21_103
timestamp 1644511149
transform 1 0 10580 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_21_119
timestamp 1644511149
transform 1 0 12052 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_21_127
timestamp 1644511149
transform 1 0 12788 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_21_135
timestamp 1644511149
transform 1 0 13524 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_21_144
timestamp 1644511149
transform 1 0 14352 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_21_164
timestamp 1644511149
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_21_174
timestamp 1644511149
transform 1 0 17112 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_21_186
timestamp 1644511149
transform 1 0 18216 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_190
timestamp 1644511149
transform 1 0 18584 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_21_195
timestamp 1644511149
transform 1 0 19044 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_21_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_21_215
timestamp 1644511149
transform 1 0 20884 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_21_230
timestamp 1644511149
transform 1 0 22264 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_238
timestamp 1644511149
transform 1 0 23000 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_21_256
timestamp 1644511149
transform 1 0 24656 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_21_264
timestamp 1644511149
transform 1 0 25392 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_21_276
timestamp 1644511149
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_21_289
timestamp 1644511149
transform 1 0 27692 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_21_311
timestamp 1644511149
transform 1 0 29716 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_315
timestamp 1644511149
transform 1 0 30084 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_21_324
timestamp 1644511149
transform 1 0 30912 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_332
timestamp 1644511149
transform 1 0 31648 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_22_13
timestamp 1644511149
transform 1 0 2300 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_22_23
timestamp 1644511149
transform 1 0 3220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_22_37
timestamp 1644511149
transform 1 0 4508 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_22_59
timestamp 1644511149
transform 1 0 6532 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_22_67
timestamp 1644511149
transform 1 0 7268 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_22_80
timestamp 1644511149
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_101
timestamp 1644511149
transform 1 0 10396 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_22_118
timestamp 1644511149
transform 1 0 11960 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_22_130
timestamp 1644511149
transform 1 0 13064 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1644511149
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_22_144
timestamp 1644511149
transform 1 0 14352 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_22_152
timestamp 1644511149
transform 1 0 15088 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_22_160
timestamp 1644511149
transform 1 0 15824 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_22_169
timestamp 1644511149
transform 1 0 16652 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_173
timestamp 1644511149
transform 1 0 17020 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_22_178
timestamp 1644511149
transform 1 0 17480 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_22_188
timestamp 1644511149
transform 1 0 18400 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_22_201
timestamp 1644511149
transform 1 0 19596 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_22_231
timestamp 1644511149
transform 1 0 22356 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_239
timestamp 1644511149
transform 1 0 23092 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_22_248
timestamp 1644511149
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_22_273
timestamp 1644511149
transform 1 0 26220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_22_283
timestamp 1644511149
transform 1 0 27140 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_22_291
timestamp 1644511149
transform 1 0 27876 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_22_304
timestamp 1644511149
transform 1 0 29072 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_22_315
timestamp 1644511149
transform 1 0 30084 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_319
timestamp 1644511149
transform 1 0 30452 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_22_328
timestamp 1644511149
transform 1 0 31280 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_332
timestamp 1644511149
transform 1 0 31648 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_23_12
timestamp 1644511149
transform 1 0 2208 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_23_34
timestamp 1644511149
transform 1 0 4232 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_23_48
timestamp 1644511149
transform 1 0 5520 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_23_68
timestamp 1644511149
transform 1 0 7360 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_23_78
timestamp 1644511149
transform 1 0 8280 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_23_85
timestamp 1644511149
transform 1 0 8924 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_23_95
timestamp 1644511149
transform 1 0 9844 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_99
timestamp 1644511149
transform 1 0 10212 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_23_108
timestamp 1644511149
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_117
timestamp 1644511149
transform 1 0 11868 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_23_124
timestamp 1644511149
transform 1 0 12512 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_23_136
timestamp 1644511149
transform 1 0 13616 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_23_143
timestamp 1644511149
transform 1 0 14260 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_23_153
timestamp 1644511149
transform 1 0 15180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_23_163
timestamp 1644511149
transform 1 0 16100 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_23_178
timestamp 1644511149
transform 1 0 17480 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1644511149
transform 1 0 17848 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_23_199
timestamp 1644511149
transform 1 0 19412 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_23_219
timestamp 1644511149
transform 1 0 21252 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_23_241
timestamp 1644511149
transform 1 0 23276 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_23_257
timestamp 1644511149
transform 1 0 24748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_23_269
timestamp 1644511149
transform 1 0 25852 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_23_276
timestamp 1644511149
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_23_287
timestamp 1644511149
transform 1 0 27508 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_295
timestamp 1644511149
transform 1 0 28244 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_23_302
timestamp 1644511149
transform 1 0 28888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_23_313
timestamp 1644511149
transform 1 0 29900 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_24_19
timestamp 1644511149
transform 1 0 2852 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_24_38
timestamp 1644511149
transform 1 0 4600 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_24_45
timestamp 1644511149
transform 1 0 5244 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_24_58
timestamp 1644511149
transform 1 0 6440 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_24_80
timestamp 1644511149
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_24_95
timestamp 1644511149
transform 1 0 9844 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_24_115
timestamp 1644511149
transform 1 0 11684 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_119
timestamp 1644511149
transform 1 0 12052 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_24_136
timestamp 1644511149
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_24_149
timestamp 1644511149
transform 1 0 14812 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_24_163
timestamp 1644511149
transform 1 0 16100 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_171
timestamp 1644511149
transform 1 0 16836 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_24_178
timestamp 1644511149
transform 1 0 17480 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_182
timestamp 1644511149
transform 1 0 17848 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_24_192
timestamp 1644511149
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_24_202
timestamp 1644511149
transform 1 0 19688 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_24_226
timestamp 1644511149
transform 1 0 21896 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_24_238
timestamp 1644511149
transform 1 0 23000 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_24_248
timestamp 1644511149
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_24_261
timestamp 1644511149
transform 1 0 25116 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_24_271
timestamp 1644511149
transform 1 0 26036 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_24_279
timestamp 1644511149
transform 1 0 26772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_24_290
timestamp 1644511149
transform 1 0 27784 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_24_304
timestamp 1644511149
transform 1 0 29072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_311
timestamp 1644511149
transform 1 0 29716 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_24_328
timestamp 1644511149
transform 1 0 31280 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_332
timestamp 1644511149
transform 1 0 31648 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_25_7
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_25_20
timestamp 1644511149
transform 1 0 2944 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_25_32
timestamp 1644511149
transform 1 0 4048 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_25_52
timestamp 1644511149
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_25_65
timestamp 1644511149
transform 1 0 7084 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_25_89
timestamp 1644511149
transform 1 0 9292 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_25_103
timestamp 1644511149
transform 1 0 10580 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_25_133
timestamp 1644511149
transform 1 0 13340 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_139
timestamp 1644511149
transform 1 0 13892 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_25_156
timestamp 1644511149
transform 1 0 15456 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_25_164
timestamp 1644511149
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_25_174
timestamp 1644511149
transform 1 0 17112 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1644511149
transform 1 0 17848 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_25_189
timestamp 1644511149
transform 1 0 18492 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_25_197
timestamp 1644511149
transform 1 0 19228 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_201
timestamp 1644511149
transform 1 0 19596 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_25_208
timestamp 1644511149
transform 1 0 20240 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_25_219
timestamp 1644511149
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_227
timestamp 1644511149
transform 1 0 21988 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_25_234
timestamp 1644511149
transform 1 0 22632 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_238
timestamp 1644511149
transform 1 0 23000 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_25_255
timestamp 1644511149
transform 1 0 24564 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_25_263
timestamp 1644511149
transform 1 0 25300 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_267
timestamp 1644511149
transform 1 0 25668 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_25_276
timestamp 1644511149
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_25_289
timestamp 1644511149
transform 1 0 27692 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_295
timestamp 1644511149
transform 1 0 28244 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_25_312
timestamp 1644511149
transform 1 0 29808 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_320
timestamp 1644511149
transform 1 0 30544 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_25_327
timestamp 1644511149
transform 1 0 31188 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_331
timestamp 1644511149
transform 1 0 31556 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_26_12
timestamp 1644511149
transform 1 0 2208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_26_22
timestamp 1644511149
transform 1 0 3128 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1644511149
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_26_38
timestamp 1644511149
transform 1 0 4600 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_26_51
timestamp 1644511149
transform 1 0 5796 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_55
timestamp 1644511149
transform 1 0 6164 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_26_73
timestamp 1644511149
transform 1 0 7820 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_26_80
timestamp 1644511149
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_26_101
timestamp 1644511149
transform 1 0 10396 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_105
timestamp 1644511149
transform 1 0 10764 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_26_113
timestamp 1644511149
transform 1 0 11500 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_26_127
timestamp 1644511149
transform 1 0 12788 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_131
timestamp 1644511149
transform 1 0 13156 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_26_136
timestamp 1644511149
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_26_178
timestamp 1644511149
transform 1 0 17480 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_26_187
timestamp 1644511149
transform 1 0 18308 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_199
timestamp 1644511149
transform 1 0 19412 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_26_208
timestamp 1644511149
transform 1 0 20240 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_212
timestamp 1644511149
transform 1 0 20608 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_26_234
timestamp 1644511149
transform 1 0 22632 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_26_248
timestamp 1644511149
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_26_260
timestamp 1644511149
transform 1 0 25024 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_264
timestamp 1644511149
transform 1 0 25392 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_26_282
timestamp 1644511149
transform 1 0 27048 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_286
timestamp 1644511149
transform 1 0 27416 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_26_294
timestamp 1644511149
transform 1 0 28152 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_26_304
timestamp 1644511149
transform 1 0 29072 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_26_317
timestamp 1644511149
transform 1 0 30268 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_26_327
timestamp 1644511149
transform 1 0 31188 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_331
timestamp 1644511149
transform 1 0 31556 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1644511149
transform 1 0 1748 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_27_24
timestamp 1644511149
transform 1 0 3312 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_28
timestamp 1644511149
transform 1 0 3680 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_27_39
timestamp 1644511149
transform 1 0 4692 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_27_52
timestamp 1644511149
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_61
timestamp 1644511149
transform 1 0 6716 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_27_70
timestamp 1644511149
transform 1 0 7544 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_27_79
timestamp 1644511149
transform 1 0 8372 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_87
timestamp 1644511149
transform 1 0 9108 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_27_94
timestamp 1644511149
transform 1 0 9752 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_27_106
timestamp 1644511149
transform 1 0 10856 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1644511149
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_115
timestamp 1644511149
transform 1 0 11684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_27_124
timestamp 1644511149
transform 1 0 12512 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_142
timestamp 1644511149
transform 1 0 14168 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_27_158
timestamp 1644511149
transform 1 0 15640 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1644511149
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_27_189
timestamp 1644511149
transform 1 0 18492 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_27_209
timestamp 1644511149
transform 1 0 20332 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_27_220
timestamp 1644511149
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_27_241
timestamp 1644511149
transform 1 0 23276 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_27_248
timestamp 1644511149
transform 1 0 23920 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_27_259
timestamp 1644511149
transform 1 0 24932 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_267
timestamp 1644511149
transform 1 0 25668 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_27_276
timestamp 1644511149
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_27_289
timestamp 1644511149
transform 1 0 27692 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_27_300
timestamp 1644511149
transform 1 0 28704 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_27_308
timestamp 1644511149
transform 1 0 29440 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_27_328
timestamp 1644511149
transform 1 0 31280 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_332
timestamp 1644511149
transform 1 0 31648 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_5
timestamp 1644511149
transform 1 0 1564 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_28_24
timestamp 1644511149
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_28_34
timestamp 1644511149
transform 1 0 4232 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_28_56
timestamp 1644511149
transform 1 0 6256 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_60
timestamp 1644511149
transform 1 0 6624 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_62
timestamp 1644511149
transform 1 0 6808 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_28_70
timestamp 1644511149
transform 1 0 7544 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_28_80
timestamp 1644511149
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_89
timestamp 1644511149
transform 1 0 9292 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_28_106
timestamp 1644511149
transform 1 0 10856 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_28_127
timestamp 1644511149
transform 1 0 12788 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_28_135
timestamp 1644511149
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_28_157
timestamp 1644511149
transform 1 0 15548 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_161
timestamp 1644511149
transform 1 0 15916 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_163
timestamp 1644511149
transform 1 0 16100 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_28_173
timestamp 1644511149
transform 1 0 17020 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_28_186
timestamp 1644511149
transform 1 0 18216 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1644511149
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_28_204
timestamp 1644511149
transform 1 0 19872 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_212
timestamp 1644511149
transform 1 0 20608 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_220
timestamp 1644511149
transform 1 0 21344 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_225
timestamp 1644511149
transform 1 0 21804 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_229
timestamp 1644511149
transform 1 0 22172 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_28_239
timestamp 1644511149
transform 1 0 23092 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_243
timestamp 1644511149
transform 1 0 23460 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_28_248
timestamp 1644511149
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_255
timestamp 1644511149
transform 1 0 24564 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_28_264
timestamp 1644511149
transform 1 0 25392 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_28_272
timestamp 1644511149
transform 1 0 26128 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1644511149
transform 1 0 26496 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_28_284
timestamp 1644511149
transform 1 0 27232 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_288
timestamp 1644511149
transform 1 0 27600 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_28_298
timestamp 1644511149
transform 1 0 28520 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_306
timestamp 1644511149
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_28_329
timestamp 1644511149
transform 1 0 31372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_29_7
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_29_14
timestamp 1644511149
transform 1 0 2392 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_29_38
timestamp 1644511149
transform 1 0 4600 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_29_48
timestamp 1644511149
transform 1 0 5520 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_29_68
timestamp 1644511149
transform 1 0 7360 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_29_101
timestamp 1644511149
transform 1 0 10396 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_29_108
timestamp 1644511149
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_29_119
timestamp 1644511149
transform 1 0 12052 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_123
timestamp 1644511149
transform 1 0 12420 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_29_140
timestamp 1644511149
transform 1 0 13984 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_29_150
timestamp 1644511149
transform 1 0 14904 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_154
timestamp 1644511149
transform 1 0 15272 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_29_164
timestamp 1644511149
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_29_175
timestamp 1644511149
transform 1 0 17204 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_29_195
timestamp 1644511149
transform 1 0 19044 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_29_203
timestamp 1644511149
transform 1 0 19780 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_29_215
timestamp 1644511149
transform 1 0 20884 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_29_232
timestamp 1644511149
transform 1 0 22448 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_236
timestamp 1644511149
transform 1 0 22816 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_238
timestamp 1644511149
transform 1 0 23000 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_29_245
timestamp 1644511149
transform 1 0 23644 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_29_255
timestamp 1644511149
transform 1 0 24564 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_29_275
timestamp 1644511149
transform 1 0 26404 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_29_284
timestamp 1644511149
transform 1 0 27232 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_29_304
timestamp 1644511149
transform 1 0 29072 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_29_311
timestamp 1644511149
transform 1 0 29716 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_29_323
timestamp 1644511149
transform 1 0 30820 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_331
timestamp 1644511149
transform 1 0 31556 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_5
timestamp 1644511149
transform 1 0 1564 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_30_12
timestamp 1644511149
transform 1 0 2208 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_16
timestamp 1644511149
transform 1 0 2576 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_30_24
timestamp 1644511149
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_30_37
timestamp 1644511149
transform 1 0 4508 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_30_46
timestamp 1644511149
transform 1 0 5336 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_30_66
timestamp 1644511149
transform 1 0 7176 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_30_79
timestamp 1644511149
transform 1 0 8372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_137
timestamp 1644511149
transform 1 0 13708 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_30_145
timestamp 1644511149
transform 1 0 14444 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_30_157
timestamp 1644511149
transform 1 0 15548 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_165
timestamp 1644511149
transform 1 0 16284 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_30_177
timestamp 1644511149
transform 1 0 17388 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_30_187
timestamp 1644511149
transform 1 0 18308 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_201
timestamp 1644511149
transform 1 0 19596 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_30_229
timestamp 1644511149
transform 1 0 22172 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_30_240
timestamp 1644511149
transform 1 0 23184 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_30_248
timestamp 1644511149
transform 1 0 23920 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_30_261
timestamp 1644511149
transform 1 0 25116 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_30_285
timestamp 1644511149
transform 1 0 27324 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_30_296
timestamp 1644511149
transform 1 0 28336 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_30_304
timestamp 1644511149
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_30_329
timestamp 1644511149
transform 1 0 31372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_31_13
timestamp 1644511149
transform 1 0 2300 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_17
timestamp 1644511149
transform 1 0 2668 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_31_24
timestamp 1644511149
transform 1 0 3312 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_28
timestamp 1644511149
transform 1 0 3680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_31_46
timestamp 1644511149
transform 1 0 5336 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1644511149
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_31_63
timestamp 1644511149
transform 1 0 6900 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_67
timestamp 1644511149
transform 1 0 7268 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_31_76
timestamp 1644511149
transform 1 0 8096 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_80
timestamp 1644511149
transform 1 0 8464 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_31_85
timestamp 1644511149
transform 1 0 8924 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_31_95
timestamp 1644511149
transform 1 0 9844 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_31_107
timestamp 1644511149
transform 1 0 10948 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_31_120
timestamp 1644511149
transform 1 0 12144 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_128
timestamp 1644511149
transform 1 0 12880 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_31_133
timestamp 1644511149
transform 1 0 13340 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_31_153
timestamp 1644511149
transform 1 0 15180 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_31_163
timestamp 1644511149
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_31_185
timestamp 1644511149
transform 1 0 18124 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_31_196
timestamp 1644511149
transform 1 0 19136 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_31_206
timestamp 1644511149
transform 1 0 20056 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_31_218
timestamp 1644511149
transform 1 0 21160 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1644511149
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_31_229
timestamp 1644511149
transform 1 0 22172 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_31_249
timestamp 1644511149
transform 1 0 24012 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_31_258
timestamp 1644511149
transform 1 0 24840 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_31_272
timestamp 1644511149
transform 1 0 26128 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_31_289
timestamp 1644511149
transform 1 0 27692 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_31_298
timestamp 1644511149
transform 1 0 28520 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_31_310
timestamp 1644511149
transform 1 0 29624 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_31_317
timestamp 1644511149
transform 1 0 30268 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_31_329
timestamp 1644511149
transform 1 0 31372 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_32_6
timestamp 1644511149
transform 1 0 1656 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_32_18
timestamp 1644511149
transform 1 0 2760 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1644511149
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_32_33
timestamp 1644511149
transform 1 0 4140 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_32_47
timestamp 1644511149
transform 1 0 5428 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_55
timestamp 1644511149
transform 1 0 6164 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_32_63
timestamp 1644511149
transform 1 0 6900 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_67
timestamp 1644511149
transform 1 0 7268 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_32_71
timestamp 1644511149
transform 1 0 7636 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_75
timestamp 1644511149
transform 1 0 8004 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_32_80
timestamp 1644511149
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_32_89
timestamp 1644511149
transform 1 0 9292 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_93
timestamp 1644511149
transform 1 0 9660 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_32_100
timestamp 1644511149
transform 1 0 10304 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_104
timestamp 1644511149
transform 1 0 10672 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_32_110
timestamp 1644511149
transform 1 0 11224 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_32_119
timestamp 1644511149
transform 1 0 12052 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_32_127
timestamp 1644511149
transform 1 0 12788 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_32_135
timestamp 1644511149
transform 1 0 13524 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_32_145
timestamp 1644511149
transform 1 0 14444 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_153
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_32_164
timestamp 1644511149
transform 1 0 16192 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_32_178
timestamp 1644511149
transform 1 0 17480 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_32_192
timestamp 1644511149
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_201
timestamp 1644511149
transform 1 0 19596 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_32_219
timestamp 1644511149
transform 1 0 21252 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_223
timestamp 1644511149
transform 1 0 21620 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_225
timestamp 1644511149
transform 1 0 21804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_32_233
timestamp 1644511149
transform 1 0 22540 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_237
timestamp 1644511149
transform 1 0 22908 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_239
timestamp 1644511149
transform 1 0 23092 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_32_248
timestamp 1644511149
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_32_264
timestamp 1644511149
transform 1 0 25392 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_32_284
timestamp 1644511149
transform 1 0 27232 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_32_297
timestamp 1644511149
transform 1 0 28428 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_32_304
timestamp 1644511149
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_32_312
timestamp 1644511149
transform 1 0 29808 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_32_324
timestamp 1644511149
transform 1 0 30912 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_332
timestamp 1644511149
transform 1 0 31648 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_33_19
timestamp 1644511149
transform 1 0 2852 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_33_31
timestamp 1644511149
transform 1 0 3956 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_33_38
timestamp 1644511149
transform 1 0 4600 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_33_52
timestamp 1644511149
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_59
timestamp 1644511149
transform 1 0 6532 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_33_67
timestamp 1644511149
transform 1 0 7268 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_33_87
timestamp 1644511149
transform 1 0 9108 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_33_94
timestamp 1644511149
transform 1 0 9752 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_98
timestamp 1644511149
transform 1 0 10120 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_33_107
timestamp 1644511149
transform 1 0 10948 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_33_129
timestamp 1644511149
transform 1 0 12972 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_33_139
timestamp 1644511149
transform 1 0 13892 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_33_151
timestamp 1644511149
transform 1 0 14996 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_33_164
timestamp 1644511149
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_33_172
timestamp 1644511149
transform 1 0 16928 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_33_184
timestamp 1644511149
transform 1 0 18032 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_33_196
timestamp 1644511149
transform 1 0 19136 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_33_210
timestamp 1644511149
transform 1 0 20424 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_33_219
timestamp 1644511149
transform 1 0 21252 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1644511149
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_33_233
timestamp 1644511149
transform 1 0 22540 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_237
timestamp 1644511149
transform 1 0 22908 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_239
timestamp 1644511149
transform 1 0 23092 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_33_247
timestamp 1644511149
transform 1 0 23828 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_33_267
timestamp 1644511149
transform 1 0 25668 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_33_276
timestamp 1644511149
transform 1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_283
timestamp 1644511149
transform 1 0 27140 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_33_290
timestamp 1644511149
transform 1 0 27784 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_33_303
timestamp 1644511149
transform 1 0 28980 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_307
timestamp 1644511149
transform 1 0 29348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_33_316
timestamp 1644511149
transform 1 0 30176 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_33_327
timestamp 1644511149
transform 1 0 31188 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_331
timestamp 1644511149
transform 1 0 31556 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_34_7
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_34_19
timestamp 1644511149
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_34_45
timestamp 1644511149
transform 1 0 5244 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_69
timestamp 1644511149
transform 1 0 7452 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_34_80
timestamp 1644511149
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_34_111
timestamp 1644511149
transform 1 0 11316 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_34_121
timestamp 1644511149
transform 1 0 12236 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_125
timestamp 1644511149
transform 1 0 12604 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_127
timestamp 1644511149
transform 1 0 12788 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_34_136
timestamp 1644511149
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_34_147
timestamp 1644511149
transform 1 0 14628 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_151
timestamp 1644511149
transform 1 0 14996 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_34_161
timestamp 1644511149
transform 1 0 15916 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_169
timestamp 1644511149
transform 1 0 16652 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_34_178
timestamp 1644511149
transform 1 0 17480 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_34_186
timestamp 1644511149
transform 1 0 18216 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1644511149
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_34_204
timestamp 1644511149
transform 1 0 19872 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_34_228
timestamp 1644511149
transform 1 0 22080 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_34_248
timestamp 1644511149
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_34_258
timestamp 1644511149
transform 1 0 24840 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_34_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_34_285
timestamp 1644511149
transform 1 0 27324 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_34_292
timestamp 1644511149
transform 1 0 27968 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_34_303
timestamp 1644511149
transform 1 0 28980 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_34_329
timestamp 1644511149
transform 1 0 31372 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_7
timestamp 1644511149
transform 1 0 1748 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_35_14
timestamp 1644511149
transform 1 0 2392 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_18
timestamp 1644511149
transform 1 0 2760 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_20
timestamp 1644511149
transform 1 0 2944 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_35_31
timestamp 1644511149
transform 1 0 3956 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_35_52
timestamp 1644511149
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_35_68
timestamp 1644511149
transform 1 0 7360 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_35_79
timestamp 1644511149
transform 1 0 8372 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_35_86
timestamp 1644511149
transform 1 0 9016 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_35_99
timestamp 1644511149
transform 1 0 10212 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_103
timestamp 1644511149
transform 1 0 10580 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_35_108
timestamp 1644511149
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_35_123
timestamp 1644511149
transform 1 0 12420 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_35_131
timestamp 1644511149
transform 1 0 13156 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_35_151
timestamp 1644511149
transform 1 0 14996 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_35_160
timestamp 1644511149
transform 1 0 15824 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_35_176
timestamp 1644511149
transform 1 0 17296 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_180
timestamp 1644511149
transform 1 0 17664 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_182
timestamp 1644511149
transform 1 0 17848 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_35_199
timestamp 1644511149
transform 1 0 19412 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_35_213
timestamp 1644511149
transform 1 0 20700 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_35_220
timestamp 1644511149
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_35_231
timestamp 1644511149
transform 1 0 22356 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_35_246
timestamp 1644511149
transform 1 0 23736 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_35_256
timestamp 1644511149
transform 1 0 24656 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_260
timestamp 1644511149
transform 1 0 25024 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_35_266
timestamp 1644511149
transform 1 0 25576 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_35_276
timestamp 1644511149
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_283
timestamp 1644511149
transform 1 0 27140 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_35_293
timestamp 1644511149
transform 1 0 28060 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_35_308
timestamp 1644511149
transform 1 0 29440 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_35_318
timestamp 1644511149
transform 1 0 30360 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_35_328
timestamp 1644511149
transform 1 0 31280 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_332
timestamp 1644511149
transform 1 0 31648 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_36_19
timestamp 1644511149
transform 1 0 2852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_36_49
timestamp 1644511149
transform 1 0 5612 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_55
timestamp 1644511149
transform 1 0 6164 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_36_63
timestamp 1644511149
transform 1 0 6900 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_71
timestamp 1644511149
transform 1 0 7636 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_36_78
timestamp 1644511149
transform 1 0 8280 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1644511149
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_36_90
timestamp 1644511149
transform 1 0 9384 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_36_100
timestamp 1644511149
transform 1 0 10304 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_36_107
timestamp 1644511149
transform 1 0 10948 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_36_132
timestamp 1644511149
transform 1 0 13248 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_36_144
timestamp 1644511149
transform 1 0 14352 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_36_164
timestamp 1644511149
transform 1 0 16192 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_36_180
timestamp 1644511149
transform 1 0 17664 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_36_192
timestamp 1644511149
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_36_205
timestamp 1644511149
transform 1 0 19964 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_209
timestamp 1644511149
transform 1 0 20332 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_36_230
timestamp 1644511149
transform 1 0 22264 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_36_243
timestamp 1644511149
transform 1 0 23460 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_36_262
timestamp 1644511149
transform 1 0 25208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_36_270
timestamp 1644511149
transform 1 0 25944 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_36_280
timestamp 1644511149
transform 1 0 26864 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_284
timestamp 1644511149
transform 1 0 27232 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_286
timestamp 1644511149
transform 1 0 27416 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_36_295
timestamp 1644511149
transform 1 0 28244 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_36_304
timestamp 1644511149
transform 1 0 29072 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_36_318
timestamp 1644511149
transform 1 0 30360 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_36_328
timestamp 1644511149
transform 1 0 31280 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_332
timestamp 1644511149
transform 1 0 31648 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_37_7
timestamp 1644511149
transform 1 0 1748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_11
timestamp 1644511149
transform 1 0 2116 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_37_35
timestamp 1644511149
transform 1 0 4324 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_37_45
timestamp 1644511149
transform 1 0 5244 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_37_52
timestamp 1644511149
transform 1 0 5888 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_37_63
timestamp 1644511149
transform 1 0 6900 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_37_78
timestamp 1644511149
transform 1 0 8280 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_86
timestamp 1644511149
transform 1 0 9016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_37_91
timestamp 1644511149
transform 1 0 9476 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_37_103
timestamp 1644511149
transform 1 0 10580 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_117
timestamp 1644511149
transform 1 0 11868 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_37_134
timestamp 1644511149
transform 1 0 13432 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_37_148
timestamp 1644511149
transform 1 0 14720 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_37_158
timestamp 1644511149
transform 1 0 15640 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1644511149
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_37_185
timestamp 1644511149
transform 1 0 18124 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_37_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_197
timestamp 1644511149
transform 1 0 19228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_37_214
timestamp 1644511149
transform 1 0 20792 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1644511149
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_37_232
timestamp 1644511149
transform 1 0 22448 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_37_245
timestamp 1644511149
transform 1 0 23644 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_253
timestamp 1644511149
transform 1 0 24380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_37_261
timestamp 1644511149
transform 1 0 25116 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_269
timestamp 1644511149
transform 1 0 25852 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_37_276
timestamp 1644511149
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_37_289
timestamp 1644511149
transform 1 0 27692 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_37_299
timestamp 1644511149
transform 1 0 28612 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_37_310
timestamp 1644511149
transform 1 0 29624 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_37_322
timestamp 1644511149
transform 1 0 30728 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_37_329
timestamp 1644511149
transform 1 0 31372 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_7
timestamp 1644511149
transform 1 0 1748 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_38_17
timestamp 1644511149
transform 1 0 2668 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_38_24
timestamp 1644511149
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_38_37
timestamp 1644511149
transform 1 0 4508 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_38_49
timestamp 1644511149
transform 1 0 5612 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_38_57
timestamp 1644511149
transform 1 0 6348 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_61
timestamp 1644511149
transform 1 0 6716 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_38_69
timestamp 1644511149
transform 1 0 7452 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_38_80
timestamp 1644511149
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_89
timestamp 1644511149
transform 1 0 9292 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_38_106
timestamp 1644511149
transform 1 0 10856 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_38_116
timestamp 1644511149
transform 1 0 11776 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_38_126
timestamp 1644511149
transform 1 0 12696 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_130
timestamp 1644511149
transform 1 0 13064 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_38_135
timestamp 1644511149
transform 1 0 13524 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_38_145
timestamp 1644511149
transform 1 0 14444 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_149
timestamp 1644511149
transform 1 0 14812 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_38_158
timestamp 1644511149
transform 1 0 15640 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_38_186
timestamp 1644511149
transform 1 0 18216 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1644511149
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_38_203
timestamp 1644511149
transform 1 0 19780 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_38_210
timestamp 1644511149
transform 1 0 20424 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_38_223
timestamp 1644511149
transform 1 0 21620 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_38_235
timestamp 1644511149
transform 1 0 22724 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_38_247
timestamp 1644511149
transform 1 0 23828 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1644511149
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_38_259
timestamp 1644511149
transform 1 0 24932 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_263
timestamp 1644511149
transform 1 0 25300 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_38_282
timestamp 1644511149
transform 1 0 27048 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_38_296
timestamp 1644511149
transform 1 0 28336 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_38_304
timestamp 1644511149
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_38_329
timestamp 1644511149
transform 1 0 31372 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_39_10
timestamp 1644511149
transform 1 0 2024 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_39_23
timestamp 1644511149
transform 1 0 3220 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_39_33
timestamp 1644511149
transform 1 0 4140 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_39_41
timestamp 1644511149
transform 1 0 4876 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_39_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_39_73
timestamp 1644511149
transform 1 0 7820 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_109
timestamp 1644511149
transform 1 0 11132 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_39_123
timestamp 1644511149
transform 1 0 12420 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_39_143
timestamp 1644511149
transform 1 0 14260 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_151
timestamp 1644511149
transform 1 0 14996 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_39_160
timestamp 1644511149
transform 1 0 15824 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_39_176
timestamp 1644511149
transform 1 0 17296 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_39_186
timestamp 1644511149
transform 1 0 18216 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_39_193
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_39_204
timestamp 1644511149
transform 1 0 19872 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_212
timestamp 1644511149
transform 1 0 20608 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_39_219
timestamp 1644511149
transform 1 0 21252 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_39_242
timestamp 1644511149
transform 1 0 23368 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_250
timestamp 1644511149
transform 1 0 24104 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_39_267
timestamp 1644511149
transform 1 0 25668 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_39_275
timestamp 1644511149
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_39_285
timestamp 1644511149
transform 1 0 27324 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_289
timestamp 1644511149
transform 1 0 27692 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_39_306
timestamp 1644511149
transform 1 0 29256 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_310
timestamp 1644511149
transform 1 0 29624 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_312
timestamp 1644511149
transform 1 0 29808 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_39_321
timestamp 1644511149
transform 1 0 30636 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_39_329
timestamp 1644511149
transform 1 0 31372 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_40_11
timestamp 1644511149
transform 1 0 2116 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_40_22
timestamp 1644511149
transform 1 0 3128 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1644511149
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_40_37
timestamp 1644511149
transform 1 0 4508 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_40_44
timestamp 1644511149
transform 1 0 5152 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_40_56
timestamp 1644511149
transform 1 0 6256 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_40_70
timestamp 1644511149
transform 1 0 7544 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_40_80
timestamp 1644511149
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_40_93
timestamp 1644511149
transform 1 0 9660 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_40_103
timestamp 1644511149
transform 1 0 10580 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_107
timestamp 1644511149
transform 1 0 10948 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_40_124
timestamp 1644511149
transform 1 0 12512 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_40_136
timestamp 1644511149
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_40_147
timestamp 1644511149
transform 1 0 14628 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_151
timestamp 1644511149
transform 1 0 14996 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_40_163
timestamp 1644511149
transform 1 0 16100 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_40_171
timestamp 1644511149
transform 1 0 16836 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_179
timestamp 1644511149
transform 1 0 17572 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_40_188
timestamp 1644511149
transform 1 0 18400 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_40_213
timestamp 1644511149
transform 1 0 20700 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_40_233
timestamp 1644511149
transform 1 0 22540 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_241
timestamp 1644511149
transform 1 0 23276 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_40_248
timestamp 1644511149
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_257
timestamp 1644511149
transform 1 0 24748 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_40_263
timestamp 1644511149
transform 1 0 25300 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_40_271
timestamp 1644511149
transform 1 0 26036 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_275
timestamp 1644511149
transform 1 0 26404 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_40_285
timestamp 1644511149
transform 1 0 27324 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_289
timestamp 1644511149
transform 1 0 27692 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_291
timestamp 1644511149
transform 1 0 27876 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_40_300
timestamp 1644511149
transform 1 0 28704 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_40_329
timestamp 1644511149
transform 1 0 31372 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_41_19
timestamp 1644511149
transform 1 0 2852 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_41_30
timestamp 1644511149
transform 1 0 3864 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_41_42
timestamp 1644511149
transform 1 0 4968 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_41_50
timestamp 1644511149
transform 1 0 5704 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_54
timestamp 1644511149
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_41_66
timestamp 1644511149
transform 1 0 7176 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_41_86
timestamp 1644511149
transform 1 0 9016 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_94
timestamp 1644511149
transform 1 0 9752 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_41_103
timestamp 1644511149
transform 1 0 10580 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_115
timestamp 1644511149
transform 1 0 11684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_129
timestamp 1644511149
transform 1 0 12972 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_41_140
timestamp 1644511149
transform 1 0 13984 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_41_160
timestamp 1644511149
transform 1 0 15824 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_41_178
timestamp 1644511149
transform 1 0 17480 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_41_206
timestamp 1644511149
transform 1 0 20056 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_41_216
timestamp 1644511149
transform 1 0 20976 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_41_230
timestamp 1644511149
transform 1 0 22264 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_234
timestamp 1644511149
transform 1 0 22632 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_41_252
timestamp 1644511149
transform 1 0 24288 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_41_268
timestamp 1644511149
transform 1 0 25760 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_41_276
timestamp 1644511149
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_41_289
timestamp 1644511149
transform 1 0 27692 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_41_303
timestamp 1644511149
transform 1 0 28980 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_41_317
timestamp 1644511149
transform 1 0 30268 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_41_327
timestamp 1644511149
transform 1 0 31188 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_331
timestamp 1644511149
transform 1 0 31556 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_5
timestamp 1644511149
transform 1 0 1564 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_42_10
timestamp 1644511149
transform 1 0 2024 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_42_24
timestamp 1644511149
transform 1 0 3312 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_42_38
timestamp 1644511149
transform 1 0 4600 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_42_48
timestamp 1644511149
transform 1 0 5520 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_52
timestamp 1644511149
transform 1 0 5888 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_42_61
timestamp 1644511149
transform 1 0 6716 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_69
timestamp 1644511149
transform 1 0 7452 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_42_73
timestamp 1644511149
transform 1 0 7820 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_42_80
timestamp 1644511149
transform 1 0 8464 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_42_89
timestamp 1644511149
transform 1 0 9292 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_42_101
timestamp 1644511149
transform 1 0 10396 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_42_111
timestamp 1644511149
transform 1 0 11316 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_115
timestamp 1644511149
transform 1 0 11684 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_42_136
timestamp 1644511149
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_42_146
timestamp 1644511149
transform 1 0 14536 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_42_156
timestamp 1644511149
transform 1 0 15456 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_42_165
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_169
timestamp 1644511149
transform 1 0 16652 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_42_187
timestamp 1644511149
transform 1 0 18308 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_42_203
timestamp 1644511149
transform 1 0 19780 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_42_210
timestamp 1644511149
transform 1 0 20424 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_42_230
timestamp 1644511149
transform 1 0 22264 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_42_243
timestamp 1644511149
transform 1 0 23460 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_42_270
timestamp 1644511149
transform 1 0 25944 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_42_290
timestamp 1644511149
transform 1 0 27784 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_42_302
timestamp 1644511149
transform 1 0 28888 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_306
timestamp 1644511149
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_313
timestamp 1644511149
transform 1 0 29900 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_42_323
timestamp 1644511149
transform 1 0 30820 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_331
timestamp 1644511149
transform 1 0 31556 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_5
timestamp 1644511149
transform 1 0 1564 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_43_12
timestamp 1644511149
transform 1 0 2208 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_43_28
timestamp 1644511149
transform 1 0 3680 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_43_48
timestamp 1644511149
transform 1 0 5520 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_43_61
timestamp 1644511149
transform 1 0 6716 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_43_102
timestamp 1644511149
transform 1 0 10488 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1644511149
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_43_123
timestamp 1644511149
transform 1 0 12420 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_43_143
timestamp 1644511149
transform 1 0 14260 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_43_151
timestamp 1644511149
transform 1 0 14996 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_159
timestamp 1644511149
transform 1 0 15732 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_43_164
timestamp 1644511149
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_43_177
timestamp 1644511149
transform 1 0 17388 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_185
timestamp 1644511149
transform 1 0 18124 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_43_193
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_43_205
timestamp 1644511149
transform 1 0 19964 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_213
timestamp 1644511149
transform 1 0 20700 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_43_220
timestamp 1644511149
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_227
timestamp 1644511149
transform 1 0 21988 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_43_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_43_246
timestamp 1644511149
transform 1 0 23736 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_43_256
timestamp 1644511149
transform 1 0 24656 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_43_268
timestamp 1644511149
transform 1 0 25760 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_43_276
timestamp 1644511149
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_43_287
timestamp 1644511149
transform 1 0 27508 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_43_297
timestamp 1644511149
transform 1 0 28428 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_301
timestamp 1644511149
transform 1 0 28796 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_303
timestamp 1644511149
transform 1 0 28980 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_43_312
timestamp 1644511149
transform 1 0 29808 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_43_324
timestamp 1644511149
transform 1 0 30912 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_332
timestamp 1644511149
transform 1 0 31648 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_44_7
timestamp 1644511149
transform 1 0 1748 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_11
timestamp 1644511149
transform 1 0 2116 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_44_22
timestamp 1644511149
transform 1 0 3128 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_26
timestamp 1644511149
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_44_33
timestamp 1644511149
transform 1 0 4140 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_44_45
timestamp 1644511149
transform 1 0 5244 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_49
timestamp 1644511149
transform 1 0 5612 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_44_54
timestamp 1644511149
transform 1 0 6072 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_44_71
timestamp 1644511149
transform 1 0 7636 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_75
timestamp 1644511149
transform 1 0 8004 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_44_80
timestamp 1644511149
transform 1 0 8464 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_44_92
timestamp 1644511149
transform 1 0 9568 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_44_99
timestamp 1644511149
transform 1 0 10212 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_103
timestamp 1644511149
transform 1 0 10580 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_44_113
timestamp 1644511149
transform 1 0 11500 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_44_125
timestamp 1644511149
transform 1 0 12604 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_44_136
timestamp 1644511149
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_44_149
timestamp 1644511149
transform 1 0 14812 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_44_159
timestamp 1644511149
transform 1 0 15732 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_163
timestamp 1644511149
transform 1 0 16100 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_44_170
timestamp 1644511149
transform 1 0 16744 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_44_180
timestamp 1644511149
transform 1 0 17664 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_44_190
timestamp 1644511149
transform 1 0 18584 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_194
timestamp 1644511149
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_44_205
timestamp 1644511149
transform 1 0 19964 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_213
timestamp 1644511149
transform 1 0 20700 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_44_223
timestamp 1644511149
transform 1 0 21620 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_44_237
timestamp 1644511149
transform 1 0 22908 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_44_248
timestamp 1644511149
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_44_261
timestamp 1644511149
transform 1 0 25116 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_265
timestamp 1644511149
transform 1 0 25484 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_267
timestamp 1644511149
transform 1 0 25668 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_44_276
timestamp 1644511149
transform 1 0 26496 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_280
timestamp 1644511149
transform 1 0 26864 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_282
timestamp 1644511149
transform 1 0 27048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_44_303
timestamp 1644511149
transform 1 0 28980 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_44_329
timestamp 1644511149
transform 1 0 31372 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_45_11
timestamp 1644511149
transform 1 0 2116 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_45_31
timestamp 1644511149
transform 1 0 3956 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_45_43
timestamp 1644511149
transform 1 0 5060 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_47
timestamp 1644511149
transform 1 0 5428 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_45_52
timestamp 1644511149
transform 1 0 5888 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_45_66
timestamp 1644511149
transform 1 0 7176 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_70
timestamp 1644511149
transform 1 0 7544 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_45_92
timestamp 1644511149
transform 1 0 9568 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_45_108
timestamp 1644511149
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_45_129
timestamp 1644511149
transform 1 0 12972 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_45_139
timestamp 1644511149
transform 1 0 13892 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_143
timestamp 1644511149
transform 1 0 14260 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_145
timestamp 1644511149
transform 1 0 14444 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_45_162
timestamp 1644511149
transform 1 0 16008 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1644511149
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_45_173
timestamp 1644511149
transform 1 0 17020 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_45_193
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_45_201
timestamp 1644511149
transform 1 0 19596 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_45_215
timestamp 1644511149
transform 1 0 20884 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_45_249
timestamp 1644511149
transform 1 0 24012 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_45_270
timestamp 1644511149
transform 1 0 25944 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_278
timestamp 1644511149
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_45_284
timestamp 1644511149
transform 1 0 27232 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_45_304
timestamp 1644511149
transform 1 0 29072 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_308
timestamp 1644511149
transform 1 0 29440 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_45_326
timestamp 1644511149
transform 1 0 31096 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_330
timestamp 1644511149
transform 1 0 31464 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_332
timestamp 1644511149
transform 1 0 31648 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_7
timestamp 1644511149
transform 1 0 1748 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_46_17
timestamp 1644511149
transform 1 0 2668 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_46_24
timestamp 1644511149
transform 1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_46_32
timestamp 1644511149
transform 1 0 4048 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_46_44
timestamp 1644511149
transform 1 0 5152 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_46_56
timestamp 1644511149
transform 1 0 6256 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_60
timestamp 1644511149
transform 1 0 6624 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_81
timestamp 1644511149
transform 1 0 8556 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_46_89
timestamp 1644511149
transform 1 0 9292 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_46_119
timestamp 1644511149
transform 1 0 12052 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_46_129
timestamp 1644511149
transform 1 0 12972 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_46_136
timestamp 1644511149
transform 1 0 13616 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_143
timestamp 1644511149
transform 1 0 14260 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_46_148
timestamp 1644511149
transform 1 0 14720 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_46_160
timestamp 1644511149
transform 1 0 15824 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_168
timestamp 1644511149
transform 1 0 16560 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_46_175
timestamp 1644511149
transform 1 0 17204 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_46_185
timestamp 1644511149
transform 1 0 18124 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_46_192
timestamp 1644511149
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_201
timestamp 1644511149
transform 1 0 19596 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_46_219
timestamp 1644511149
transform 1 0 21252 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_46_231
timestamp 1644511149
transform 1 0 22356 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_46_238
timestamp 1644511149
transform 1 0 23000 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_46_248
timestamp 1644511149
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_46_261
timestamp 1644511149
transform 1 0 25116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_46_281
timestamp 1644511149
transform 1 0 26956 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_285
timestamp 1644511149
transform 1 0 27324 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_287
timestamp 1644511149
transform 1 0 27508 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_46_304
timestamp 1644511149
transform 1 0 29072 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_46_315
timestamp 1644511149
transform 1 0 30084 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_46_325
timestamp 1644511149
transform 1 0 31004 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_47_19
timestamp 1644511149
transform 1 0 2852 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_47_45
timestamp 1644511149
transform 1 0 5244 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_47_52
timestamp 1644511149
transform 1 0 5888 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_47_62
timestamp 1644511149
transform 1 0 6808 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_47_72
timestamp 1644511149
transform 1 0 7728 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_47_92
timestamp 1644511149
transform 1 0 9568 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_100
timestamp 1644511149
transform 1 0 10304 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_47_108
timestamp 1644511149
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_47_121
timestamp 1644511149
transform 1 0 12236 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_47_130
timestamp 1644511149
transform 1 0 13064 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_134
timestamp 1644511149
transform 1 0 13432 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_47_141
timestamp 1644511149
transform 1 0 14076 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_47_149
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_157
timestamp 1644511149
transform 1 0 15548 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_47_164
timestamp 1644511149
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_171
timestamp 1644511149
transform 1 0 16836 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_47_176
timestamp 1644511149
transform 1 0 17296 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_47_186
timestamp 1644511149
transform 1 0 18216 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_47_197
timestamp 1644511149
transform 1 0 19228 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_201
timestamp 1644511149
transform 1 0 19596 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_203
timestamp 1644511149
transform 1 0 19780 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_47_210
timestamp 1644511149
transform 1 0 20424 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_47_220
timestamp 1644511149
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_47_241
timestamp 1644511149
transform 1 0 23276 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_249
timestamp 1644511149
transform 1 0 24012 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_47_266
timestamp 1644511149
transform 1 0 25576 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_47_276
timestamp 1644511149
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_47_289
timestamp 1644511149
transform 1 0 27692 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_47_299
timestamp 1644511149
transform 1 0 28612 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_47_309
timestamp 1644511149
transform 1 0 29532 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_317
timestamp 1644511149
transform 1 0 30268 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_47_324
timestamp 1644511149
transform 1 0 30912 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_332
timestamp 1644511149
transform 1 0 31648 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_5
timestamp 1644511149
transform 1 0 1564 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_48_12
timestamp 1644511149
transform 1 0 2208 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_48_22
timestamp 1644511149
transform 1 0 3128 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_26
timestamp 1644511149
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_48_37
timestamp 1644511149
transform 1 0 4508 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_48_57
timestamp 1644511149
transform 1 0 6348 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_61
timestamp 1644511149
transform 1 0 6716 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_48_68
timestamp 1644511149
transform 1 0 7360 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_48_80
timestamp 1644511149
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_48_91
timestamp 1644511149
transform 1 0 9476 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_48_105
timestamp 1644511149
transform 1 0 10764 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_48_119
timestamp 1644511149
transform 1 0 12052 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_48_131
timestamp 1644511149
transform 1 0 13156 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_145
timestamp 1644511149
transform 1 0 14444 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_48_163
timestamp 1644511149
transform 1 0 16100 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_167
timestamp 1644511149
transform 1 0 16468 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_48_172
timestamp 1644511149
transform 1 0 16928 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_48_192
timestamp 1644511149
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_48_205
timestamp 1644511149
transform 1 0 19964 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_48_216
timestamp 1644511149
transform 1 0 20976 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_48_223
timestamp 1644511149
transform 1 0 21620 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_48_231
timestamp 1644511149
transform 1 0 22356 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_48_245
timestamp 1644511149
transform 1 0 23644 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_249
timestamp 1644511149
transform 1 0 24012 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_48_257
timestamp 1644511149
transform 1 0 24748 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_261
timestamp 1644511149
transform 1 0 25116 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_48_266
timestamp 1644511149
transform 1 0 25576 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_48_274
timestamp 1644511149
transform 1 0 26312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_48_294
timestamp 1644511149
transform 1 0 28152 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_48_304
timestamp 1644511149
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_48_329
timestamp 1644511149
transform 1 0 31372 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_49_7
timestamp 1644511149
transform 1 0 1748 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_11
timestamp 1644511149
transform 1 0 2116 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_49_16
timestamp 1644511149
transform 1 0 2576 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_49_40
timestamp 1644511149
transform 1 0 4784 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_49_50
timestamp 1644511149
transform 1 0 5704 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_54
timestamp 1644511149
transform 1 0 6072 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_49_73
timestamp 1644511149
transform 1 0 7820 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_49_85
timestamp 1644511149
transform 1 0 8924 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_49_101
timestamp 1644511149
transform 1 0 10396 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_49_108
timestamp 1644511149
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_49_131
timestamp 1644511149
transform 1 0 13156 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_49_151
timestamp 1644511149
transform 1 0 14996 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_49_164
timestamp 1644511149
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_173
timestamp 1644511149
transform 1 0 17020 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_49_183
timestamp 1644511149
transform 1 0 17940 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_49_191
timestamp 1644511149
transform 1 0 18676 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_195
timestamp 1644511149
transform 1 0 19044 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_49_206
timestamp 1644511149
transform 1 0 20056 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_210
timestamp 1644511149
transform 1 0 20424 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_49_220
timestamp 1644511149
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_49_229
timestamp 1644511149
transform 1 0 22172 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_233
timestamp 1644511149
transform 1 0 22540 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_49_242
timestamp 1644511149
transform 1 0 23368 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_250
timestamp 1644511149
transform 1 0 24104 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_49_260
timestamp 1644511149
transform 1 0 25024 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_268
timestamp 1644511149
transform 1 0 25760 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_49_276
timestamp 1644511149
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_49_287
timestamp 1644511149
transform 1 0 27508 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_49_300
timestamp 1644511149
transform 1 0 28704 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_49_312
timestamp 1644511149
transform 1 0 29808 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_316
timestamp 1644511149
transform 1 0 30176 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_49_325
timestamp 1644511149
transform 1 0 31004 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_7
timestamp 1644511149
transform 1 0 1748 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_50_24
timestamp 1644511149
transform 1 0 3312 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_50_39
timestamp 1644511149
transform 1 0 4692 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_50_64
timestamp 1644511149
transform 1 0 6992 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_50_80
timestamp 1644511149
transform 1 0 8464 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_50_92
timestamp 1644511149
transform 1 0 9568 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_96
timestamp 1644511149
transform 1 0 9936 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_50_105
timestamp 1644511149
transform 1 0 10764 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_50_115
timestamp 1644511149
transform 1 0 11684 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_50_127
timestamp 1644511149
transform 1 0 12788 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_131
timestamp 1644511149
transform 1 0 13156 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_50_136
timestamp 1644511149
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_50_149
timestamp 1644511149
transform 1 0 14812 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_50_163
timestamp 1644511149
transform 1 0 16100 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_50_183
timestamp 1644511149
transform 1 0 17940 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_187
timestamp 1644511149
transform 1 0 18308 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_50_192
timestamp 1644511149
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_50_213
timestamp 1644511149
transform 1 0 20700 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_50_224
timestamp 1644511149
transform 1 0 21712 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_232
timestamp 1644511149
transform 1 0 22448 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_50_242
timestamp 1644511149
transform 1 0 23368 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_250
timestamp 1644511149
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_50_262
timestamp 1644511149
transform 1 0 25208 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_50_271
timestamp 1644511149
transform 1 0 26036 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_275
timestamp 1644511149
transform 1 0 26404 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_50_283
timestamp 1644511149
transform 1 0 27140 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_287
timestamp 1644511149
transform 1 0 27508 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_50_304
timestamp 1644511149
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_50_329
timestamp 1644511149
transform 1 0 31372 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_51_8
timestamp 1644511149
transform 1 0 1840 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_51_18
timestamp 1644511149
transform 1 0 2760 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_51_30
timestamp 1644511149
transform 1 0 3864 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_34
timestamp 1644511149
transform 1 0 4232 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_51_52
timestamp 1644511149
transform 1 0 5888 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_59
timestamp 1644511149
transform 1 0 6532 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_51_68
timestamp 1644511149
transform 1 0 7360 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_51_79
timestamp 1644511149
transform 1 0 8372 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_87
timestamp 1644511149
transform 1 0 9108 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_109
timestamp 1644511149
transform 1 0 11132 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_51_123
timestamp 1644511149
transform 1 0 12420 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_127
timestamp 1644511149
transform 1 0 12788 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_51_135
timestamp 1644511149
transform 1 0 13524 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_139
timestamp 1644511149
transform 1 0 13892 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_51_146
timestamp 1644511149
transform 1 0 14536 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_51_158
timestamp 1644511149
transform 1 0 15640 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1644511149
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_173
timestamp 1644511149
transform 1 0 17020 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_51_180
timestamp 1644511149
transform 1 0 17664 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_188
timestamp 1644511149
transform 1 0 18400 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_51_210
timestamp 1644511149
transform 1 0 20424 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_214
timestamp 1644511149
transform 1 0 20792 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_51_219
timestamp 1644511149
transform 1 0 21252 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_51_231
timestamp 1644511149
transform 1 0 22356 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_51_240
timestamp 1644511149
transform 1 0 23184 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_248
timestamp 1644511149
transform 1 0 23920 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_51_259
timestamp 1644511149
transform 1 0 24932 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_263
timestamp 1644511149
transform 1 0 25300 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_51_271
timestamp 1644511149
transform 1 0 26036 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_51_292
timestamp 1644511149
transform 1 0 27968 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_51_300
timestamp 1644511149
transform 1 0 28704 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_304
timestamp 1644511149
transform 1 0 29072 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_51_326
timestamp 1644511149
transform 1 0 31096 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_330
timestamp 1644511149
transform 1 0 31464 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_332
timestamp 1644511149
transform 1 0 31648 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_52_19
timestamp 1644511149
transform 1 0 2852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_52_37
timestamp 1644511149
transform 1 0 4508 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_52_51
timestamp 1644511149
transform 1 0 5796 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_55
timestamp 1644511149
transform 1 0 6164 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_52_61
timestamp 1644511149
transform 1 0 6716 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_52_75
timestamp 1644511149
transform 1 0 8004 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_52_93
timestamp 1644511149
transform 1 0 9660 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_99
timestamp 1644511149
transform 1 0 10212 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_52_116
timestamp 1644511149
transform 1 0 11776 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_52_136
timestamp 1644511149
transform 1 0 13616 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_52_148
timestamp 1644511149
transform 1 0 14720 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_152
timestamp 1644511149
transform 1 0 15088 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_154
timestamp 1644511149
transform 1 0 15272 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_52_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_52_173
timestamp 1644511149
transform 1 0 17020 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_177
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_52_186
timestamp 1644511149
transform 1 0 18216 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1644511149
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_201
timestamp 1644511149
transform 1 0 19596 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_52_207
timestamp 1644511149
transform 1 0 20148 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_211
timestamp 1644511149
transform 1 0 20516 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_213
timestamp 1644511149
transform 1 0 20700 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_52_218
timestamp 1644511149
transform 1 0 21160 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_222
timestamp 1644511149
transform 1 0 21528 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_224
timestamp 1644511149
transform 1 0 21712 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_52_241
timestamp 1644511149
transform 1 0 23276 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_52_248
timestamp 1644511149
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_52_261
timestamp 1644511149
transform 1 0 25116 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_52_272
timestamp 1644511149
transform 1 0 26128 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_52_292
timestamp 1644511149
transform 1 0 27968 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_296
timestamp 1644511149
transform 1 0 28336 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_52_304
timestamp 1644511149
transform 1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_52_329
timestamp 1644511149
transform 1 0 31372 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_7
timestamp 1644511149
transform 1 0 1748 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_53_16
timestamp 1644511149
transform 1 0 2576 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_53_28
timestamp 1644511149
transform 1 0 3680 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_32
timestamp 1644511149
transform 1 0 4048 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_53_50
timestamp 1644511149
transform 1 0 5704 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_54
timestamp 1644511149
transform 1 0 6072 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_61
timestamp 1644511149
transform 1 0 6716 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_53_84
timestamp 1644511149
transform 1 0 8832 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_88
timestamp 1644511149
transform 1 0 9200 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_53_92
timestamp 1644511149
transform 1 0 9568 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_53_106
timestamp 1644511149
transform 1 0 10856 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1644511149
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_53_119
timestamp 1644511149
transform 1 0 12052 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_53_127
timestamp 1644511149
transform 1 0 12788 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_53_155
timestamp 1644511149
transform 1 0 15364 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_53_163
timestamp 1644511149
transform 1 0 16100 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1644511149
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_53_173
timestamp 1644511149
transform 1 0 17020 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_177
timestamp 1644511149
transform 1 0 17388 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_53_186
timestamp 1644511149
transform 1 0 18216 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_53_200
timestamp 1644511149
transform 1 0 19504 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_53_208
timestamp 1644511149
transform 1 0 20240 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_53_218
timestamp 1644511149
transform 1 0 21160 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1644511149
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_227
timestamp 1644511149
transform 1 0 21988 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_53_234
timestamp 1644511149
transform 1 0 22632 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_53_241
timestamp 1644511149
transform 1 0 23276 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_53_251
timestamp 1644511149
transform 1 0 24196 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_255
timestamp 1644511149
transform 1 0 24564 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_257
timestamp 1644511149
transform 1 0 24748 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_53_264
timestamp 1644511149
transform 1 0 25392 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_53_276
timestamp 1644511149
transform 1 0 26496 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_53_291
timestamp 1644511149
transform 1 0 27876 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_53_315
timestamp 1644511149
transform 1 0 30084 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_53_327
timestamp 1644511149
transform 1 0 31188 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_331
timestamp 1644511149
transform 1 0 31556 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_54_20
timestamp 1644511149
transform 1 0 2944 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_33
timestamp 1644511149
transform 1 0 4140 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_54_42
timestamp 1644511149
transform 1 0 4968 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_46
timestamp 1644511149
transform 1 0 5336 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_54_51
timestamp 1644511149
transform 1 0 5796 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_54_62
timestamp 1644511149
transform 1 0 6808 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_54_69
timestamp 1644511149
transform 1 0 7452 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_54_80
timestamp 1644511149
transform 1 0 8464 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_54_90
timestamp 1644511149
transform 1 0 9384 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_54_110
timestamp 1644511149
transform 1 0 11224 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_114
timestamp 1644511149
transform 1 0 11592 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_116
timestamp 1644511149
transform 1 0 11776 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_54_120
timestamp 1644511149
transform 1 0 12144 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_54_129
timestamp 1644511149
transform 1 0 12972 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_54_136
timestamp 1644511149
transform 1 0 13616 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_54_148
timestamp 1644511149
transform 1 0 14720 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_152
timestamp 1644511149
transform 1 0 15088 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_54_169
timestamp 1644511149
transform 1 0 16652 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_193
timestamp 1644511149
transform 1 0 18860 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_54_205
timestamp 1644511149
transform 1 0 19964 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_54_225
timestamp 1644511149
transform 1 0 21804 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_54_245
timestamp 1644511149
transform 1 0 23644 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_249
timestamp 1644511149
transform 1 0 24012 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_54_269
timestamp 1644511149
transform 1 0 25852 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_54_281
timestamp 1644511149
transform 1 0 26956 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_289
timestamp 1644511149
transform 1 0 27692 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_54_294
timestamp 1644511149
transform 1 0 28152 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_54_304
timestamp 1644511149
transform 1 0 29072 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_54_317
timestamp 1644511149
transform 1 0 30268 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_54_329
timestamp 1644511149
transform 1 0 31372 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_11
timestamp 1644511149
transform 1 0 2116 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_13
timestamp 1644511149
transform 1 0 2300 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_55_20
timestamp 1644511149
transform 1 0 2944 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_55_31
timestamp 1644511149
transform 1 0 3956 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_55_41
timestamp 1644511149
transform 1 0 4876 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_55_52
timestamp 1644511149
transform 1 0 5888 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_55_68
timestamp 1644511149
transform 1 0 7360 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_76
timestamp 1644511149
transform 1 0 8096 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_55_85
timestamp 1644511149
transform 1 0 8924 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_55_97
timestamp 1644511149
transform 1 0 10028 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_55_107
timestamp 1644511149
transform 1 0 10948 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_55_121
timestamp 1644511149
transform 1 0 12236 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_55_133
timestamp 1644511149
transform 1 0 13340 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_55_148
timestamp 1644511149
transform 1 0 14720 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_152
timestamp 1644511149
transform 1 0 15088 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_55_162
timestamp 1644511149
transform 1 0 16008 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1644511149
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_55_175
timestamp 1644511149
transform 1 0 17204 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_55_187
timestamp 1644511149
transform 1 0 18308 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_191
timestamp 1644511149
transform 1 0 18676 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_193
timestamp 1644511149
transform 1 0 18860 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_55_202
timestamp 1644511149
transform 1 0 19688 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_210
timestamp 1644511149
transform 1 0 20424 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_55_216
timestamp 1644511149
transform 1 0 20976 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_55_231
timestamp 1644511149
transform 1 0 22356 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_239
timestamp 1644511149
transform 1 0 23092 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_55_246
timestamp 1644511149
transform 1 0 23736 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_55_254
timestamp 1644511149
transform 1 0 24472 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_258
timestamp 1644511149
transform 1 0 24840 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_55_266
timestamp 1644511149
transform 1 0 25576 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_55_274
timestamp 1644511149
transform 1 0 26312 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_278
timestamp 1644511149
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_55_291
timestamp 1644511149
transform 1 0 27876 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_295
timestamp 1644511149
transform 1 0 28244 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_55_302
timestamp 1644511149
transform 1 0 28888 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_55_309
timestamp 1644511149
transform 1 0 29532 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_55_329
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_5
timestamp 1644511149
transform 1 0 1564 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_56_10
timestamp 1644511149
transform 1 0 2024 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_56_20
timestamp 1644511149
transform 1 0 2944 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_56_37
timestamp 1644511149
transform 1 0 4508 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_56_52
timestamp 1644511149
transform 1 0 5888 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_56
timestamp 1644511149
transform 1 0 6256 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_56_66
timestamp 1644511149
transform 1 0 7176 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_56_78
timestamp 1644511149
transform 1 0 8280 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_82
timestamp 1644511149
transform 1 0 8648 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_56_95
timestamp 1644511149
transform 1 0 9844 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_99
timestamp 1644511149
transform 1 0 10212 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_56_106
timestamp 1644511149
transform 1 0 10856 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_110
timestamp 1644511149
transform 1 0 11224 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_56_116
timestamp 1644511149
transform 1 0 11776 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_56_128
timestamp 1644511149
transform 1 0 12880 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_56_136
timestamp 1644511149
transform 1 0 13616 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_56_150
timestamp 1644511149
transform 1 0 14904 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_154
timestamp 1644511149
transform 1 0 15272 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_56_162
timestamp 1644511149
transform 1 0 16008 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_166
timestamp 1644511149
transform 1 0 16376 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_56_171
timestamp 1644511149
transform 1 0 16836 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_56_184
timestamp 1644511149
transform 1 0 18032 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_56_192
timestamp 1644511149
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_56_213
timestamp 1644511149
transform 1 0 20700 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_56_225
timestamp 1644511149
transform 1 0 21804 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_56_236
timestamp 1644511149
transform 1 0 22816 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_56_244
timestamp 1644511149
transform 1 0 23552 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_56_260
timestamp 1644511149
transform 1 0 25024 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_56_272
timestamp 1644511149
transform 1 0 26128 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_56_292
timestamp 1644511149
transform 1 0 27968 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_296
timestamp 1644511149
transform 1 0 28336 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_56_304
timestamp 1644511149
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_313
timestamp 1644511149
transform 1 0 29900 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_56_321
timestamp 1644511149
transform 1 0 30636 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_56_329
timestamp 1644511149
transform 1 0 31372 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_57_19
timestamp 1644511149
transform 1 0 2852 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_57_31
timestamp 1644511149
transform 1 0 3956 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_35
timestamp 1644511149
transform 1 0 4324 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_57_52
timestamp 1644511149
transform 1 0 5888 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_57_65
timestamp 1644511149
transform 1 0 7084 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_57_74
timestamp 1644511149
transform 1 0 7912 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_57_87
timestamp 1644511149
transform 1 0 9108 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_57_107
timestamp 1644511149
transform 1 0 10948 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_57_120
timestamp 1644511149
transform 1 0 12144 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_124
timestamp 1644511149
transform 1 0 12512 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_57_141
timestamp 1644511149
transform 1 0 14076 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_57_153
timestamp 1644511149
transform 1 0 15180 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_157
timestamp 1644511149
transform 1 0 15548 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_57_164
timestamp 1644511149
transform 1 0 16192 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_57_178
timestamp 1644511149
transform 1 0 17480 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_57_188
timestamp 1644511149
transform 1 0 18400 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_57_202
timestamp 1644511149
transform 1 0 19688 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_206
timestamp 1644511149
transform 1 0 20056 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_57_212
timestamp 1644511149
transform 1 0 20608 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_57_220
timestamp 1644511149
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_57_229
timestamp 1644511149
transform 1 0 22172 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_57_249
timestamp 1644511149
transform 1 0 24012 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_57_269
timestamp 1644511149
transform 1 0 25852 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_57_276
timestamp 1644511149
transform 1 0 26496 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_57_304
timestamp 1644511149
transform 1 0 29072 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_57_329
timestamp 1644511149
transform 1 0 31372 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_5
timestamp 1644511149
transform 1 0 1564 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_58_12
timestamp 1644511149
transform 1 0 2208 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_58_24
timestamp 1644511149
transform 1 0 3312 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_58_32
timestamp 1644511149
transform 1 0 4048 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_58_46
timestamp 1644511149
transform 1 0 5336 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_58_56
timestamp 1644511149
transform 1 0 6256 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_60
timestamp 1644511149
transform 1 0 6624 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_58_68
timestamp 1644511149
transform 1 0 7360 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_58_78
timestamp 1644511149
transform 1 0 8280 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_82
timestamp 1644511149
transform 1 0 8648 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_58_90
timestamp 1644511149
transform 1 0 9384 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_94
timestamp 1644511149
transform 1 0 9752 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_58_102
timestamp 1644511149
transform 1 0 10488 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_58_122
timestamp 1644511149
transform 1 0 12328 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_58_129
timestamp 1644511149
transform 1 0 12972 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_58_136
timestamp 1644511149
transform 1 0 13616 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_58_147
timestamp 1644511149
transform 1 0 14628 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_151
timestamp 1644511149
transform 1 0 14996 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_58_168
timestamp 1644511149
transform 1 0 16560 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_58_185
timestamp 1644511149
transform 1 0 18124 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_58_192
timestamp 1644511149
transform 1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_58_201
timestamp 1644511149
transform 1 0 19596 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_58_208
timestamp 1644511149
transform 1 0 20240 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_58_228
timestamp 1644511149
transform 1 0 22080 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_58_237
timestamp 1644511149
transform 1 0 22908 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_58_248
timestamp 1644511149
transform 1 0 23920 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_58_263
timestamp 1644511149
transform 1 0 25300 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_58_273
timestamp 1644511149
transform 1 0 26220 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_58_285
timestamp 1644511149
transform 1 0 27324 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_289
timestamp 1644511149
transform 1 0 27692 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_58_294
timestamp 1644511149
transform 1 0 28152 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_58_304
timestamp 1644511149
transform 1 0 29072 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_58_329
timestamp 1644511149
transform 1 0 31372 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_59_19
timestamp 1644511149
transform 1 0 2852 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_59
timestamp 1644511149
transform 1 0 6532 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_59_66
timestamp 1644511149
transform 1 0 7176 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_59_76
timestamp 1644511149
transform 1 0 8096 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_80
timestamp 1644511149
transform 1 0 8464 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_82
timestamp 1644511149
transform 1 0 8648 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_59_91
timestamp 1644511149
transform 1 0 9476 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_95
timestamp 1644511149
transform 1 0 9844 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_97
timestamp 1644511149
transform 1 0 10028 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_59_101
timestamp 1644511149
transform 1 0 10396 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_59_108
timestamp 1644511149
transform 1 0 11040 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_59_117
timestamp 1644511149
transform 1 0 11868 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_121
timestamp 1644511149
transform 1 0 12236 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_123
timestamp 1644511149
transform 1 0 12420 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_59_127
timestamp 1644511149
transform 1 0 12788 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_59_147
timestamp 1644511149
transform 1 0 14628 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_59_164
timestamp 1644511149
transform 1 0 16192 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_59_187
timestamp 1644511149
transform 1 0 18308 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_59_207
timestamp 1644511149
transform 1 0 20148 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_59_215
timestamp 1644511149
transform 1 0 20884 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_59_230
timestamp 1644511149
transform 1 0 22264 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_59_237
timestamp 1644511149
transform 1 0 22908 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_59_249
timestamp 1644511149
transform 1 0 24012 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_253
timestamp 1644511149
transform 1 0 24380 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_59_261
timestamp 1644511149
transform 1 0 25116 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_59_270
timestamp 1644511149
transform 1 0 25944 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_278
timestamp 1644511149
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_59_289
timestamp 1644511149
transform 1 0 27692 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_59_311
timestamp 1644511149
transform 1 0 29716 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_315
timestamp 1644511149
transform 1 0 30084 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_59_325
timestamp 1644511149
transform 1 0 31004 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_7
timestamp 1644511149
transform 1 0 1748 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_60_14
timestamp 1644511149
transform 1 0 2392 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_60_24
timestamp 1644511149
transform 1 0 3312 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_61
timestamp 1644511149
transform 1 0 6716 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_60_79
timestamp 1644511149
transform 1 0 8372 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_60_93
timestamp 1644511149
transform 1 0 9660 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_60_103
timestamp 1644511149
transform 1 0 10580 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_107
timestamp 1644511149
transform 1 0 10948 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_60_111
timestamp 1644511149
transform 1 0 11316 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_60_119
timestamp 1644511149
transform 1 0 12052 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_127
timestamp 1644511149
transform 1 0 12788 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_60_132
timestamp 1644511149
transform 1 0 13248 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_60_149
timestamp 1644511149
transform 1 0 14812 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_60_161
timestamp 1644511149
transform 1 0 15916 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_60_170
timestamp 1644511149
transform 1 0 16744 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_174
timestamp 1644511149
transform 1 0 17112 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_176
timestamp 1644511149
transform 1 0 17296 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_60_181
timestamp 1644511149
transform 1 0 17756 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_185
timestamp 1644511149
transform 1 0 18124 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_60_192
timestamp 1644511149
transform 1 0 18768 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_60_214
timestamp 1644511149
transform 1 0 20792 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_60_224
timestamp 1644511149
transform 1 0 21712 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_60_245
timestamp 1644511149
transform 1 0 23644 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_249
timestamp 1644511149
transform 1 0 24012 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_60_269
timestamp 1644511149
transform 1 0 25852 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_273
timestamp 1644511149
transform 1 0 26220 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_60_290
timestamp 1644511149
transform 1 0 27784 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_60_304
timestamp 1644511149
transform 1 0 29072 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_60_317
timestamp 1644511149
transform 1 0 30268 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_60_327
timestamp 1644511149
transform 1 0 31188 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_331
timestamp 1644511149
transform 1 0 31556 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_7 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1748 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_61_25
timestamp 1644511149
transform 1 0 3404 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_61_45
timestamp 1644511149
transform 1 0 5244 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_61_52
timestamp 1644511149
transform 1 0 5888 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_61_73
timestamp 1644511149
transform 1 0 7820 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_61_102
timestamp 1644511149
transform 1 0 10488 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_110
timestamp 1644511149
transform 1 0 11224 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_61_120
timestamp 1644511149
transform 1 0 12144 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_128
timestamp 1644511149
transform 1 0 12880 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_61_135
timestamp 1644511149
transform 1 0 13524 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_139
timestamp 1644511149
transform 1 0 13892 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_61_143
timestamp 1644511149
transform 1 0 14260 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_61_150
timestamp 1644511149
transform 1 0 14904 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_61_160
timestamp 1644511149
transform 1 0 15824 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_61_173
timestamp 1644511149
transform 1 0 17020 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_61_180
timestamp 1644511149
transform 1 0 17664 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_184
timestamp 1644511149
transform 1 0 18032 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_61_190
timestamp 1644511149
transform 1 0 18584 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_198
timestamp 1644511149
transform 1 0 19320 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_61_220
timestamp 1644511149
transform 1 0 21344 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_227
timestamp 1644511149
transform 1 0 21988 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_61_231
timestamp 1644511149
transform 1 0 22356 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_61_241
timestamp 1644511149
transform 1 0 23276 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_61_248
timestamp 1644511149
transform 1 0 23920 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_61_264
timestamp 1644511149
transform 1 0 25392 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_268
timestamp 1644511149
transform 1 0 25760 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_61_276
timestamp 1644511149
transform 1 0 26496 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_61_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_61_301
timestamp 1644511149
transform 1 0 28796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_61_315
timestamp 1644511149
transform 1 0 30084 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_61_327
timestamp 1644511149
transform 1 0 31188 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_331
timestamp 1644511149
transform 1 0 31556 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_7
timestamp 1644511149
transform 1 0 1748 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_62_14
timestamp 1644511149
transform 1 0 2392 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_62_24
timestamp 1644511149
transform 1 0 3312 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_45
timestamp 1644511149
transform 1 0 5244 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_57
timestamp 1644511149
transform 1 0 6348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_62_66
timestamp 1644511149
transform 1 0 7176 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_62_78
timestamp 1644511149
transform 1 0 8280 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_82
timestamp 1644511149
transform 1 0 8648 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_62_91
timestamp 1644511149
transform 1 0 9476 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_62_111
timestamp 1644511149
transform 1 0 11316 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_62_122
timestamp 1644511149
transform 1 0 12328 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_130
timestamp 1644511149
transform 1 0 13064 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_62_136
timestamp 1644511149
transform 1 0 13616 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_145
timestamp 1644511149
transform 1 0 14444 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_62_151
timestamp 1644511149
transform 1 0 14996 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_62_159
timestamp 1644511149
transform 1 0 15732 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_167
timestamp 1644511149
transform 1 0 16468 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_62_175
timestamp 1644511149
transform 1 0 17204 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_62_182
timestamp 1644511149
transform 1 0 17848 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_186
timestamp 1644511149
transform 1 0 18216 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_188
timestamp 1644511149
transform 1 0 18400 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_62_192
timestamp 1644511149
transform 1 0 18768 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_62_203
timestamp 1644511149
transform 1 0 19780 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_62_210
timestamp 1644511149
transform 1 0 20424 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_62_231
timestamp 1644511149
transform 1 0 22356 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_235
timestamp 1644511149
transform 1 0 22724 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_62_237
timestamp 1644511149
transform 1 0 22908 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_62_244
timestamp 1644511149
transform 1 0 23552 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_257
timestamp 1644511149
transform 1 0 24748 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_62_267
timestamp 1644511149
transform 1 0 25668 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_62_277
timestamp 1644511149
transform 1 0 26588 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_62_284
timestamp 1644511149
transform 1 0 27232 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_62_304
timestamp 1644511149
transform 1 0 29072 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_62_313
timestamp 1644511149
transform 1 0 29900 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_62_325
timestamp 1644511149
transform 1 0 31004 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_63_19
timestamp 1644511149
transform 1 0 2852 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_23
timestamp 1644511149
transform 1 0 3220 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_63_45
timestamp 1644511149
transform 1 0 5244 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_53
timestamp 1644511149
transform 1 0 5980 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_63_65
timestamp 1644511149
transform 1 0 7084 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_63_87
timestamp 1644511149
transform 1 0 9108 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_63_101
timestamp 1644511149
transform 1 0 10396 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_63_108
timestamp 1644511149
transform 1 0 11040 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_63_129
timestamp 1644511149
transform 1 0 12972 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_63_139
timestamp 1644511149
transform 1 0 13892 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_143
timestamp 1644511149
transform 1 0 14260 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_145
timestamp 1644511149
transform 1 0 14444 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_63_151
timestamp 1644511149
transform 1 0 14996 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_63_164
timestamp 1644511149
transform 1 0 16192 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_63_187
timestamp 1644511149
transform 1 0 18308 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_63_207
timestamp 1644511149
transform 1 0 20148 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_211
timestamp 1644511149
transform 1 0 20516 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_213
timestamp 1644511149
transform 1 0 20700 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_63_220
timestamp 1644511149
transform 1 0 21344 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_63_228
timestamp 1644511149
transform 1 0 22080 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_63_248
timestamp 1644511149
transform 1 0 23920 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_252
timestamp 1644511149
transform 1 0 24288 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_63_269
timestamp 1644511149
transform 1 0 25852 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_63_276
timestamp 1644511149
transform 1 0 26496 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_63_289
timestamp 1644511149
transform 1 0 27692 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_63_297
timestamp 1644511149
transform 1 0 28428 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_63_309
timestamp 1644511149
transform 1 0 29532 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_63_329
timestamp 1644511149
transform 1 0 31372 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_64_7
timestamp 1644511149
transform 1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_11
timestamp 1644511149
transform 1 0 2116 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_64_21
timestamp 1644511149
transform 1 0 3036 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_25
timestamp 1644511149
transform 1 0 3404 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_64_37
timestamp 1644511149
transform 1 0 4508 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_45
timestamp 1644511149
transform 1 0 5244 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_47
timestamp 1644511149
transform 1 0 5428 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_64_64
timestamp 1644511149
transform 1 0 6992 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_64_71
timestamp 1644511149
transform 1 0 7636 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_64_80
timestamp 1644511149
transform 1 0 8464 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_64_94
timestamp 1644511149
transform 1 0 9752 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_64_108
timestamp 1644511149
transform 1 0 11040 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_64_115
timestamp 1644511149
transform 1 0 11684 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_119
timestamp 1644511149
transform 1 0 12052 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_64_136
timestamp 1644511149
transform 1 0 13616 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_145
timestamp 1644511149
transform 1 0 14444 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_64_151
timestamp 1644511149
transform 1 0 14996 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_155
timestamp 1644511149
transform 1 0 15364 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_64_163
timestamp 1644511149
transform 1 0 16100 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_64_174
timestamp 1644511149
transform 1 0 17112 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_178
timestamp 1644511149
transform 1 0 17480 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_180
timestamp 1644511149
transform 1 0 17664 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_193
timestamp 1644511149
transform 1 0 18860 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_64_205
timestamp 1644511149
transform 1 0 19964 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_213
timestamp 1644511149
transform 1 0 20700 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_64_230
timestamp 1644511149
transform 1 0 22264 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_64_240
timestamp 1644511149
transform 1 0 23184 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_64_247
timestamp 1644511149
transform 1 0 23828 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_64_261
timestamp 1644511149
transform 1 0 25116 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_267
timestamp 1644511149
transform 1 0 25668 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_64_284
timestamp 1644511149
transform 1 0 27232 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_64_296
timestamp 1644511149
transform 1 0 28336 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_64_304
timestamp 1644511149
transform 1 0 29072 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_64_325
timestamp 1644511149
transform 1 0 31004 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_65_9
timestamp 1644511149
transform 1 0 1932 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_65_21
timestamp 1644511149
transform 1 0 3036 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_25
timestamp 1644511149
transform 1 0 3404 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_65_35
timestamp 1644511149
transform 1 0 4324 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_65_46
timestamp 1644511149
transform 1 0 5336 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_54
timestamp 1644511149
transform 1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_65_63
timestamp 1644511149
transform 1 0 6900 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_71
timestamp 1644511149
transform 1 0 7636 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_65_77
timestamp 1644511149
transform 1 0 8188 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_65_86
timestamp 1644511149
transform 1 0 9016 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_65_95
timestamp 1644511149
transform 1 0 9844 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_65_104
timestamp 1644511149
transform 1 0 10672 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_65_120
timestamp 1644511149
transform 1 0 12144 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_124
timestamp 1644511149
transform 1 0 12512 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_65_133
timestamp 1644511149
transform 1 0 13340 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_65_148
timestamp 1644511149
transform 1 0 14720 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_152
timestamp 1644511149
transform 1 0 15088 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_154
timestamp 1644511149
transform 1 0 15272 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_65_164
timestamp 1644511149
transform 1 0 16192 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_65_173
timestamp 1644511149
transform 1 0 17020 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_65_183
timestamp 1644511149
transform 1 0 17940 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_187
timestamp 1644511149
transform 1 0 18308 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_189
timestamp 1644511149
transform 1 0 18492 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_65_198
timestamp 1644511149
transform 1 0 19320 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_65_210
timestamp 1644511149
transform 1 0 20424 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_65_218
timestamp 1644511149
transform 1 0 21160 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_222
timestamp 1644511149
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_65_232
timestamp 1644511149
transform 1 0 22448 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_65_240
timestamp 1644511149
transform 1 0 23184 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_248
timestamp 1644511149
transform 1 0 23920 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_65_254
timestamp 1644511149
transform 1 0 24472 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_258
timestamp 1644511149
transform 1 0 24840 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_65_266
timestamp 1644511149
transform 1 0 25576 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_65_276
timestamp 1644511149
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_283
timestamp 1644511149
transform 1 0 27140 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_65_300
timestamp 1644511149
transform 1 0 28704 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_65_310
timestamp 1644511149
transform 1 0 29624 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_314
timestamp 1644511149
transform 1 0 29992 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_65_324
timestamp 1644511149
transform 1 0 30912 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_332
timestamp 1644511149
transform 1 0 31648 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_66_19
timestamp 1644511149
transform 1 0 2852 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_33
timestamp 1644511149
transform 1 0 4140 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_66_43
timestamp 1644511149
transform 1 0 5060 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_66_56
timestamp 1644511149
transform 1 0 6256 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_66_66
timestamp 1644511149
transform 1 0 7176 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_66_76
timestamp 1644511149
transform 1 0 8096 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_66_91
timestamp 1644511149
transform 1 0 9476 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_99
timestamp 1644511149
transform 1 0 10212 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_66_108
timestamp 1644511149
transform 1 0 11040 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_66_116
timestamp 1644511149
transform 1 0 11776 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_66_136
timestamp 1644511149
transform 1 0 13616 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_145
timestamp 1644511149
transform 1 0 14444 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_66_154
timestamp 1644511149
transform 1 0 15272 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_66_163
timestamp 1644511149
transform 1 0 16100 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_66_171
timestamp 1644511149
transform 1 0 16836 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_179
timestamp 1644511149
transform 1 0 17572 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_66_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_193
timestamp 1644511149
transform 1 0 18860 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_66_208
timestamp 1644511149
transform 1 0 20240 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_66_218
timestamp 1644511149
transform 1 0 21160 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_66_226
timestamp 1644511149
transform 1 0 21896 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_234
timestamp 1644511149
transform 1 0 22632 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_66_239
timestamp 1644511149
transform 1 0 23092 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_66_248
timestamp 1644511149
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_66_260
timestamp 1644511149
transform 1 0 25024 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_66_274
timestamp 1644511149
transform 1 0 26312 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_66_281
timestamp 1644511149
transform 1 0 26956 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_66_292
timestamp 1644511149
transform 1 0 27968 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_66_304
timestamp 1644511149
transform 1 0 29072 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_66_329
timestamp 1644511149
transform 1 0 31372 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_67_13
timestamp 1644511149
transform 1 0 2300 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_67_25
timestamp 1644511149
transform 1 0 3404 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_29
timestamp 1644511149
transform 1 0 3772 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_31
timestamp 1644511149
transform 1 0 3956 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_67_42
timestamp 1644511149
transform 1 0 4968 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_46
timestamp 1644511149
transform 1 0 5336 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_67_52
timestamp 1644511149
transform 1 0 5888 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_67_60
timestamp 1644511149
transform 1 0 6624 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_67_80
timestamp 1644511149
transform 1 0 8464 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_88
timestamp 1644511149
transform 1 0 9200 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_90
timestamp 1644511149
transform 1 0 9384 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_67_108
timestamp 1644511149
transform 1 0 11040 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_67_121
timestamp 1644511149
transform 1 0 12236 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_67_135
timestamp 1644511149
transform 1 0 13524 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_139
timestamp 1644511149
transform 1 0 13892 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_67_148
timestamp 1644511149
transform 1 0 14720 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_67_160
timestamp 1644511149
transform 1 0 15824 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_67_189
timestamp 1644511149
transform 1 0 18492 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_67_199
timestamp 1644511149
transform 1 0 19412 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_67_220
timestamp 1644511149
transform 1 0 21344 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_227
timestamp 1644511149
transform 1 0 21988 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_67_234
timestamp 1644511149
transform 1 0 22632 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_238
timestamp 1644511149
transform 1 0 23000 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_67_244
timestamp 1644511149
transform 1 0 23552 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_248
timestamp 1644511149
transform 1 0 23920 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_67_256
timestamp 1644511149
transform 1 0 24656 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_260
timestamp 1644511149
transform 1 0 25024 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_262
timestamp 1644511149
transform 1 0 25208 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_67_271
timestamp 1644511149
transform 1 0 26036 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1644511149
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_67_289
timestamp 1644511149
transform 1 0 27692 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_67_309
timestamp 1644511149
transform 1 0 29532 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_67_329
timestamp 1644511149
transform 1 0 31372 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_7
timestamp 1644511149
transform 1 0 1748 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_68_24
timestamp 1644511149
transform 1 0 3312 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_31
timestamp 1644511149
transform 1 0 3956 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_68_39
timestamp 1644511149
transform 1 0 4692 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_43
timestamp 1644511149
transform 1 0 5060 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_45
timestamp 1644511149
transform 1 0 5244 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_68_51
timestamp 1644511149
transform 1 0 5796 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_55
timestamp 1644511149
transform 1 0 6164 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_68_72
timestamp 1644511149
transform 1 0 7728 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_68_80
timestamp 1644511149
transform 1 0 8464 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_68_92
timestamp 1644511149
transform 1 0 9568 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_68_99
timestamp 1644511149
transform 1 0 10212 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_68_123
timestamp 1644511149
transform 1 0 12420 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_68_135
timestamp 1644511149
transform 1 0 13524 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_68_146
timestamp 1644511149
transform 1 0 14536 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_150
timestamp 1644511149
transform 1 0 14904 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_68_171
timestamp 1644511149
transform 1 0 16836 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_68_182
timestamp 1644511149
transform 1 0 17848 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_68_192
timestamp 1644511149
transform 1 0 18768 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_201
timestamp 1644511149
transform 1 0 19596 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_68_219
timestamp 1644511149
transform 1 0 21252 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_68_239
timestamp 1644511149
transform 1 0 23092 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_243
timestamp 1644511149
transform 1 0 23460 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_68_248
timestamp 1644511149
transform 1 0 23920 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_68_261
timestamp 1644511149
transform 1 0 25116 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_68_273
timestamp 1644511149
transform 1 0 26220 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_68_284
timestamp 1644511149
transform 1 0 27232 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_68_295
timestamp 1644511149
transform 1 0 28244 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_68_304
timestamp 1644511149
transform 1 0 29072 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_68_317
timestamp 1644511149
transform 1 0 30268 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_68_327
timestamp 1644511149
transform 1 0 31188 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_331
timestamp 1644511149
transform 1 0 31556 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_11
timestamp 1644511149
transform 1 0 2116 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_69_18
timestamp 1644511149
transform 1 0 2760 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_69_30
timestamp 1644511149
transform 1 0 3864 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_34
timestamp 1644511149
transform 1 0 4232 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_69_60
timestamp 1644511149
transform 1 0 6624 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_69_72
timestamp 1644511149
transform 1 0 7728 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_69_84
timestamp 1644511149
transform 1 0 8832 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_69_94
timestamp 1644511149
transform 1 0 9752 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_98
timestamp 1644511149
transform 1 0 10120 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_69_108
timestamp 1644511149
transform 1 0 11040 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_69_133
timestamp 1644511149
transform 1 0 13340 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_139
timestamp 1644511149
transform 1 0 13892 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_69_156
timestamp 1644511149
transform 1 0 15456 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_69_164
timestamp 1644511149
transform 1 0 16192 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_173
timestamp 1644511149
transform 1 0 17020 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_69_182
timestamp 1644511149
transform 1 0 17848 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_69_202
timestamp 1644511149
transform 1 0 19688 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_206
timestamp 1644511149
transform 1 0 20056 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_69_217
timestamp 1644511149
transform 1 0 21068 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_221
timestamp 1644511149
transform 1 0 21436 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1644511149
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_69_233
timestamp 1644511149
transform 1 0 22540 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_69_245
timestamp 1644511149
transform 1 0 23644 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_69_252
timestamp 1644511149
transform 1 0 24288 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_69_276
timestamp 1644511149
transform 1 0 26496 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_283
timestamp 1644511149
transform 1 0 27140 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_69_291
timestamp 1644511149
transform 1 0 27876 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_69_301
timestamp 1644511149
transform 1 0 28796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_69_315
timestamp 1644511149
transform 1 0 30084 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_69_325
timestamp 1644511149
transform 1 0 31004 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_70_5
timestamp 1644511149
transform 1 0 1564 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_70_12
timestamp 1644511149
transform 1 0 2208 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_70_22
timestamp 1644511149
transform 1 0 3128 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_26
timestamp 1644511149
transform 1 0 3496 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_33
timestamp 1644511149
transform 1 0 4140 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_70_45
timestamp 1644511149
transform 1 0 5244 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_70_56
timestamp 1644511149
transform 1 0 6256 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_60
timestamp 1644511149
transform 1 0 6624 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_70_68
timestamp 1644511149
transform 1 0 7360 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_70_80
timestamp 1644511149
transform 1 0 8464 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_70_95
timestamp 1644511149
transform 1 0 9844 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_99
timestamp 1644511149
transform 1 0 10212 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_70_107
timestamp 1644511149
transform 1 0 10948 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_115
timestamp 1644511149
transform 1 0 11684 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_70_123
timestamp 1644511149
transform 1 0 12420 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_70_135
timestamp 1644511149
transform 1 0 13524 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_70_151
timestamp 1644511149
transform 1 0 14996 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_70_161
timestamp 1644511149
transform 1 0 15916 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_169
timestamp 1644511149
transform 1 0 16652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_70_176
timestamp 1644511149
transform 1 0 17296 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_70_192
timestamp 1644511149
transform 1 0 18768 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_70_203
timestamp 1644511149
transform 1 0 19780 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_211
timestamp 1644511149
transform 1 0 20516 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_70_232
timestamp 1644511149
transform 1 0 22448 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_70_244
timestamp 1644511149
transform 1 0 23552 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_70_259
timestamp 1644511149
transform 1 0 24932 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_267
timestamp 1644511149
transform 1 0 25668 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_70_276
timestamp 1644511149
transform 1 0 26496 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_284
timestamp 1644511149
transform 1 0 27232 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_70_295
timestamp 1644511149
transform 1 0 28244 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_70_302
timestamp 1644511149
transform 1 0 28888 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_306
timestamp 1644511149
transform 1 0 29256 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_70_329
timestamp 1644511149
transform 1 0 31372 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_71_19
timestamp 1644511149
transform 1 0 2852 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_23
timestamp 1644511149
transform 1 0 3220 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_71_32
timestamp 1644511149
transform 1 0 4048 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_71_52
timestamp 1644511149
transform 1 0 5888 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_71_66
timestamp 1644511149
transform 1 0 7176 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_71_78
timestamp 1644511149
transform 1 0 8280 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_82
timestamp 1644511149
transform 1 0 8648 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_71_92
timestamp 1644511149
transform 1 0 9568 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_71_102
timestamp 1644511149
transform 1 0 10488 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_110
timestamp 1644511149
transform 1 0 11224 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_71_121
timestamp 1644511149
transform 1 0 12236 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_71_131
timestamp 1644511149
transform 1 0 13156 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_71_138
timestamp 1644511149
transform 1 0 13800 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_71_150
timestamp 1644511149
transform 1 0 14904 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_71_160
timestamp 1644511149
transform 1 0 15824 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_71_177
timestamp 1644511149
transform 1 0 17388 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_71_184
timestamp 1644511149
transform 1 0 18032 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_71_198
timestamp 1644511149
transform 1 0 19320 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_71_205
timestamp 1644511149
transform 1 0 19964 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_71_219
timestamp 1644511149
transform 1 0 21252 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_71_231
timestamp 1644511149
transform 1 0 22356 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_235
timestamp 1644511149
transform 1 0 22724 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_71_244
timestamp 1644511149
transform 1 0 23552 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_248
timestamp 1644511149
transform 1 0 23920 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_71_260
timestamp 1644511149
transform 1 0 25024 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_71_272
timestamp 1644511149
transform 1 0 26128 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_71_289
timestamp 1644511149
transform 1 0 27692 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_71_301
timestamp 1644511149
transform 1 0 28796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_71_313
timestamp 1644511149
transform 1 0 29900 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_71_325
timestamp 1644511149
transform 1 0 31004 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_5
timestamp 1644511149
transform 1 0 1564 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_72_12
timestamp 1644511149
transform 1 0 2208 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_72_24
timestamp 1644511149
transform 1 0 3312 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_37
timestamp 1644511149
transform 1 0 4508 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_49
timestamp 1644511149
transform 1 0 5612 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_72_70
timestamp 1644511149
transform 1 0 7544 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_72_80
timestamp 1644511149
transform 1 0 8464 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_89
timestamp 1644511149
transform 1 0 9292 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_72_106
timestamp 1644511149
transform 1 0 10856 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_72_118
timestamp 1644511149
transform 1 0 11960 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_126
timestamp 1644511149
transform 1 0 12696 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_72_135
timestamp 1644511149
transform 1 0 13524 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_145
timestamp 1644511149
transform 1 0 14444 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_72_162
timestamp 1644511149
transform 1 0 16008 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_72_174
timestamp 1644511149
transform 1 0 17112 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_72_186
timestamp 1644511149
transform 1 0 18216 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_194
timestamp 1644511149
transform 1 0 18952 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_72_213
timestamp 1644511149
transform 1 0 20700 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_221
timestamp 1644511149
transform 1 0 21436 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_72_225
timestamp 1644511149
transform 1 0 21804 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_72_237
timestamp 1644511149
transform 1 0 22908 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_72_247
timestamp 1644511149
transform 1 0 23828 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_72_269
timestamp 1644511149
transform 1 0 25852 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_72_281
timestamp 1644511149
transform 1 0 26956 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_72_293
timestamp 1644511149
transform 1 0 28060 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_72_303
timestamp 1644511149
transform 1 0 28980 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1644511149
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_72_325
timestamp 1644511149
transform 1 0 31004 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILLER_73_19
timestamp 1644511149
transform 1 0 2852 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_27
timestamp 1644511149
transform 1 0 3588 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_73_45
timestamp 1644511149
transform 1 0 5244 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_53
timestamp 1644511149
transform 1 0 5980 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_73_73
timestamp 1644511149
transform 1 0 7820 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_77
timestamp 1644511149
transform 1 0 8188 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_73_95
timestamp 1644511149
transform 1 0 9844 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_99
timestamp 1644511149
transform 1 0 10212 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_73_106
timestamp 1644511149
transform 1 0 10856 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_110
timestamp 1644511149
transform 1 0 11224 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_73_130
timestamp 1644511149
transform 1 0 13064 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_73_142
timestamp 1644511149
transform 1 0 14168 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_73_154
timestamp 1644511149
transform 1 0 15272 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_73_164
timestamp 1644511149
transform 1 0 16192 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_73_185
timestamp 1644511149
transform 1 0 18124 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_73_205
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_209
timestamp 1644511149
transform 1 0 20332 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_73_213
timestamp 1644511149
transform 1 0 20700 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_73_220
timestamp 1644511149
transform 1 0 21344 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_73_241
timestamp 1644511149
transform 1 0 23276 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_73_251
timestamp 1644511149
transform 1 0 24196 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_259
timestamp 1644511149
transform 1 0 24932 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_73_276
timestamp 1644511149
transform 1 0 26496 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_73_297
timestamp 1644511149
transform 1 0 28428 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_73_317
timestamp 1644511149
transform 1 0 30268 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_73_324
timestamp 1644511149
transform 1 0 30912 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_332
timestamp 1644511149
transform 1 0 31648 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_7
timestamp 1644511149
transform 1 0 1748 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_74_24
timestamp 1644511149
transform 1 0 3312 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_74_35
timestamp 1644511149
transform 1 0 4324 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_74_47
timestamp 1644511149
transform 1 0 5428 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_74_57
timestamp 1644511149
transform 1 0 6348 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_61
timestamp 1644511149
transform 1 0 6716 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_63
timestamp 1644511149
transform 1 0 6900 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_74_80
timestamp 1644511149
transform 1 0 8464 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_74_91
timestamp 1644511149
transform 1 0 9476 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_95
timestamp 1644511149
transform 1 0 9844 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_74_113
timestamp 1644511149
transform 1 0 11500 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_117
timestamp 1644511149
transform 1 0 11868 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_74_135
timestamp 1644511149
transform 1 0 13524 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_74_157
timestamp 1644511149
transform 1 0 15548 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_181
timestamp 1644511149
transform 1 0 17756 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_183
timestamp 1644511149
transform 1 0 17940 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_74_192
timestamp 1644511149
transform 1 0 18768 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_74_203
timestamp 1644511149
transform 1 0 19780 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_211
timestamp 1644511149
transform 1 0 20516 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_74_228
timestamp 1644511149
transform 1 0 22080 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_74_248
timestamp 1644511149
transform 1 0 23920 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_74_269
timestamp 1644511149
transform 1 0 25852 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_74_279
timestamp 1644511149
transform 1 0 26772 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_287
timestamp 1644511149
transform 1 0 27508 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_74_304
timestamp 1644511149
transform 1 0 29072 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_74_315
timestamp 1644511149
transform 1 0 30084 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_74_322
timestamp 1644511149
transform 1 0 30728 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_74_329
timestamp 1644511149
transform 1 0 31372 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_75_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_75_13
timestamp 1644511149
transform 1 0 2300 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_75_23
timestamp 1644511149
transform 1 0 3220 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_27
timestamp 1644511149
transform 1 0 3588 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_75_29
timestamp 1644511149
transform 1 0 3772 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1644511149
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_75_51
timestamp 1644511149
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_75_72
timestamp 1644511149
transform 1 0 7728 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_75_80
timestamp 1644511149
transform 1 0 8464 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_75_91
timestamp 1644511149
transform 1 0 9476 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_98
timestamp 1644511149
transform 1 0 10120 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_110
timestamp 1644511149
transform 1 0 11224 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_8  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_121
timestamp 1644511149
transform 1 0 12236 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_123
timestamp 1644511149
transform 1 0 12420 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILLER_75_130
timestamp 1644511149
transform 1 0 13064 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_138
timestamp 1644511149
transform 1 0 13800 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_141
timestamp 1644511149
transform 1 0 14076 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_4  FILLER_75_156
timestamp 1644511149
transform 1 0 15456 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_75_164
timestamp 1644511149
transform 1 0 16192 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_75_175
timestamp 1644511149
transform 1 0 17204 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILLER_75_189
timestamp 1644511149
transform 1 0 18492 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_195
timestamp 1644511149
transform 1 0 19044 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_75_197
timestamp 1644511149
transform 1 0 19228 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_201
timestamp 1644511149
transform 1 0 19596 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_75_219
timestamp 1644511149
transform 1 0 21252 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_229
timestamp 1644511149
transform 1 0 22172 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_75_233
timestamp 1644511149
transform 1 0 22540 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_75_240
timestamp 1644511149
transform 1 0 23184 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_75_248
timestamp 1644511149
transform 1 0 23920 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_75_256
timestamp 1644511149
transform 1 0 24656 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_264
timestamp 1644511149
transform 1 0 25392 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_75_269
timestamp 1644511149
transform 1 0 25852 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_75_276
timestamp 1644511149
transform 1 0 26496 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILLER_75_287
timestamp 1644511149
transform 1 0 27508 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_295
timestamp 1644511149
transform 1 0 28244 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILLER_75_303
timestamp 1644511149
transform 1 0 28980 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_307
timestamp 1644511149
transform 1 0 29348 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_75_312
timestamp 1644511149
transform 1 0 29808 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_4  FILLER_75_319
timestamp 1644511149
transform 1 0 30452 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_323
timestamp 1644511149
transform 1 0 30820 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_325
timestamp 1644511149
transform 1 0 31004 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_4  FILLER_75_329
timestamp 1644511149
transform 1 0 31372 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 32016 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 32016 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 32016 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 32016 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 32016 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 32016 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 32016 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 32016 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 32016 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 32016 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 32016 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 32016 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 32016 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 32016 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 32016 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 32016 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 32016 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 32016 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 32016 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 32016 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 32016 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 32016 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 32016 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 32016 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 32016 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 32016 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 32016 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 32016 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 32016 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 32016 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 32016 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 32016 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 32016 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 32016 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 32016 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 32016 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 32016 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 32016 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 32016 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 32016 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 32016 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 32016 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 32016 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 32016 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 32016 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 32016 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 32016 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 32016 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 32016 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 32016 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 32016 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 32016 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 32016 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 32016 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 32016 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 32016 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 32016 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 32016 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 32016 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 32016 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 32016 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 32016 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 32016 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 32016 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 32016 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 32016 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 32016 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 32016 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 32016 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 32016 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 32016 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 32016 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 32016 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 32016 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 32016 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 32016 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 26864 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 29440 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 26864 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 3680 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 8832 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 13984 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 19136 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 24288 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 29440 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__and3b_1  _1311_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1312_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7544 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1313_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8740 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1314_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7544 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1315_
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1316_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7544 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_2  _1317_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6440 0 1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__and2_1  _1318_
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1319_
timestamp 1644511149
transform 1 0 3772 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1320_
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1321_
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1322_
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1323_
timestamp 1644511149
transform 1 0 1656 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_2  _1324_
timestamp 1644511149
transform 1 0 1656 0 1 16320
box -38 -48 1694 592
use sky130_fd_sc_hd__buf_2  _1325_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1326_
timestamp 1644511149
transform 1 0 16192 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1327_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17388 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1328_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1329_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12420 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1330_
timestamp 1644511149
transform 1 0 12880 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1331_
timestamp 1644511149
transform 1 0 13248 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _1332_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22632 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1333_
timestamp 1644511149
transform 1 0 9108 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1334_
timestamp 1644511149
transform 1 0 7636 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1335_
timestamp 1644511149
transform 1 0 7636 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1336_
timestamp 1644511149
transform 1 0 6532 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1337_
timestamp 1644511149
transform 1 0 7728 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_2  _1338_
timestamp 1644511149
transform 1 0 6808 0 1 14144
box -38 -48 1694 592
use sky130_fd_sc_hd__and2_1  _1339_
timestamp 1644511149
transform 1 0 15824 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1340_
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1341_
timestamp 1644511149
transform 1 0 1932 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1342_
timestamp 1644511149
transform 1 0 2024 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__and3b_1  _1343_
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1344_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1840 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1345_
timestamp 1644511149
transform 1 0 2576 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1346_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2944 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1347_
timestamp 1644511149
transform 1 0 5428 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1348_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3312 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _1349_
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1350_
timestamp 1644511149
transform 1 0 18860 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1351_
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1352_
timestamp 1644511149
transform 1 0 15272 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1353_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1354_
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1355_
timestamp 1644511149
transform 1 0 6716 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1356_
timestamp 1644511149
transform 1 0 9384 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1357_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1358_
timestamp 1644511149
transform 1 0 7912 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1359_
timestamp 1644511149
transform 1 0 7728 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1360_
timestamp 1644511149
transform 1 0 8188 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _1361_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _1362_
timestamp 1644511149
transform 1 0 15364 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1363_
timestamp 1644511149
transform 1 0 4600 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1364_
timestamp 1644511149
transform 1 0 1748 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1365_
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1366_
timestamp 1644511149
transform 1 0 2116 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1367_
timestamp 1644511149
transform 1 0 2576 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_2  _1368_
timestamp 1644511149
transform 1 0 2576 0 -1 14144
box -38 -48 1694 592
use sky130_fd_sc_hd__buf_2  _1369_
timestamp 1644511149
transform 1 0 19320 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1370_
timestamp 1644511149
transform 1 0 15364 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1371_
timestamp 1644511149
transform 1 0 15088 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1372_
timestamp 1644511149
transform 1 0 11960 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _1373_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14352 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1374_
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1375_
timestamp 1644511149
transform 1 0 6348 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1376_
timestamp 1644511149
transform 1 0 5612 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1377_
timestamp 1644511149
transform 1 0 4784 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1378_
timestamp 1644511149
transform 1 0 3956 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_2  _1379_
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__and2_1  _1380_
timestamp 1644511149
transform 1 0 16192 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1381_
timestamp 1644511149
transform 1 0 4968 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1382_
timestamp 1644511149
transform 1 0 7912 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1383_
timestamp 1644511149
transform 1 0 5060 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1384_
timestamp 1644511149
transform 1 0 4968 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1385_
timestamp 1644511149
transform 1 0 4968 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_2  _1386_
timestamp 1644511149
transform 1 0 4600 0 1 16320
box -38 -48 1694 592
use sky130_fd_sc_hd__mux2_1  _1387_
timestamp 1644511149
transform 1 0 16652 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1388_
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1389_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1390_
timestamp 1644511149
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1391_
timestamp 1644511149
transform 1 0 15732 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1392_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15364 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1393_
timestamp 1644511149
transform 1 0 15088 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1394_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14628 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1395_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1396_
timestamp 1644511149
transform 1 0 15640 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1397_
timestamp 1644511149
transform 1 0 16744 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1398_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16928 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1399_
timestamp 1644511149
transform 1 0 15548 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1400_
timestamp 1644511149
transform 1 0 16652 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1401_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16560 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1402_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16744 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1403_
timestamp 1644511149
transform 1 0 17664 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_2  _1404_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21252 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1405_
timestamp 1644511149
transform 1 0 22816 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1406_
timestamp 1644511149
transform 1 0 24104 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1407_
timestamp 1644511149
transform 1 0 24196 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1408_
timestamp 1644511149
transform 1 0 25576 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1409_
timestamp 1644511149
transform 1 0 24104 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1410_
timestamp 1644511149
transform 1 0 25668 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1411_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22172 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_4  _1412_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1413_
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1414_
timestamp 1644511149
transform 1 0 12788 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1415_
timestamp 1644511149
transform 1 0 17848 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1416_
timestamp 1644511149
transform 1 0 23552 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1417_
timestamp 1644511149
transform 1 0 23276 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _1418_
timestamp 1644511149
transform 1 0 23184 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_4  _1419_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23368 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_4  _1420_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1421_
timestamp 1644511149
transform 1 0 29256 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_2  _1422_
timestamp 1644511149
transform 1 0 30544 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_4  _1423_
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1424_
timestamp 1644511149
transform 1 0 23644 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1425_
timestamp 1644511149
transform 1 0 19964 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1426_
timestamp 1644511149
transform 1 0 19320 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1427_
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _1428_
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _1429_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23276 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1430_
timestamp 1644511149
transform 1 0 15732 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1431_
timestamp 1644511149
transform 1 0 16652 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1432_
timestamp 1644511149
transform 1 0 4140 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1433_
timestamp 1644511149
transform 1 0 1932 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1434_
timestamp 1644511149
transform 1 0 3036 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1435_
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1436_
timestamp 1644511149
transform 1 0 2760 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_2  _1437_
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__or2_1  _1438_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20516 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1439_
timestamp 1644511149
transform 1 0 21068 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1440_
timestamp 1644511149
transform 1 0 22172 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1441_
timestamp 1644511149
transform 1 0 23276 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1442_
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1443_
timestamp 1644511149
transform 1 0 6716 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1444_
timestamp 1644511149
transform 1 0 7544 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1445_
timestamp 1644511149
transform 1 0 6716 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1446_
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1447_
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1448_
timestamp 1644511149
transform 1 0 6256 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1449_
timestamp 1644511149
transform 1 0 6900 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1450_
timestamp 1644511149
transform 1 0 6900 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _1451_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7728 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1452_
timestamp 1644511149
transform 1 0 22632 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1453_
timestamp 1644511149
transform 1 0 22080 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1454_
timestamp 1644511149
transform 1 0 22816 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1455_
timestamp 1644511149
transform 1 0 24012 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1456_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23460 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1457_
timestamp 1644511149
transform 1 0 23552 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1458_
timestamp 1644511149
transform 1 0 26680 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1459_
timestamp 1644511149
transform 1 0 23092 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1460_
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1461_
timestamp 1644511149
transform 1 0 15732 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1462_
timestamp 1644511149
transform 1 0 17204 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _1463_
timestamp 1644511149
transform 1 0 17296 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1464_
timestamp 1644511149
transform 1 0 24012 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1465_
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1466_
timestamp 1644511149
transform 1 0 18308 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1467_
timestamp 1644511149
transform 1 0 18492 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_2  _1468_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17112 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1469_
timestamp 1644511149
transform 1 0 28612 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1470_
timestamp 1644511149
transform 1 0 25760 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _1471_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1472_
timestamp 1644511149
transform 1 0 25852 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1473_
timestamp 1644511149
transform 1 0 26588 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1474_
timestamp 1644511149
transform 1 0 27232 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1475_
timestamp 1644511149
transform 1 0 27600 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1476_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28612 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1477_
timestamp 1644511149
transform 1 0 27324 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1478_
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1479_
timestamp 1644511149
transform 1 0 25300 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1480_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25484 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1481_
timestamp 1644511149
transform 1 0 25484 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_2  _1482_
timestamp 1644511149
transform 1 0 23276 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1483_
timestamp 1644511149
transform 1 0 23276 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1484_
timestamp 1644511149
transform 1 0 23276 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1485_
timestamp 1644511149
transform 1 0 23644 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1486_
timestamp 1644511149
transform 1 0 11040 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1487_
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1488_
timestamp 1644511149
transform 1 0 20148 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1489_
timestamp 1644511149
transform 1 0 9568 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1490_
timestamp 1644511149
transform 1 0 11500 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1491_
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1492_
timestamp 1644511149
transform 1 0 6900 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1493_
timestamp 1644511149
transform 1 0 7452 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_2  _1494_
timestamp 1644511149
transform 1 0 7544 0 -1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__and2_1  _1495_
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1496_
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1497_
timestamp 1644511149
transform 1 0 15364 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1498_
timestamp 1644511149
transform 1 0 6900 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1499_
timestamp 1644511149
transform 1 0 8004 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1500_
timestamp 1644511149
transform 1 0 6716 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1501_
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1502_
timestamp 1644511149
transform 1 0 6256 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_2  _1503_
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__a21oi_1  _1504_
timestamp 1644511149
transform 1 0 13248 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1505_
timestamp 1644511149
transform 1 0 7360 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1506_
timestamp 1644511149
transform 1 0 4968 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1507_
timestamp 1644511149
transform 1 0 6532 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1508_
timestamp 1644511149
transform 1 0 6624 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1509_
timestamp 1644511149
transform 1 0 8740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1510_
timestamp 1644511149
transform 1 0 7728 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1511_
timestamp 1644511149
transform 1 0 5060 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1512_
timestamp 1644511149
transform 1 0 6256 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1513_
timestamp 1644511149
transform 1 0 6256 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _1514_
timestamp 1644511149
transform 1 0 11684 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1515_
timestamp 1644511149
transform 1 0 11868 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1516_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_2  _1517_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1518_
timestamp 1644511149
transform 1 0 14536 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1519_
timestamp 1644511149
transform 1 0 14628 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1520_
timestamp 1644511149
transform 1 0 13984 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1521_
timestamp 1644511149
transform 1 0 14536 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1522_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14536 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1523_
timestamp 1644511149
transform 1 0 14076 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1524_
timestamp 1644511149
transform 1 0 15088 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1525_
timestamp 1644511149
transform 1 0 14076 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1526_
timestamp 1644511149
transform 1 0 14536 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1527_
timestamp 1644511149
transform 1 0 15548 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1528_
timestamp 1644511149
transform 1 0 2392 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1529_
timestamp 1644511149
transform 1 0 2392 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1530_
timestamp 1644511149
transform 1 0 3220 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1531_
timestamp 1644511149
transform 1 0 2576 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1532_
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1533_
timestamp 1644511149
transform 1 0 1656 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1534_
timestamp 1644511149
transform 1 0 2300 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  _1535_
timestamp 1644511149
transform 1 0 2576 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1536_
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1537_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15364 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1538_
timestamp 1644511149
transform 1 0 18492 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1539_
timestamp 1644511149
transform 1 0 15364 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_2  _1540_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15364 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1541_
timestamp 1644511149
transform 1 0 17204 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  _1542_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17204 0 -1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1543_
timestamp 1644511149
transform 1 0 16560 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1544_
timestamp 1644511149
transform 1 0 16468 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1545_
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1546_
timestamp 1644511149
transform 1 0 15548 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1547_
timestamp 1644511149
transform 1 0 12696 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1548_
timestamp 1644511149
transform 1 0 9936 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1549_
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1550_
timestamp 1644511149
transform 1 0 6624 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__and3b_1  _1551_
timestamp 1644511149
transform 1 0 6072 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1552_
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1553_
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1554_
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1555_
timestamp 1644511149
transform 1 0 5704 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1556_
timestamp 1644511149
transform 1 0 6440 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1557_
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1558_
timestamp 1644511149
transform 1 0 13340 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1559_
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_2  _1560_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12880 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1561_
timestamp 1644511149
transform 1 0 9108 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1562_
timestamp 1644511149
transform 1 0 9752 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1563_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10304 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1564_
timestamp 1644511149
transform 1 0 9752 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_2  _1565_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9384 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1566_
timestamp 1644511149
transform 1 0 6900 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1567_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7912 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1568_
timestamp 1644511149
transform 1 0 7820 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1569_
timestamp 1644511149
transform 1 0 7636 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _1570_
timestamp 1644511149
transform 1 0 6808 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1571_
timestamp 1644511149
transform 1 0 12420 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1572_
timestamp 1644511149
transform 1 0 12972 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1573_
timestamp 1644511149
transform 1 0 10672 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1574_
timestamp 1644511149
transform 1 0 12052 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o221ai_4  _1575_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11316 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _1576_
timestamp 1644511149
transform 1 0 6624 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1577_
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1578_
timestamp 1644511149
transform 1 0 6256 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a32oi_4  _1579_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9292 0 1 19584
box -38 -48 2062 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1580_
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__nor3_2  _1581_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8188 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1582_
timestamp 1644511149
transform 1 0 6716 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1583_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6716 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1584_
timestamp 1644511149
transform 1 0 6164 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1585_
timestamp 1644511149
transform 1 0 6440 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_2  _1586_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11592 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1587_
timestamp 1644511149
transform 1 0 7728 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1588_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7544 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1589_
timestamp 1644511149
transform 1 0 6348 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _1590_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6624 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1591_
timestamp 1644511149
transform 1 0 7728 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _1592_
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1593_
timestamp 1644511149
transform 1 0 8188 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1594_
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1595_
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1596_
timestamp 1644511149
transform 1 0 7820 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1597_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9292 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1598_
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1599_
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1600_
timestamp 1644511149
transform 1 0 10304 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_2  _1601_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__and3b_1  _1602_
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1603_
timestamp 1644511149
transform 1 0 12512 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _1604_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12144 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _1605_
timestamp 1644511149
transform 1 0 12696 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1606_
timestamp 1644511149
transform 1 0 12972 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1607_
timestamp 1644511149
transform 1 0 15364 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_2  _1608_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _1609_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20792 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_4  _1610_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20792 0 1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_1  _1611_
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1612_
timestamp 1644511149
transform 1 0 24104 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1613_
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1614_
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _1615_
timestamp 1644511149
transform 1 0 10396 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1616_
timestamp 1644511149
transform 1 0 9016 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1617_
timestamp 1644511149
transform 1 0 11316 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1618_
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1619_
timestamp 1644511149
transform 1 0 9660 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a31oi_4  _1620_
timestamp 1644511149
transform 1 0 8924 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1621_
timestamp 1644511149
transform 1 0 8740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1622_
timestamp 1644511149
transform 1 0 7636 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1623_
timestamp 1644511149
transform 1 0 9384 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and3b_1  _1624_
timestamp 1644511149
transform 1 0 7820 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1625_
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1626_
timestamp 1644511149
transform 1 0 7544 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1627_
timestamp 1644511149
transform 1 0 9108 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1628_
timestamp 1644511149
transform 1 0 7912 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_4  _1629_
timestamp 1644511149
transform 1 0 8648 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1630_
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1631_
timestamp 1644511149
transform 1 0 13156 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1632_
timestamp 1644511149
transform 1 0 11776 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1633_
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1634_
timestamp 1644511149
transform 1 0 20148 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1635_
timestamp 1644511149
transform 1 0 5612 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1636_
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1637_
timestamp 1644511149
transform 1 0 12972 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1638_
timestamp 1644511149
transform 1 0 9384 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1639_
timestamp 1644511149
transform 1 0 9016 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1640_
timestamp 1644511149
transform 1 0 11408 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1641_
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1642_
timestamp 1644511149
transform 1 0 6716 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1643_
timestamp 1644511149
transform 1 0 9292 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1644_
timestamp 1644511149
transform 1 0 10212 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1645_
timestamp 1644511149
transform 1 0 7728 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1646_
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1647_
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _1648_
timestamp 1644511149
transform 1 0 5520 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1649_
timestamp 1644511149
transform 1 0 5612 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1650_
timestamp 1644511149
transform 1 0 4048 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1651_
timestamp 1644511149
transform 1 0 5336 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _1652_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10304 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1653_
timestamp 1644511149
transform 1 0 6532 0 -1 40256
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1654_
timestamp 1644511149
transform 1 0 5060 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1655_
timestamp 1644511149
transform 1 0 4692 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1656_
timestamp 1644511149
transform 1 0 4324 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1657_
timestamp 1644511149
transform 1 0 5428 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1658_
timestamp 1644511149
transform 1 0 8004 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1659_
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1660_
timestamp 1644511149
transform 1 0 11684 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _1661_
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1662_
timestamp 1644511149
transform 1 0 21344 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1663_
timestamp 1644511149
transform 1 0 22724 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1664_
timestamp 1644511149
transform 1 0 16928 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1665_
timestamp 1644511149
transform 1 0 22724 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1666_
timestamp 1644511149
transform 1 0 22632 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1667_
timestamp 1644511149
transform 1 0 22724 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1668_
timestamp 1644511149
transform 1 0 18308 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1669_
timestamp 1644511149
transform 1 0 20148 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1670_
timestamp 1644511149
transform 1 0 19228 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1671_
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1672_
timestamp 1644511149
transform 1 0 25944 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1673_
timestamp 1644511149
transform 1 0 23000 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1674_
timestamp 1644511149
transform 1 0 18584 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1675_
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1676_
timestamp 1644511149
transform 1 0 18584 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1677_
timestamp 1644511149
transform 1 0 25576 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1678_
timestamp 1644511149
transform 1 0 25208 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  _1679_
timestamp 1644511149
transform 1 0 29440 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _1680_
timestamp 1644511149
transform 1 0 29164 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  _1681_
timestamp 1644511149
transform 1 0 23644 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1682_
timestamp 1644511149
transform 1 0 20516 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1683_
timestamp 1644511149
transform 1 0 20608 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _1684_
timestamp 1644511149
transform 1 0 21068 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1685_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1686_
timestamp 1644511149
transform 1 0 27876 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _1687_
timestamp 1644511149
transform 1 0 27140 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__a31oi_1  _1688_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22724 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1689_
timestamp 1644511149
transform 1 0 24748 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1690_
timestamp 1644511149
transform 1 0 25392 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1691_
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1692_
timestamp 1644511149
transform 1 0 26496 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1693_
timestamp 1644511149
transform 1 0 25852 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1694_
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a2111o_1  _1695_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24196 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__o2111a_1  _1696_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24104 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1697_
timestamp 1644511149
transform 1 0 26036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1698_
timestamp 1644511149
transform 1 0 20792 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1699_
timestamp 1644511149
transform 1 0 22632 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1700_
timestamp 1644511149
transform 1 0 20792 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1701_
timestamp 1644511149
transform 1 0 25116 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1702_
timestamp 1644511149
transform 1 0 22816 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1703_
timestamp 1644511149
transform 1 0 23092 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1704_
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1705_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26036 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1706_
timestamp 1644511149
transform 1 0 27232 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1707_
timestamp 1644511149
transform 1 0 28612 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _1708_
timestamp 1644511149
transform 1 0 24564 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1709_
timestamp 1644511149
transform 1 0 27692 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1710_
timestamp 1644511149
transform 1 0 18492 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1711_
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1712_
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_2  _1713_
timestamp 1644511149
transform 1 0 16836 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1714_
timestamp 1644511149
transform 1 0 31096 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1715_
timestamp 1644511149
transform 1 0 27508 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1716_
timestamp 1644511149
transform 1 0 24840 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1717_
timestamp 1644511149
transform 1 0 28980 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1718_
timestamp 1644511149
transform 1 0 28796 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1719_
timestamp 1644511149
transform 1 0 28336 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1720_
timestamp 1644511149
transform 1 0 28060 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1721_
timestamp 1644511149
transform 1 0 24380 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1722_
timestamp 1644511149
transform 1 0 29808 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1723_
timestamp 1644511149
transform 1 0 29624 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1724_
timestamp 1644511149
transform 1 0 28060 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1725_
timestamp 1644511149
transform 1 0 29532 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1726_
timestamp 1644511149
transform 1 0 30544 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1727_
timestamp 1644511149
transform 1 0 28152 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1728_
timestamp 1644511149
transform 1 0 18216 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1729_
timestamp 1644511149
transform 1 0 21068 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1730_
timestamp 1644511149
transform 1 0 18492 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1731_
timestamp 1644511149
transform 1 0 19412 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1732_
timestamp 1644511149
transform 1 0 27600 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1733_
timestamp 1644511149
transform 1 0 28612 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1734_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1735_
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1736_
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1737_
timestamp 1644511149
transform 1 0 17756 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1738_
timestamp 1644511149
transform 1 0 17940 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1739_
timestamp 1644511149
transform 1 0 24748 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1740_
timestamp 1644511149
transform 1 0 19504 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1741_
timestamp 1644511149
transform 1 0 19688 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1742_
timestamp 1644511149
transform 1 0 20700 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1743_
timestamp 1644511149
transform 1 0 25208 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _1744_
timestamp 1644511149
transform 1 0 27140 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__and2b_1  _1745_
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1746_
timestamp 1644511149
transform 1 0 25576 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1747_
timestamp 1644511149
transform 1 0 24932 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1748_
timestamp 1644511149
transform 1 0 26220 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1749_
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1750_
timestamp 1644511149
transform 1 0 27048 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1751_
timestamp 1644511149
transform 1 0 21528 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1752_
timestamp 1644511149
transform 1 0 20792 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1753_
timestamp 1644511149
transform 1 0 19780 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1754_
timestamp 1644511149
transform 1 0 20700 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1755_
timestamp 1644511149
transform 1 0 20608 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1756_
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1757_
timestamp 1644511149
transform 1 0 25944 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1758_
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1759_
timestamp 1644511149
transform 1 0 25576 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1760_
timestamp 1644511149
transform 1 0 25760 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1761_
timestamp 1644511149
transform 1 0 25668 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1762_
timestamp 1644511149
transform 1 0 26128 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1763_
timestamp 1644511149
transform 1 0 25208 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1764_
timestamp 1644511149
transform 1 0 21988 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1765_
timestamp 1644511149
transform 1 0 21896 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1766_
timestamp 1644511149
transform 1 0 22540 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1767_
timestamp 1644511149
transform 1 0 25024 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1768_
timestamp 1644511149
transform 1 0 23920 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1769_
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1770_
timestamp 1644511149
transform 1 0 24380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _1771_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23092 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_2  _1772_
timestamp 1644511149
transform 1 0 23368 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1773_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27048 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1774_
timestamp 1644511149
transform 1 0 27140 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1775_
timestamp 1644511149
transform 1 0 27508 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1776_
timestamp 1644511149
transform 1 0 27508 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1777_
timestamp 1644511149
transform 1 0 27416 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1778_
timestamp 1644511149
transform 1 0 28520 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1779_
timestamp 1644511149
transform 1 0 31096 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _1780_
timestamp 1644511149
transform 1 0 28520 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1781_
timestamp 1644511149
transform 1 0 27048 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1782_
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1783_
timestamp 1644511149
transform 1 0 28796 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _1784_
timestamp 1644511149
transform 1 0 23184 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1785_
timestamp 1644511149
transform 1 0 23184 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1786_
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1787_
timestamp 1644511149
transform 1 0 27692 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1788_
timestamp 1644511149
transform 1 0 25852 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1789_
timestamp 1644511149
transform 1 0 25024 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1790_
timestamp 1644511149
transform 1 0 24748 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1791_
timestamp 1644511149
transform 1 0 25024 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1792_
timestamp 1644511149
transform 1 0 31096 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _1793_
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1794_
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1795_
timestamp 1644511149
transform 1 0 24288 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1796_
timestamp 1644511149
transform 1 0 15640 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1797_
timestamp 1644511149
transform 1 0 7360 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1798_
timestamp 1644511149
transform 1 0 14720 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1799_
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1800_
timestamp 1644511149
transform 1 0 15824 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1801_
timestamp 1644511149
transform 1 0 16192 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1802_
timestamp 1644511149
transform 1 0 9936 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1803_
timestamp 1644511149
transform 1 0 17848 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1804_
timestamp 1644511149
transform 1 0 15824 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1805_
timestamp 1644511149
transform 1 0 9844 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1806_
timestamp 1644511149
transform 1 0 12972 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1807_
timestamp 1644511149
transform 1 0 12420 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1808_
timestamp 1644511149
transform 1 0 9292 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1809_
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1810_
timestamp 1644511149
transform 1 0 10396 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1811_
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1812_
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1813_
timestamp 1644511149
transform 1 0 7728 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1814_
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1815_
timestamp 1644511149
transform 1 0 8188 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1816_
timestamp 1644511149
transform 1 0 6808 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1817_
timestamp 1644511149
transform 1 0 7728 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1818_
timestamp 1644511149
transform 1 0 7176 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1819_
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1820_
timestamp 1644511149
transform 1 0 5060 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1821_
timestamp 1644511149
transform 1 0 13156 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1822_
timestamp 1644511149
transform 1 0 8096 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1823_
timestamp 1644511149
transform 1 0 3680 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1824_
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1825_
timestamp 1644511149
transform 1 0 4140 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1826_
timestamp 1644511149
transform 1 0 4232 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1827_
timestamp 1644511149
transform 1 0 4324 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1828_
timestamp 1644511149
transform 1 0 3128 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1829_
timestamp 1644511149
transform 1 0 2208 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1830_
timestamp 1644511149
transform 1 0 2944 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1831_
timestamp 1644511149
transform 1 0 2576 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1832_
timestamp 1644511149
transform 1 0 1840 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1833_
timestamp 1644511149
transform 1 0 2392 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1834_
timestamp 1644511149
transform 1 0 4968 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1835_
timestamp 1644511149
transform 1 0 17848 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1836_
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1837_
timestamp 1644511149
transform 1 0 4416 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1838_
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1839_
timestamp 1644511149
transform 1 0 3220 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1840_
timestamp 1644511149
transform 1 0 2392 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1841_
timestamp 1644511149
transform 1 0 2576 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1842_
timestamp 1644511149
transform 1 0 1656 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1843_
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1844_
timestamp 1644511149
transform 1 0 2760 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1845_
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1846_
timestamp 1644511149
transform 1 0 5704 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1847_
timestamp 1644511149
transform 1 0 5060 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1848_
timestamp 1644511149
transform 1 0 2852 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1849_
timestamp 1644511149
transform 1 0 7544 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1850_
timestamp 1644511149
transform 1 0 9476 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1851_
timestamp 1644511149
transform 1 0 5612 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1852_
timestamp 1644511149
transform 1 0 6440 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1853_
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1854_
timestamp 1644511149
transform 1 0 7544 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1855_
timestamp 1644511149
transform 1 0 7544 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1856_
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1857_
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1858_
timestamp 1644511149
transform 1 0 8740 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1859_
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1860_
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1861_
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1862_
timestamp 1644511149
transform 1 0 9108 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1863_
timestamp 1644511149
transform 1 0 16560 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1864_
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1865_
timestamp 1644511149
transform 1 0 9936 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1866_
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_1  _1867_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1868_
timestamp 1644511149
transform 1 0 16928 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1869_
timestamp 1644511149
transform 1 0 16468 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1870_
timestamp 1644511149
transform 1 0 11408 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1871_
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1872_
timestamp 1644511149
transform 1 0 6624 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1873_
timestamp 1644511149
transform 1 0 4048 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1874_
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1875_
timestamp 1644511149
transform 1 0 3588 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1876_
timestamp 1644511149
transform 1 0 1840 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1877_
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1878_
timestamp 1644511149
transform 1 0 2760 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1879_
timestamp 1644511149
transform 1 0 2300 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1880_
timestamp 1644511149
transform 1 0 1840 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1881_
timestamp 1644511149
transform 1 0 2300 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1882_
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1883_
timestamp 1644511149
transform 1 0 4324 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1884_
timestamp 1644511149
transform 1 0 2668 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1885_
timestamp 1644511149
transform 1 0 2208 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1886_
timestamp 1644511149
transform 1 0 4324 0 1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1887_
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1888_
timestamp 1644511149
transform 1 0 3128 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1889_
timestamp 1644511149
transform 1 0 2576 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1890_
timestamp 1644511149
transform 1 0 2576 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1891_
timestamp 1644511149
transform 1 0 1656 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1892_
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1893_
timestamp 1644511149
transform 1 0 2668 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1894_
timestamp 1644511149
transform 1 0 3312 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1895_
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1896_
timestamp 1644511149
transform 1 0 8096 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1897_
timestamp 1644511149
transform 1 0 4692 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1898_
timestamp 1644511149
transform 1 0 5796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1899_
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1900_
timestamp 1644511149
transform 1 0 8188 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1901_
timestamp 1644511149
transform 1 0 9844 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1902_
timestamp 1644511149
transform 1 0 7544 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1903_
timestamp 1644511149
transform 1 0 7912 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1904_
timestamp 1644511149
transform 1 0 6992 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1905_
timestamp 1644511149
transform 1 0 9200 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1906_
timestamp 1644511149
transform 1 0 8096 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1907_
timestamp 1644511149
transform 1 0 7544 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1908_
timestamp 1644511149
transform 1 0 7728 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1909_
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1910_
timestamp 1644511149
transform 1 0 15824 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1911_
timestamp 1644511149
transform 1 0 8832 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1912_
timestamp 1644511149
transform 1 0 8924 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1913_
timestamp 1644511149
transform 1 0 16836 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1914_
timestamp 1644511149
transform 1 0 20792 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1915_
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1916_
timestamp 1644511149
transform 1 0 13524 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1917_
timestamp 1644511149
transform 1 0 11224 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1918_
timestamp 1644511149
transform 1 0 9936 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1919_
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1920_
timestamp 1644511149
transform 1 0 10304 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1921_
timestamp 1644511149
transform 1 0 10304 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1922_
timestamp 1644511149
transform 1 0 10396 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1923_
timestamp 1644511149
transform 1 0 11684 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1924_
timestamp 1644511149
transform 1 0 10488 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1925_
timestamp 1644511149
transform 1 0 22448 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1926_
timestamp 1644511149
transform 1 0 22632 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1927_
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _1928_
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1929_
timestamp 1644511149
transform 1 0 13340 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1930_
timestamp 1644511149
transform 1 0 12788 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1931_
timestamp 1644511149
transform 1 0 11684 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1932_
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1933_
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1934_
timestamp 1644511149
transform 1 0 12788 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1935_
timestamp 1644511149
transform 1 0 11868 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1936_
timestamp 1644511149
transform 1 0 12788 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1937_
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1938_
timestamp 1644511149
transform 1 0 13432 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1939_
timestamp 1644511149
transform 1 0 12512 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1940_
timestamp 1644511149
transform 1 0 20148 0 -1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1941_
timestamp 1644511149
transform 1 0 15824 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1942_
timestamp 1644511149
transform 1 0 14536 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1943_
timestamp 1644511149
transform 1 0 15640 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1944_
timestamp 1644511149
transform 1 0 14168 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1945_
timestamp 1644511149
transform 1 0 15364 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1946_
timestamp 1644511149
transform 1 0 18400 0 -1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1947_
timestamp 1644511149
transform 1 0 19688 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1948_
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1949_
timestamp 1644511149
transform 1 0 15272 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1950_
timestamp 1644511149
transform 1 0 16376 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1951_
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1952_
timestamp 1644511149
transform 1 0 17480 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1953_
timestamp 1644511149
transform 1 0 16744 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1954_
timestamp 1644511149
transform 1 0 21528 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1955_
timestamp 1644511149
transform 1 0 18032 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1956_
timestamp 1644511149
transform 1 0 17940 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1957_
timestamp 1644511149
transform 1 0 18032 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1958_
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1959_
timestamp 1644511149
transform 1 0 19320 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1960_
timestamp 1644511149
transform 1 0 17572 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1961_
timestamp 1644511149
transform 1 0 18584 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1962_
timestamp 1644511149
transform 1 0 18860 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1963_
timestamp 1644511149
transform 1 0 17756 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1964_
timestamp 1644511149
transform 1 0 18216 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1965_
timestamp 1644511149
transform 1 0 17756 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1966_
timestamp 1644511149
transform 1 0 17388 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1967_
timestamp 1644511149
transform 1 0 23552 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1968_
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1969_
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1970_
timestamp 1644511149
transform 1 0 18216 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1971_
timestamp 1644511149
transform 1 0 18216 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _1972_
timestamp 1644511149
transform 1 0 17112 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1973_
timestamp 1644511149
transform 1 0 20516 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1974_
timestamp 1644511149
transform 1 0 21160 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1975_
timestamp 1644511149
transform 1 0 19688 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1976_
timestamp 1644511149
transform 1 0 20608 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1977_
timestamp 1644511149
transform 1 0 20332 0 -1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _1978_
timestamp 1644511149
transform 1 0 13156 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1979_
timestamp 1644511149
transform 1 0 24748 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1980_
timestamp 1644511149
transform 1 0 24380 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1981_
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1982_
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1983_
timestamp 1644511149
transform 1 0 23460 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1984_
timestamp 1644511149
transform 1 0 23644 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1985_
timestamp 1644511149
transform 1 0 23552 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1986_
timestamp 1644511149
transform 1 0 22908 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1987_
timestamp 1644511149
transform 1 0 22080 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1988_
timestamp 1644511149
transform 1 0 22816 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1989_
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1990_
timestamp 1644511149
transform 1 0 22172 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1991_
timestamp 1644511149
transform 1 0 23644 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1992_
timestamp 1644511149
transform 1 0 22816 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1993_
timestamp 1644511149
transform 1 0 23276 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1994_
timestamp 1644511149
transform 1 0 28428 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1995_
timestamp 1644511149
transform 1 0 27324 0 1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1996_
timestamp 1644511149
transform 1 0 26220 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1997_
timestamp 1644511149
transform 1 0 25392 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1998_
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1999_
timestamp 1644511149
transform 1 0 24104 0 -1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _2000_
timestamp 1644511149
transform 1 0 26220 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2001_
timestamp 1644511149
transform 1 0 28244 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2002_
timestamp 1644511149
transform 1 0 27324 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2003_
timestamp 1644511149
transform 1 0 26220 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2004_
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2005_
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2006_
timestamp 1644511149
transform 1 0 28060 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2007_
timestamp 1644511149
transform 1 0 28428 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2008_
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _2009_
timestamp 1644511149
transform 1 0 30636 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2010_
timestamp 1644511149
transform 1 0 29164 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2011_
timestamp 1644511149
transform 1 0 28428 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2012_
timestamp 1644511149
transform 1 0 28060 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2013_
timestamp 1644511149
transform 1 0 28704 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2014_
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2015_
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2016_
timestamp 1644511149
transform 1 0 30268 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2017_
timestamp 1644511149
transform 1 0 30452 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2018_
timestamp 1644511149
transform 1 0 30176 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2019_
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2020_
timestamp 1644511149
transform 1 0 28336 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2021_
timestamp 1644511149
transform 1 0 29072 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2022_
timestamp 1644511149
transform 1 0 27140 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _2023_
timestamp 1644511149
transform 1 0 26220 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2024_
timestamp 1644511149
transform 1 0 27600 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2025_
timestamp 1644511149
transform 1 0 25944 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2026_
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2027_
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2028_
timestamp 1644511149
transform 1 0 26036 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2029_
timestamp 1644511149
transform 1 0 24932 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2030_
timestamp 1644511149
transform 1 0 25024 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2031_
timestamp 1644511149
transform 1 0 24656 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2032_
timestamp 1644511149
transform 1 0 24564 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2033_
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2034_
timestamp 1644511149
transform 1 0 22724 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2035_
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2036_
timestamp 1644511149
transform 1 0 23000 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2037_
timestamp 1644511149
transform 1 0 28428 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2038_
timestamp 1644511149
transform 1 0 29440 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2039_
timestamp 1644511149
transform 1 0 27784 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2040_
timestamp 1644511149
transform 1 0 31004 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _2041_
timestamp 1644511149
transform 1 0 29256 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2042_
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2043_
timestamp 1644511149
transform 1 0 30360 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2044_
timestamp 1644511149
transform 1 0 30452 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2045_
timestamp 1644511149
transform 1 0 28520 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2046_
timestamp 1644511149
transform 1 0 29072 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2047_
timestamp 1644511149
transform 1 0 28520 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2048_
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2049_
timestamp 1644511149
transform 1 0 28520 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2050_
timestamp 1644511149
transform 1 0 30636 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2051_
timestamp 1644511149
transform 1 0 30084 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2052_
timestamp 1644511149
transform 1 0 27784 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2053_
timestamp 1644511149
transform 1 0 29164 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _2054_
timestamp 1644511149
transform 1 0 25944 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _2055_
timestamp 1644511149
transform 1 0 26220 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2056_
timestamp 1644511149
transform 1 0 30268 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2057_
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2058_
timestamp 1644511149
transform 1 0 30268 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2059_
timestamp 1644511149
transform 1 0 28520 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2060_
timestamp 1644511149
transform 1 0 30452 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2061_
timestamp 1644511149
transform 1 0 28520 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2062_
timestamp 1644511149
transform 1 0 28796 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2063_
timestamp 1644511149
transform 1 0 25944 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2064_
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2065_
timestamp 1644511149
transform 1 0 28520 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2066_
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2067_
timestamp 1644511149
transform 1 0 27048 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2068_
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _2069_
timestamp 1644511149
transform 1 0 26956 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2070_
timestamp 1644511149
transform 1 0 26588 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2071_
timestamp 1644511149
transform 1 0 25668 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2072_
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2073_
timestamp 1644511149
transform 1 0 28336 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2074_
timestamp 1644511149
transform 1 0 25392 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2075_
timestamp 1644511149
transform 1 0 24748 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2076_
timestamp 1644511149
transform 1 0 26220 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2077_
timestamp 1644511149
transform 1 0 25024 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2078_
timestamp 1644511149
transform 1 0 25760 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2079_
timestamp 1644511149
transform 1 0 24840 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2080_
timestamp 1644511149
transform 1 0 28704 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2081_
timestamp 1644511149
transform 1 0 26128 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2082_
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _2083_
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2084_
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2085_
timestamp 1644511149
transform 1 0 25944 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2086_
timestamp 1644511149
transform 1 0 25760 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2087_
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2088_
timestamp 1644511149
transform 1 0 25024 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2089_
timestamp 1644511149
transform 1 0 24104 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2090_
timestamp 1644511149
transform 1 0 17572 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2091_
timestamp 1644511149
transform 1 0 21988 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2092_
timestamp 1644511149
transform 1 0 22356 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2093_
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2094_
timestamp 1644511149
transform 1 0 23368 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2095_
timestamp 1644511149
transform 1 0 22356 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2096_
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2097_
timestamp 1644511149
transform 1 0 27416 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _2098_
timestamp 1644511149
transform 1 0 25024 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2099_
timestamp 1644511149
transform 1 0 24564 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2100_
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _2101_
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2102_
timestamp 1644511149
transform 1 0 26588 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2103_
timestamp 1644511149
transform 1 0 25944 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2104_
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2105_
timestamp 1644511149
transform 1 0 26312 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2106_
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2107_
timestamp 1644511149
transform 1 0 27876 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2108_
timestamp 1644511149
transform 1 0 27968 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2109_
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2110_
timestamp 1644511149
transform 1 0 28704 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2111_
timestamp 1644511149
transform 1 0 28152 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2112_
timestamp 1644511149
transform 1 0 28980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2113_
timestamp 1644511149
transform 1 0 29348 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _2114_
timestamp 1644511149
transform 1 0 29992 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2115_
timestamp 1644511149
transform 1 0 29072 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2116_
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2117_
timestamp 1644511149
transform 1 0 30176 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2118_
timestamp 1644511149
transform 1 0 30452 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2119_
timestamp 1644511149
transform 1 0 30084 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2120_
timestamp 1644511149
transform 1 0 30636 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2121_
timestamp 1644511149
transform 1 0 29900 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2122_
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2123_
timestamp 1644511149
transform 1 0 29072 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2124_
timestamp 1644511149
transform 1 0 29992 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2125_
timestamp 1644511149
transform 1 0 30728 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2126_
timestamp 1644511149
transform 1 0 31004 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2127_
timestamp 1644511149
transform 1 0 26036 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _2128_
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2129_
timestamp 1644511149
transform 1 0 30176 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2130_
timestamp 1644511149
transform 1 0 30728 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2131_
timestamp 1644511149
transform 1 0 30084 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2132_
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2133_
timestamp 1644511149
transform 1 0 30636 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2134_
timestamp 1644511149
transform 1 0 30636 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2135_
timestamp 1644511149
transform 1 0 28888 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2136_
timestamp 1644511149
transform 1 0 27232 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2137_
timestamp 1644511149
transform 1 0 26404 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2138_
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2139_
timestamp 1644511149
transform 1 0 28520 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2140_
timestamp 1644511149
transform 1 0 24748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2141_
timestamp 1644511149
transform 1 0 29440 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _2142_
timestamp 1644511149
transform 1 0 28612 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2143_
timestamp 1644511149
transform 1 0 28888 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2144_
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2145_
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2146_
timestamp 1644511149
transform 1 0 28520 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2147_
timestamp 1644511149
transform 1 0 30544 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2148_
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2149_
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2150_
timestamp 1644511149
transform 1 0 30360 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2151_
timestamp 1644511149
transform 1 0 20884 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2152_
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2153_
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2154_
timestamp 1644511149
transform 1 0 28060 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _2155_
timestamp 1644511149
transform 1 0 28336 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2156_
timestamp 1644511149
transform 1 0 27416 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2157_
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _2158_
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2159_
timestamp 1644511149
transform 1 0 29716 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2160_
timestamp 1644511149
transform 1 0 27692 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2161_
timestamp 1644511149
transform 1 0 30452 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2162_
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2163_
timestamp 1644511149
transform 1 0 30452 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2164_
timestamp 1644511149
transform 1 0 30820 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2165_
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2166_
timestamp 1644511149
transform 1 0 30820 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2167_
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2168_
timestamp 1644511149
transform 1 0 28336 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2169_
timestamp 1644511149
transform 1 0 29348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2170_
timestamp 1644511149
transform 1 0 28152 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _2171_
timestamp 1644511149
transform 1 0 27508 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2172_
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2173_
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2174_
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2175_
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2176_
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2177_
timestamp 1644511149
transform 1 0 30636 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2178_
timestamp 1644511149
transform 1 0 28152 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2179_
timestamp 1644511149
transform 1 0 27876 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2180_
timestamp 1644511149
transform 1 0 26220 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _2181_
timestamp 1644511149
transform 1 0 27416 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2182_
timestamp 1644511149
transform 1 0 25944 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2183_
timestamp 1644511149
transform 1 0 24564 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _2184_
timestamp 1644511149
transform 1 0 26404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2185_
timestamp 1644511149
transform 1 0 25300 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2186_
timestamp 1644511149
transform 1 0 25760 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2187_
timestamp 1644511149
transform 1 0 24748 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2188_
timestamp 1644511149
transform 1 0 24656 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2189_
timestamp 1644511149
transform 1 0 25116 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2190_
timestamp 1644511149
transform 1 0 23368 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2191_
timestamp 1644511149
transform 1 0 24380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2192_
timestamp 1644511149
transform 1 0 23460 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2193_
timestamp 1644511149
transform 1 0 22540 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _2194_
timestamp 1644511149
transform 1 0 23184 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2195_
timestamp 1644511149
transform 1 0 23368 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2196_
timestamp 1644511149
transform 1 0 23828 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _2197_
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _2198_
timestamp 1644511149
transform 1 0 19228 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2199_
timestamp 1644511149
transform 1 0 22080 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2200_
timestamp 1644511149
transform 1 0 22448 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2201_
timestamp 1644511149
transform 1 0 22080 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2202_
timestamp 1644511149
transform 1 0 19504 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2203_
timestamp 1644511149
transform 1 0 23092 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2204_
timestamp 1644511149
transform 1 0 22264 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2205_
timestamp 1644511149
transform 1 0 20976 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2206_
timestamp 1644511149
transform 1 0 20792 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2207_
timestamp 1644511149
transform 1 0 21068 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2208_
timestamp 1644511149
transform 1 0 20424 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2209_
timestamp 1644511149
transform 1 0 19872 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2210_
timestamp 1644511149
transform 1 0 19872 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2211_
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2212_
timestamp 1644511149
transform 1 0 19964 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2213_
timestamp 1644511149
transform 1 0 16928 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _2214_
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2215_
timestamp 1644511149
transform 1 0 18124 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2216_
timestamp 1644511149
transform 1 0 18216 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2217_
timestamp 1644511149
transform 1 0 18032 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2218_
timestamp 1644511149
transform 1 0 18216 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2219_
timestamp 1644511149
transform 1 0 18124 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2220_
timestamp 1644511149
transform 1 0 18216 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2221_
timestamp 1644511149
transform 1 0 13248 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2222_
timestamp 1644511149
transform 1 0 15364 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _2223_
timestamp 1644511149
transform 1 0 16836 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2224_
timestamp 1644511149
transform 1 0 16652 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2225_
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2226_
timestamp 1644511149
transform 1 0 15640 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2227_
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _2228_
timestamp 1644511149
transform 1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2229_
timestamp 1644511149
transform 1 0 14628 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2230_
timestamp 1644511149
transform 1 0 14720 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2231_
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2232_
timestamp 1644511149
transform 1 0 13340 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2233_
timestamp 1644511149
transform 1 0 14076 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2234_
timestamp 1644511149
transform 1 0 13064 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2235_
timestamp 1644511149
transform 1 0 12696 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _2236_
timestamp 1644511149
transform 1 0 15180 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2237_
timestamp 1644511149
transform 1 0 12604 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2238_
timestamp 1644511149
transform 1 0 13984 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2239_
timestamp 1644511149
transform 1 0 11776 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2240_
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _2241_
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2242_
timestamp 1644511149
transform 1 0 13432 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2243_
timestamp 1644511149
transform 1 0 12236 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2244_
timestamp 1644511149
transform 1 0 14536 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2245_
timestamp 1644511149
transform 1 0 12328 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2246_
timestamp 1644511149
transform 1 0 13616 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2247_
timestamp 1644511149
transform 1 0 15640 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2248_
timestamp 1644511149
transform 1 0 15272 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _2249_
timestamp 1644511149
transform 1 0 15364 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2250_
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2251_
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2252_
timestamp 1644511149
transform 1 0 16468 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2253_
timestamp 1644511149
transform 1 0 13248 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _2254_
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2255_
timestamp 1644511149
transform 1 0 18952 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2256_
timestamp 1644511149
transform 1 0 18032 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2257_
timestamp 1644511149
transform 1 0 20056 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2258_
timestamp 1644511149
transform 1 0 19320 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2259_
timestamp 1644511149
transform 1 0 20148 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2260_
timestamp 1644511149
transform 1 0 19320 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2261_
timestamp 1644511149
transform 1 0 13984 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2262_
timestamp 1644511149
transform 1 0 22632 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _2263_
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _2264_
timestamp 1644511149
transform 1 0 22448 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2265_
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2266_
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2267_
timestamp 1644511149
transform 1 0 12604 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2268_
timestamp 1644511149
transform 1 0 15272 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2269_
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2270_
timestamp 1644511149
transform 1 0 8648 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2271_
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2272_
timestamp 1644511149
transform 1 0 21252 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2273_
timestamp 1644511149
transform 1 0 24196 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2274_
timestamp 1644511149
transform 1 0 22632 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2275_
timestamp 1644511149
transform 1 0 22724 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _2276_
timestamp 1644511149
transform 1 0 23552 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2277_
timestamp 1644511149
transform 1 0 25208 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _2278_
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2279_
timestamp 1644511149
transform 1 0 26128 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2280_
timestamp 1644511149
transform 1 0 25484 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2281_
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2282_
timestamp 1644511149
transform 1 0 20700 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2283_
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2284_
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2285_
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2286_
timestamp 1644511149
transform 1 0 25760 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2287_
timestamp 1644511149
transform 1 0 25760 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2288_
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2289_
timestamp 1644511149
transform 1 0 25944 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2290_
timestamp 1644511149
transform 1 0 24472 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _2291_
timestamp 1644511149
transform 1 0 25760 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2292_
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _2293_
timestamp 1644511149
transform 1 0 13156 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2294_
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2295_
timestamp 1644511149
transform 1 0 23092 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2296_
timestamp 1644511149
transform 1 0 18400 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2297_
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2298_
timestamp 1644511149
transform 1 0 24012 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2299_
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2300_
timestamp 1644511149
transform 1 0 24196 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2301_
timestamp 1644511149
transform 1 0 18676 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2302_
timestamp 1644511149
transform 1 0 24656 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2303_
timestamp 1644511149
transform 1 0 23368 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2304_
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2305_
timestamp 1644511149
transform 1 0 23368 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _2306_
timestamp 1644511149
transform 1 0 6532 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2307_
timestamp 1644511149
transform 1 0 23184 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2308_
timestamp 1644511149
transform 1 0 23368 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2309_
timestamp 1644511149
transform 1 0 22264 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2310_
timestamp 1644511149
transform 1 0 21804 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2311_
timestamp 1644511149
transform 1 0 22356 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2312_
timestamp 1644511149
transform 1 0 22080 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2313_
timestamp 1644511149
transform 1 0 13156 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2314_
timestamp 1644511149
transform 1 0 17940 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _2315_
timestamp 1644511149
transform 1 0 17940 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _2316_
timestamp 1644511149
transform 1 0 4140 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _2317_
timestamp 1644511149
transform 1 0 18952 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _2318_
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2319_
timestamp 1644511149
transform 1 0 4968 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2320_
timestamp 1644511149
transform 1 0 8464 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2321_
timestamp 1644511149
transform 1 0 4508 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _2322_
timestamp 1644511149
transform 1 0 13892 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _2323_
timestamp 1644511149
transform 1 0 10212 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2324_
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2325_
timestamp 1644511149
transform 1 0 5520 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2326_
timestamp 1644511149
transform 1 0 5152 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2327_
timestamp 1644511149
transform 1 0 14996 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _2328_
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _2329_
timestamp 1644511149
transform 1 0 7176 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2330_
timestamp 1644511149
transform 1 0 5520 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2331_
timestamp 1644511149
transform 1 0 5244 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _2332_
timestamp 1644511149
transform 1 0 5612 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2333_
timestamp 1644511149
transform 1 0 4508 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2334_
timestamp 1644511149
transform 1 0 4968 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2335_
timestamp 1644511149
transform 1 0 4416 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2336_
timestamp 1644511149
transform 1 0 3956 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2337_
timestamp 1644511149
transform 1 0 4232 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2338_
timestamp 1644511149
transform 1 0 3956 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2339_
timestamp 1644511149
transform 1 0 4324 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2340_
timestamp 1644511149
transform 1 0 5336 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2341_
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2342_
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2343_
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2344_
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2345_
timestamp 1644511149
transform 1 0 3036 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _2346_
timestamp 1644511149
transform 1 0 1932 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2347_
timestamp 1644511149
transform 1 0 1472 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2348_
timestamp 1644511149
transform 1 0 1932 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2349_
timestamp 1644511149
transform 1 0 1564 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2350_
timestamp 1644511149
transform 1 0 4324 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2351_
timestamp 1644511149
transform 1 0 1656 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2352_
timestamp 1644511149
transform 1 0 4508 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _2353_
timestamp 1644511149
transform 1 0 7452 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2354_
timestamp 1644511149
transform 1 0 3220 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2355_
timestamp 1644511149
transform 1 0 2760 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2356_
timestamp 1644511149
transform 1 0 2024 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2357_
timestamp 1644511149
transform 1 0 1748 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2358_
timestamp 1644511149
transform 1 0 11316 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2359_
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _2360_
timestamp 1644511149
transform 1 0 2116 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2361_
timestamp 1644511149
transform 1 0 1840 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2362_
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2363_
timestamp 1644511149
transform 1 0 2760 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2364_
timestamp 1644511149
transform 1 0 6900 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2365_
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2366_
timestamp 1644511149
transform 1 0 8096 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2367_
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2368_
timestamp 1644511149
transform 1 0 7636 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2369_
timestamp 1644511149
transform 1 0 9476 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2370_
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2371_
timestamp 1644511149
transform 1 0 3312 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2372_
timestamp 1644511149
transform 1 0 1748 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2373_
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2374_
timestamp 1644511149
transform 1 0 2024 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2375_
timestamp 1644511149
transform 1 0 2116 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2376_
timestamp 1644511149
transform 1 0 2668 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2377_
timestamp 1644511149
transform 1 0 2300 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2378_
timestamp 1644511149
transform 1 0 3220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _2379_
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2380_
timestamp 1644511149
transform 1 0 3036 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2381_
timestamp 1644511149
transform 1 0 3128 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2382_
timestamp 1644511149
transform 1 0 1932 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2383_
timestamp 1644511149
transform 1 0 2116 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2384_
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2385_
timestamp 1644511149
transform 1 0 1932 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2386_
timestamp 1644511149
transform 1 0 1840 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2387_
timestamp 1644511149
transform 1 0 4600 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2388_
timestamp 1644511149
transform 1 0 2024 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2389_
timestamp 1644511149
transform 1 0 1748 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2390_
timestamp 1644511149
transform 1 0 2024 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2391_
timestamp 1644511149
transform 1 0 1748 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _2392_
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2393_
timestamp 1644511149
transform 1 0 3496 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2394_
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2395_
timestamp 1644511149
transform 1 0 4600 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2396_
timestamp 1644511149
transform 1 0 5060 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2397_
timestamp 1644511149
transform 1 0 9016 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2398_
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2399_
timestamp 1644511149
transform 1 0 7912 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2400_
timestamp 1644511149
transform 1 0 7728 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2401_
timestamp 1644511149
transform 1 0 2116 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2402_
timestamp 1644511149
transform 1 0 4508 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2403_
timestamp 1644511149
transform 1 0 4876 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2404_
timestamp 1644511149
transform 1 0 5060 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _2405_
timestamp 1644511149
transform 1 0 4784 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2406_
timestamp 1644511149
transform 1 0 5888 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2407_
timestamp 1644511149
transform 1 0 4692 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2408_
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2409_
timestamp 1644511149
transform 1 0 6624 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _2410_
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2411_
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2412_
timestamp 1644511149
transform 1 0 8096 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2413_
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2414_
timestamp 1644511149
transform 1 0 5336 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2415_
timestamp 1644511149
transform 1 0 5152 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2416_
timestamp 1644511149
transform 1 0 5428 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2417_
timestamp 1644511149
transform 1 0 8464 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2418_
timestamp 1644511149
transform 1 0 6440 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2419_
timestamp 1644511149
transform 1 0 7268 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2420_
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2421_
timestamp 1644511149
transform 1 0 2760 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2422_
timestamp 1644511149
transform 1 0 7912 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _2423_
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2424_
timestamp 1644511149
transform 1 0 6348 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2425_
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2426_
timestamp 1644511149
transform 1 0 9200 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2427_
timestamp 1644511149
transform 1 0 10304 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2428_
timestamp 1644511149
transform 1 0 9016 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2429_
timestamp 1644511149
transform 1 0 10212 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2430_
timestamp 1644511149
transform 1 0 10764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2431_
timestamp 1644511149
transform 1 0 10120 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2432_
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2433_
timestamp 1644511149
transform 1 0 9200 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2434_
timestamp 1644511149
transform 1 0 10304 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2435_
timestamp 1644511149
transform 1 0 10672 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _2436_
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2437_
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2438_
timestamp 1644511149
transform 1 0 10212 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2439_
timestamp 1644511149
transform 1 0 12236 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2440_
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2441_
timestamp 1644511149
transform 1 0 10396 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2442_
timestamp 1644511149
transform 1 0 9660 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2443_
timestamp 1644511149
transform 1 0 9292 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2444_
timestamp 1644511149
transform 1 0 10764 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _2445_
timestamp 1644511149
transform 1 0 10212 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2446_
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2447_
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2448_
timestamp 1644511149
transform 1 0 10488 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _2449_
timestamp 1644511149
transform 1 0 5612 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2450_
timestamp 1644511149
transform 1 0 12328 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2451_
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2452_
timestamp 1644511149
transform 1 0 10304 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2453_
timestamp 1644511149
transform 1 0 9292 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2454_
timestamp 1644511149
transform 1 0 9844 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2455_
timestamp 1644511149
transform 1 0 9292 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2456_
timestamp 1644511149
transform 1 0 13616 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _2457_
timestamp 1644511149
transform 1 0 12512 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _2458_
timestamp 1644511149
transform 1 0 12328 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2459_
timestamp 1644511149
transform 1 0 1472 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _2460_
timestamp 1644511149
transform 1 0 11592 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2461_
timestamp 1644511149
transform 1 0 11868 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _2462_
timestamp 1644511149
transform 1 0 12880 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2463_
timestamp 1644511149
transform 1 0 11960 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2464_
timestamp 1644511149
transform 1 0 20884 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _2465_
timestamp 1644511149
transform 1 0 17848 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _2466_
timestamp 1644511149
transform 1 0 17572 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2467_
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2468_
timestamp 1644511149
transform 1 0 10948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2469_
timestamp 1644511149
transform 1 0 13248 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _2470_
timestamp 1644511149
transform 1 0 4324 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2471_
timestamp 1644511149
transform 1 0 12604 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2472_
timestamp 1644511149
transform 1 0 14352 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2473_
timestamp 1644511149
transform 1 0 11500 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2474_
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2475_
timestamp 1644511149
transform 1 0 11776 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2476_
timestamp 1644511149
transform 1 0 11592 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2477_
timestamp 1644511149
transform 1 0 13156 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2478_
timestamp 1644511149
transform 1 0 10212 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2479_
timestamp 1644511149
transform 1 0 9292 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2480_
timestamp 1644511149
transform 1 0 10120 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2481_
timestamp 1644511149
transform 1 0 9200 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2482_
timestamp 1644511149
transform 1 0 19228 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2483_
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _2484_
timestamp 1644511149
transform 1 0 7544 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2485_
timestamp 1644511149
transform 1 0 10028 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2486_
timestamp 1644511149
transform 1 0 9108 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2487_
timestamp 1644511149
transform 1 0 9844 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2488_
timestamp 1644511149
transform 1 0 11224 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2489_
timestamp 1644511149
transform 1 0 9844 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2490_
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2491_
timestamp 1644511149
transform 1 0 18400 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2492_
timestamp 1644511149
transform 1 0 14352 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2493_
timestamp 1644511149
transform 1 0 10764 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2494_
timestamp 1644511149
transform 1 0 10764 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2495_
timestamp 1644511149
transform 1 0 14444 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2496_
timestamp 1644511149
transform 1 0 11500 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2497_
timestamp 1644511149
transform 1 0 10304 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2498_
timestamp 1644511149
transform 1 0 12420 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2499_
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2500_
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _2501_
timestamp 1644511149
transform 1 0 12880 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2502_
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2503_
timestamp 1644511149
transform 1 0 11868 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2504_
timestamp 1644511149
transform 1 0 12144 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2505_
timestamp 1644511149
transform 1 0 14628 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2506_
timestamp 1644511149
transform 1 0 12420 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2507_
timestamp 1644511149
transform 1 0 11500 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2508_
timestamp 1644511149
transform 1 0 16468 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2509_
timestamp 1644511149
transform 1 0 13340 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2510_
timestamp 1644511149
transform 1 0 15732 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2511_
timestamp 1644511149
transform 1 0 16652 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2512_
timestamp 1644511149
transform 1 0 14168 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2513_
timestamp 1644511149
transform 1 0 12052 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2514_
timestamp 1644511149
transform 1 0 12972 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2515_
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2516_
timestamp 1644511149
transform 1 0 13524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2517_
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2518_
timestamp 1644511149
transform 1 0 15364 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _2519_
timestamp 1644511149
transform 1 0 12972 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _2520_
timestamp 1644511149
transform 1 0 17388 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2521_
timestamp 1644511149
transform 1 0 14904 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2522_
timestamp 1644511149
transform 1 0 13984 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2523_
timestamp 1644511149
transform 1 0 14444 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2524_
timestamp 1644511149
transform 1 0 14260 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2525_
timestamp 1644511149
transform 1 0 14168 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2526_
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2527_
timestamp 1644511149
transform 1 0 15272 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2528_
timestamp 1644511149
transform 1 0 15456 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2529_
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2530_
timestamp 1644511149
transform 1 0 15272 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2531_
timestamp 1644511149
transform 1 0 19780 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2532_
timestamp 1644511149
transform 1 0 18584 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _2533_
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2534_
timestamp 1644511149
transform 1 0 17480 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2535_
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2536_
timestamp 1644511149
transform 1 0 17480 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2537_
timestamp 1644511149
transform 1 0 17112 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2538_
timestamp 1644511149
transform 1 0 18952 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2539_
timestamp 1644511149
transform 1 0 19136 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2540_
timestamp 1644511149
transform 1 0 17572 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2541_
timestamp 1644511149
transform 1 0 17848 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _2542_
timestamp 1644511149
transform 1 0 19872 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2543_
timestamp 1644511149
transform 1 0 20792 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2544_
timestamp 1644511149
transform 1 0 20608 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2545_
timestamp 1644511149
transform 1 0 20884 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2546_
timestamp 1644511149
transform 1 0 20976 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2547_
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2548_
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2549_
timestamp 1644511149
transform 1 0 22080 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2550_
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _2551_
timestamp 1644511149
transform 1 0 22080 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2552_
timestamp 1644511149
transform 1 0 20884 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2553_
timestamp 1644511149
transform 1 0 20792 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2554_
timestamp 1644511149
transform 1 0 21620 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2555_
timestamp 1644511149
transform 1 0 20792 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2556_
timestamp 1644511149
transform 1 0 23184 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2557_
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2558_
timestamp 1644511149
transform 1 0 19228 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2559_
timestamp 1644511149
transform 1 0 12512 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2560_
timestamp 1644511149
transform 1 0 19412 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2561_
timestamp 1644511149
transform 1 0 10672 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2562_
timestamp 1644511149
transform 1 0 20148 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2563_
timestamp 1644511149
transform 1 0 19872 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2564_
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2565_
timestamp 1644511149
transform 1 0 18032 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2566_
timestamp 1644511149
transform 1 0 18400 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2567_
timestamp 1644511149
transform 1 0 17664 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2568_
timestamp 1644511149
transform 1 0 19228 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2569_
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2570_
timestamp 1644511149
transform 1 0 19780 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _2571_
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2572_
timestamp 1644511149
transform 1 0 17664 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2573_
timestamp 1644511149
transform 1 0 17664 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2574_
timestamp 1644511149
transform 1 0 9108 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2575_
timestamp 1644511149
transform 1 0 17296 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2576_
timestamp 1644511149
transform 1 0 16928 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2577_
timestamp 1644511149
transform 1 0 18400 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2578_
timestamp 1644511149
transform 1 0 17756 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2579_
timestamp 1644511149
transform 1 0 18032 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2580_
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2581_
timestamp 1644511149
transform 1 0 16928 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2582_
timestamp 1644511149
transform 1 0 16744 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2583_
timestamp 1644511149
transform 1 0 25760 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2584_
timestamp 1644511149
transform 1 0 19504 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _2585_
timestamp 1644511149
transform 1 0 21988 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2586_
timestamp 1644511149
transform 1 0 20700 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2587_
timestamp 1644511149
transform 1 0 24932 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2588_
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2589_
timestamp 1644511149
transform 1 0 20424 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2590_
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2591_
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2592_
timestamp 1644511149
transform 1 0 23092 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2593_
timestamp 1644511149
transform 1 0 21896 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2594_
timestamp 1644511149
transform 1 0 20424 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2595_
timestamp 1644511149
transform 1 0 19504 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2596_
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2597_
timestamp 1644511149
transform 1 0 16468 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__o21ba_1  _2598_
timestamp 1644511149
transform 1 0 20148 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2599_
timestamp 1644511149
transform 1 0 19780 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2600_
timestamp 1644511149
transform 1 0 17112 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2601_
timestamp 1644511149
transform 1 0 16744 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2602_
timestamp 1644511149
transform 1 0 19412 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2603_
timestamp 1644511149
transform 1 0 19504 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2604_
timestamp 1644511149
transform 1 0 19320 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2605_
timestamp 1644511149
transform 1 0 18216 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2606_
timestamp 1644511149
transform 1 0 16836 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2607_
timestamp 1644511149
transform 1 0 19596 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2608_
timestamp 1644511149
transform 1 0 20332 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2609_
timestamp 1644511149
transform 1 0 17480 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2610_
timestamp 1644511149
transform 1 0 16836 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2611_
timestamp 1644511149
transform 1 0 10856 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2612_
timestamp 1644511149
transform 1 0 15824 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2613_
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2614_
timestamp 1644511149
transform 1 0 15272 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _2615_
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2616_
timestamp 1644511149
transform 1 0 14904 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2617_
timestamp 1644511149
transform 1 0 14628 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2618_
timestamp 1644511149
transform 1 0 15364 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2619_
timestamp 1644511149
transform 1 0 15548 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2620_
timestamp 1644511149
transform 1 0 14812 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2621_
timestamp 1644511149
transform 1 0 15548 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2622_
timestamp 1644511149
transform 1 0 15456 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2623_
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2624_
timestamp 1644511149
transform 1 0 16468 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _2625_
timestamp 1644511149
transform 1 0 14260 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2626_
timestamp 1644511149
transform 1 0 15088 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2627_
timestamp 1644511149
transform 1 0 14904 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2628_
timestamp 1644511149
transform 1 0 14168 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2629_
timestamp 1644511149
transform 1 0 15088 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2630_
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2631_
timestamp 1644511149
transform 1 0 15088 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2632_
timestamp 1644511149
transform 1 0 14904 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2633_
timestamp 1644511149
transform 1 0 19872 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _2634_
timestamp 1644511149
transform 1 0 20608 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _2635_
timestamp 1644511149
transform 1 0 20056 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _2636_
timestamp 1644511149
transform 1 0 12604 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _2637_
timestamp 1644511149
transform 1 0 14076 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _2638_
timestamp 1644511149
transform 1 0 8280 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2639_
timestamp 1644511149
transform 1 0 6532 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2640_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2641_
timestamp 1644511149
transform 1 0 9752 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2642_
timestamp 1644511149
transform 1 0 9292 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2643_
timestamp 1644511149
transform 1 0 8096 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2644_
timestamp 1644511149
transform 1 0 6716 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2645_
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2646_
timestamp 1644511149
transform 1 0 4416 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2647_
timestamp 1644511149
transform 1 0 4232 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2648_
timestamp 1644511149
transform 1 0 1840 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2649_
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2650_
timestamp 1644511149
transform 1 0 1472 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2651_
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2652_
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2653_
timestamp 1644511149
transform 1 0 3220 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2654_
timestamp 1644511149
transform 1 0 4416 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2655_
timestamp 1644511149
transform 1 0 4508 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2656_
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2657_
timestamp 1644511149
transform 1 0 6900 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2658_
timestamp 1644511149
transform 1 0 7636 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2659_ pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 -1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2660_
timestamp 1644511149
transform 1 0 10856 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2661_
timestamp 1644511149
transform 1 0 20792 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2662_
timestamp 1644511149
transform 1 0 5520 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2663_
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2664_
timestamp 1644511149
transform 1 0 3772 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2665_
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2666_
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2667_
timestamp 1644511149
transform 1 0 1840 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2668_
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2669_
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2670_
timestamp 1644511149
transform 1 0 1840 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2671_
timestamp 1644511149
transform 1 0 3772 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2672_
timestamp 1644511149
transform 1 0 4416 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2673_
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2674_
timestamp 1644511149
transform 1 0 6256 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2675_
timestamp 1644511149
transform 1 0 6992 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2676_
timestamp 1644511149
transform 1 0 6992 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2677_
timestamp 1644511149
transform 1 0 8372 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2678_
timestamp 1644511149
transform 1 0 9384 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2679_
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2680_
timestamp 1644511149
transform 1 0 9476 0 -1 38080
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2681_
timestamp 1644511149
transform 1 0 9844 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2682_
timestamp 1644511149
transform 1 0 22540 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2683_
timestamp 1644511149
transform 1 0 12144 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2684_
timestamp 1644511149
transform 1 0 12144 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2685_
timestamp 1644511149
transform 1 0 11868 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2686_
timestamp 1644511149
transform 1 0 11592 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2687_
timestamp 1644511149
transform 1 0 12052 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2688_
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2689_
timestamp 1644511149
transform 1 0 13984 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2690_
timestamp 1644511149
transform 1 0 14536 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2691_
timestamp 1644511149
transform 1 0 15916 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2692_
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2693_
timestamp 1644511149
transform 1 0 18492 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2694_
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2695_
timestamp 1644511149
transform 1 0 18216 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2696_
timestamp 1644511149
transform 1 0 17020 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2697_
timestamp 1644511149
transform 1 0 16836 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2698_
timestamp 1644511149
transform 1 0 18676 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2699_
timestamp 1644511149
transform 1 0 18676 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2700_
timestamp 1644511149
transform 1 0 19320 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2701_
timestamp 1644511149
transform 1 0 19780 0 -1 38080
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2702_
timestamp 1644511149
transform 1 0 19780 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2703_
timestamp 1644511149
transform 1 0 22816 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2704_
timestamp 1644511149
transform 1 0 21620 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2705_
timestamp 1644511149
transform 1 0 20608 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2706_
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2707_
timestamp 1644511149
transform 1 0 22448 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2708_
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2709_
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2710_
timestamp 1644511149
transform 1 0 25024 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2711_
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2712_
timestamp 1644511149
transform 1 0 28796 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2713_
timestamp 1644511149
transform 1 0 27600 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2714_
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2715_
timestamp 1644511149
transform 1 0 29900 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2716_
timestamp 1644511149
transform 1 0 29900 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2717_
timestamp 1644511149
transform 1 0 28060 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2718_
timestamp 1644511149
transform 1 0 27232 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2719_
timestamp 1644511149
transform 1 0 25760 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2720_
timestamp 1644511149
transform 1 0 24380 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2721_
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2722_
timestamp 1644511149
transform 1 0 22080 0 1 33728
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2723_
timestamp 1644511149
transform 1 0 22448 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2724_
timestamp 1644511149
transform 1 0 29808 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2725_
timestamp 1644511149
transform 1 0 29900 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2726_
timestamp 1644511149
transform 1 0 29900 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2727_
timestamp 1644511149
transform 1 0 27600 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2728_
timestamp 1644511149
transform 1 0 29900 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2729_
timestamp 1644511149
transform 1 0 29900 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2730_
timestamp 1644511149
transform 1 0 29900 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2731_
timestamp 1644511149
transform 1 0 29900 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2732_
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2733_
timestamp 1644511149
transform 1 0 27600 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2734_
timestamp 1644511149
transform 1 0 28244 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2735_
timestamp 1644511149
transform 1 0 26312 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2736_
timestamp 1644511149
transform 1 0 26496 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2737_
timestamp 1644511149
transform 1 0 24380 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2738_
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2739_
timestamp 1644511149
transform 1 0 26496 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2740_
timestamp 1644511149
transform 1 0 26680 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2741_
timestamp 1644511149
transform 1 0 25484 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2742_
timestamp 1644511149
transform 1 0 24472 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2743_
timestamp 1644511149
transform 1 0 24380 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2744_
timestamp 1644511149
transform 1 0 24104 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2745_
timestamp 1644511149
transform 1 0 22356 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2746_
timestamp 1644511149
transform 1 0 24196 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2747_
timestamp 1644511149
transform 1 0 25576 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2748_
timestamp 1644511149
transform 1 0 25852 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2749_
timestamp 1644511149
transform 1 0 26312 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2750_
timestamp 1644511149
transform 1 0 27784 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2751_
timestamp 1644511149
transform 1 0 27600 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2752_
timestamp 1644511149
transform 1 0 27600 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2753_
timestamp 1644511149
transform 1 0 29624 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2754_
timestamp 1644511149
transform 1 0 29900 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2755_
timestamp 1644511149
transform 1 0 29900 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2756_
timestamp 1644511149
transform 1 0 29900 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2757_
timestamp 1644511149
transform 1 0 29900 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2758_
timestamp 1644511149
transform 1 0 29900 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2759_
timestamp 1644511149
transform 1 0 29808 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2760_
timestamp 1644511149
transform 1 0 27600 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2761_
timestamp 1644511149
transform 1 0 28336 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2762_
timestamp 1644511149
transform 1 0 28244 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2763_
timestamp 1644511149
transform 1 0 28704 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2764_
timestamp 1644511149
transform 1 0 29808 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2765_
timestamp 1644511149
transform 1 0 29900 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2766_
timestamp 1644511149
transform 1 0 20240 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2767_
timestamp 1644511149
transform 1 0 27600 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2768_
timestamp 1644511149
transform 1 0 27876 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2769_
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2770_
timestamp 1644511149
transform 1 0 29900 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2771_
timestamp 1644511149
transform 1 0 29900 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2772_
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2773_
timestamp 1644511149
transform 1 0 27692 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2774_
timestamp 1644511149
transform 1 0 29348 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2775_
timestamp 1644511149
transform 1 0 29256 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2776_
timestamp 1644511149
transform 1 0 27416 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2777_
timestamp 1644511149
transform 1 0 26312 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2778_
timestamp 1644511149
transform 1 0 24472 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2779_
timestamp 1644511149
transform 1 0 24012 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2780_
timestamp 1644511149
transform 1 0 24564 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2781_
timestamp 1644511149
transform 1 0 23920 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2782_
timestamp 1644511149
transform 1 0 23184 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2783_
timestamp 1644511149
transform 1 0 21896 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2784_
timestamp 1644511149
transform 1 0 21344 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2785_
timestamp 1644511149
transform 1 0 21804 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2786_
timestamp 1644511149
transform 1 0 21988 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2787_
timestamp 1644511149
transform 1 0 19872 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2788_
timestamp 1644511149
transform 1 0 19872 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2789_
timestamp 1644511149
transform 1 0 18124 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2790_
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2791_
timestamp 1644511149
transform 1 0 18032 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2792_
timestamp 1644511149
transform 1 0 16376 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2793_
timestamp 1644511149
transform 1 0 14536 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2794_
timestamp 1644511149
transform 1 0 14536 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2795_
timestamp 1644511149
transform 1 0 12788 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2796_
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2797_
timestamp 1644511149
transform 1 0 11500 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2798_
timestamp 1644511149
transform 1 0 11500 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2799_
timestamp 1644511149
transform 1 0 11316 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2800_
timestamp 1644511149
transform 1 0 11592 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2801_
timestamp 1644511149
transform 1 0 12972 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2802_
timestamp 1644511149
transform 1 0 14628 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2803_
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2804_
timestamp 1644511149
transform 1 0 18032 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2805_
timestamp 1644511149
transform 1 0 19320 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2806_
timestamp 1644511149
transform 1 0 20240 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2807_
timestamp 1644511149
transform 1 0 11500 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2808_
timestamp 1644511149
transform 1 0 20792 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2809_
timestamp 1644511149
transform 1 0 19964 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2810_
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2811_
timestamp 1644511149
transform 1 0 21988 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2812_
timestamp 1644511149
transform 1 0 26220 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2813_
timestamp 1644511149
transform 1 0 24932 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2814_
timestamp 1644511149
transform 1 0 26680 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2815_
timestamp 1644511149
transform 1 0 26680 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2816_
timestamp 1644511149
transform 1 0 25760 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2817_
timestamp 1644511149
transform 1 0 25576 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2818_
timestamp 1644511149
transform 1 0 22540 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2819_
timestamp 1644511149
transform 1 0 24196 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2820_
timestamp 1644511149
transform 1 0 24748 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2821_
timestamp 1644511149
transform 1 0 24932 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2822_
timestamp 1644511149
transform 1 0 23092 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2823_
timestamp 1644511149
transform 1 0 23184 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2824_
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2825_
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2826_
timestamp 1644511149
transform 1 0 17940 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2827_
timestamp 1644511149
transform 1 0 14076 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2828_
timestamp 1644511149
transform 1 0 9568 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2829_
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2830_
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2831_
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2832_
timestamp 1644511149
transform 1 0 4048 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2833_
timestamp 1644511149
transform 1 0 3772 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2834_
timestamp 1644511149
transform 1 0 3864 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2835_
timestamp 1644511149
transform 1 0 2852 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2836_
timestamp 1644511149
transform 1 0 4140 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2837_
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2838_
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2839_
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2840_
timestamp 1644511149
transform 1 0 1840 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2841_
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2842_
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2843_
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2844_
timestamp 1644511149
transform 1 0 5612 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2845_
timestamp 1644511149
transform 1 0 7636 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2846_
timestamp 1644511149
transform 1 0 2668 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2847_
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2848_
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2849_
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2850_
timestamp 1644511149
transform 1 0 1564 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2851_
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2852_
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2853_
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2854_
timestamp 1644511149
transform 1 0 2760 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2855_
timestamp 1644511149
transform 1 0 4416 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2856_
timestamp 1644511149
transform 1 0 5704 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2857_
timestamp 1644511149
transform 1 0 7820 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2858_
timestamp 1644511149
transform 1 0 4508 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2859_
timestamp 1644511149
transform 1 0 4140 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2860_
timestamp 1644511149
transform 1 0 4140 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2861_
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2862_
timestamp 1644511149
transform 1 0 5060 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2863_
timestamp 1644511149
transform 1 0 4232 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2864_
timestamp 1644511149
transform 1 0 7176 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2865_
timestamp 1644511149
transform 1 0 4416 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2866_
timestamp 1644511149
transform 1 0 4416 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2867_
timestamp 1644511149
transform 1 0 9476 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2868_
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2869_
timestamp 1644511149
transform 1 0 9568 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2870_
timestamp 1644511149
transform 1 0 7360 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2871_
timestamp 1644511149
transform 1 0 9568 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2872_
timestamp 1644511149
transform 1 0 10120 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2873_
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2874_
timestamp 1644511149
transform 1 0 9752 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2875_
timestamp 1644511149
transform 1 0 10488 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2876_
timestamp 1644511149
transform 1 0 10488 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2877_
timestamp 1644511149
transform 1 0 10212 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2878_
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2879_
timestamp 1644511149
transform 1 0 11776 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2880_
timestamp 1644511149
transform 1 0 14444 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2881_
timestamp 1644511149
transform 1 0 19780 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2882_
timestamp 1644511149
transform 1 0 12144 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2883_
timestamp 1644511149
transform 1 0 17020 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2884_
timestamp 1644511149
transform 1 0 11868 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2885_
timestamp 1644511149
transform 1 0 12512 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2886_
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2887_
timestamp 1644511149
transform 1 0 11224 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2888_
timestamp 1644511149
transform 1 0 8924 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2889_
timestamp 1644511149
transform 1 0 9384 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2890_
timestamp 1644511149
transform 1 0 8188 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2891_
timestamp 1644511149
transform 1 0 9384 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2892_
timestamp 1644511149
transform 1 0 7084 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2893_
timestamp 1644511149
transform 1 0 7544 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2894_
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2895_
timestamp 1644511149
transform 1 0 9660 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2896_
timestamp 1644511149
transform 1 0 12788 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2897_
timestamp 1644511149
transform 1 0 11040 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2898_
timestamp 1644511149
transform 1 0 11684 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2899_
timestamp 1644511149
transform 1 0 12788 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2900_
timestamp 1644511149
transform 1 0 12144 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2901_
timestamp 1644511149
transform 1 0 10304 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2902_
timestamp 1644511149
transform 1 0 13524 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2903_
timestamp 1644511149
transform 1 0 14628 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2904_
timestamp 1644511149
transform 1 0 13156 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2905_
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2906_
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2907_
timestamp 1644511149
transform 1 0 15088 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2908_
timestamp 1644511149
transform 1 0 17020 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2909_
timestamp 1644511149
transform 1 0 16468 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2910_
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2911_
timestamp 1644511149
transform 1 0 16836 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2912_
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2913_
timestamp 1644511149
transform 1 0 20608 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2914_
timestamp 1644511149
transform 1 0 22172 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2915_
timestamp 1644511149
transform 1 0 20792 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2916_
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2917_
timestamp 1644511149
transform 1 0 21804 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2918_
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2919_
timestamp 1644511149
transform 1 0 19780 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2920_
timestamp 1644511149
transform 1 0 17388 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2921_
timestamp 1644511149
transform 1 0 17296 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2922_
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2923_
timestamp 1644511149
transform 1 0 16836 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2924_
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2925_
timestamp 1644511149
transform 1 0 17572 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2926_
timestamp 1644511149
transform 1 0 17940 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2927_
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2928_
timestamp 1644511149
transform 1 0 21068 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2929_
timestamp 1644511149
transform 1 0 19320 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2930_
timestamp 1644511149
transform 1 0 22448 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2931_
timestamp 1644511149
transform 1 0 21896 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2932_
timestamp 1644511149
transform 1 0 19780 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2933_
timestamp 1644511149
transform 1 0 20700 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2934_
timestamp 1644511149
transform 1 0 19780 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2935_
timestamp 1644511149
transform 1 0 18860 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2936_
timestamp 1644511149
transform 1 0 17848 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2937_
timestamp 1644511149
transform 1 0 19320 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2938_
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2939_
timestamp 1644511149
transform 1 0 16652 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2940_
timestamp 1644511149
transform 1 0 13984 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2941_
timestamp 1644511149
transform 1 0 14720 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2942_
timestamp 1644511149
transform 1 0 13708 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2943_
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2944_
timestamp 1644511149
transform 1 0 14720 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2945_
timestamp 1644511149
transform 1 0 13524 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2946_
timestamp 1644511149
transform 1 0 14536 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2947_
timestamp 1644511149
transform 1 0 14352 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2948_
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2949_
timestamp 1644511149
transform 1 0 11776 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2950_
timestamp 1644511149
transform 1 0 9476 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2951_
timestamp 1644511149
transform 1 0 17020 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _2952_
timestamp 1644511149
transform 1 0 30452 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2953_
timestamp 1644511149
transform 1 0 3036 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2954_
timestamp 1644511149
transform 1 0 31096 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2955_
timestamp 1644511149
transform 1 0 26220 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2956_
timestamp 1644511149
transform 1 0 28704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2957_
timestamp 1644511149
transform 1 0 29532 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2958_
timestamp 1644511149
transform 1 0 3864 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2959_
timestamp 1644511149
transform 1 0 31096 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2960_
timestamp 1644511149
transform 1 0 29532 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2961_
timestamp 1644511149
transform 1 0 31096 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20424 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk
timestamp 1644511149
transform 1 0 16376 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_prog_clk
timestamp 1644511149
transform 1 0 15456 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1644511149
transform 1 0 20792 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_prog_clk
timestamp 1644511149
transform 1 0 13248 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1644511149
transform 1 0 18216 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_prog_clk
timestamp 1644511149
transform 1 0 13156 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_prog_clk
timestamp 1644511149
transform 1 0 25852 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_prog_clk
timestamp 1644511149
transform 1 0 11868 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_prog_clk
timestamp 1644511149
transform 1 0 20240 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_0_prog_clk
timestamp 1644511149
transform 1 0 9292 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_1_prog_clk
timestamp 1644511149
transform 1 0 11776 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_2_prog_clk
timestamp 1644511149
transform 1 0 7728 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_3_prog_clk
timestamp 1644511149
transform 1 0 2944 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_4_prog_clk
timestamp 1644511149
transform 1 0 3404 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_5_prog_clk
timestamp 1644511149
transform 1 0 5704 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_6_prog_clk
timestamp 1644511149
transform 1 0 10580 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_7_prog_clk
timestamp 1644511149
transform 1 0 14996 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_8_prog_clk
timestamp 1644511149
transform 1 0 13524 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_9_prog_clk
timestamp 1644511149
transform 1 0 18584 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_10_prog_clk
timestamp 1644511149
transform 1 0 19504 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_11_prog_clk
timestamp 1644511149
transform 1 0 20608 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_12_prog_clk
timestamp 1644511149
transform 1 0 24656 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_13_prog_clk
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_14_prog_clk
timestamp 1644511149
transform 1 0 28244 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_15_prog_clk
timestamp 1644511149
transform 1 0 27140 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_16_prog_clk
timestamp 1644511149
transform 1 0 22172 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_17_prog_clk
timestamp 1644511149
transform 1 0 20240 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_18_prog_clk
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_19_prog_clk
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_20_prog_clk
timestamp 1644511149
transform 1 0 28612 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_21_prog_clk
timestamp 1644511149
transform 1 0 26956 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_22_prog_clk
timestamp 1644511149
transform 1 0 21712 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_23_prog_clk
timestamp 1644511149
transform 1 0 18400 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_24_prog_clk
timestamp 1644511149
transform 1 0 20056 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_25_prog_clk
timestamp 1644511149
transform 1 0 14444 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_26_prog_clk
timestamp 1644511149
transform 1 0 14444 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_27_prog_clk
timestamp 1644511149
transform 1 0 11868 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_28_prog_clk
timestamp 1644511149
transform 1 0 6624 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_29_prog_clk
timestamp 1644511149
transform 1 0 3220 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_30_prog_clk
timestamp 1644511149
transform 1 0 2760 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1644511149
transform 1 0 1748 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1644511149
transform 1 0 1748 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input3
timestamp 1644511149
transform 1 0 1748 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1644511149
transform 1 0 5612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1644511149
transform 1 0 4508 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1644511149
transform 1 0 1564 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1644511149
transform 1 0 1748 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input10
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1644511149
transform 1 0 1472 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input12
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1644511149
transform 1 0 1380 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input14
timestamp 1644511149
transform 1 0 1656 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input15
timestamp 1644511149
transform 1 0 4140 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 1644511149
transform 1 0 2484 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1644511149
transform 1 0 3772 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input20
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1644511149
transform 1 0 1656 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input22
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1644511149
transform 1 0 1656 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input24
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1644511149
transform 1 0 8924 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1644511149
transform 1 0 19412 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform 1 0 8188 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1644511149
transform 1 0 21804 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output29
timestamp 1644511149
transform 1 0 28796 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output30
timestamp 1644511149
transform 1 0 25576 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output31
timestamp 1644511149
transform 1 0 30452 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output32
timestamp 1644511149
transform 1 0 27232 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output33
timestamp 1644511149
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output34
timestamp 1644511149
transform 1 0 6532 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output35
timestamp 1644511149
transform 1 0 2208 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output36
timestamp 1644511149
transform 1 0 5612 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output37
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output38
timestamp 1644511149
transform 1 0 30176 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output39
timestamp 1644511149
transform 1 0 7176 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output40
timestamp 1644511149
transform 1 0 21528 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output41
timestamp 1644511149
transform 1 0 5612 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output42
timestamp 1644511149
transform 1 0 22908 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output43
timestamp 1644511149
transform 1 0 22264 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output44
timestamp 1644511149
transform 1 0 3036 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output45
timestamp 1644511149
transform 1 0 2300 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output46
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output47
timestamp 1644511149
transform 1 0 10120 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output48
timestamp 1644511149
transform 1 0 5520 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output49
timestamp 1644511149
transform 1 0 5612 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output50
timestamp 1644511149
transform 1 0 21068 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output51
timestamp 1644511149
transform 1 0 20424 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output52
timestamp 1644511149
transform 1 0 9936 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output53
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output54
timestamp 1644511149
transform 1 0 15180 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  repeater1
timestamp 1644511149
transform 1 0 28336 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  repeater2
timestamp 1644511149
transform 1 0 14720 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  repeater3
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 406 592
<< labels >>
rlabel metal1 s 0 890 800 946 6 bi_u1y0n_L1[0]
port 0 nsew signal input
rlabel metal1 s 0 37134 800 37190 6 bi_u1y0n_L1[10]
port 1 nsew signal input
rlabel metal1 s 0 40738 800 40794 6 bi_u1y0n_L1[11]
port 2 nsew signal input
rlabel metal1 s 0 4494 800 4550 6 bi_u1y0n_L1[1]
port 3 nsew signal input
rlabel metal1 s 0 8098 800 8154 6 bi_u1y0n_L1[2]
port 4 nsew signal input
rlabel metal1 s 0 11770 800 11826 6 bi_u1y0n_L1[3]
port 5 nsew signal input
rlabel metal1 s 0 15374 800 15430 6 bi_u1y0n_L1[4]
port 6 nsew signal input
rlabel metal1 s 0 18978 800 19034 6 bi_u1y0n_L1[5]
port 7 nsew signal input
rlabel metal1 s 0 22650 800 22706 6 bi_u1y0n_L1[6]
port 8 nsew signal input
rlabel metal1 s 0 26254 800 26310 6 bi_u1y0n_L1[7]
port 9 nsew signal input
rlabel metal1 s 0 29858 800 29914 6 bi_u1y0n_L1[8]
port 10 nsew signal input
rlabel metal1 s 0 33530 800 33586 6 bi_u1y0n_L1[9]
port 11 nsew signal input
rlabel metal1 s 0 2658 800 2714 6 bi_u1y0s_L1[0]
port 12 nsew signal input
rlabel metal1 s 0 38970 800 39026 6 bi_u1y0s_L1[10]
port 13 nsew signal input
rlabel metal1 s 0 42574 800 42630 6 bi_u1y0s_L1[11]
port 14 nsew signal input
rlabel metal1 s 0 6330 800 6386 6 bi_u1y0s_L1[1]
port 15 nsew signal input
rlabel metal1 s 0 9934 800 9990 6 bi_u1y0s_L1[2]
port 16 nsew signal input
rlabel metal1 s 0 13538 800 13594 6 bi_u1y0s_L1[3]
port 17 nsew signal input
rlabel metal1 s 0 17210 800 17266 6 bi_u1y0s_L1[4]
port 18 nsew signal input
rlabel metal1 s 0 20814 800 20870 6 bi_u1y0s_L1[5]
port 19 nsew signal input
rlabel metal1 s 0 24418 800 24474 6 bi_u1y0s_L1[6]
port 20 nsew signal input
rlabel metal1 s 0 28090 800 28146 6 bi_u1y0s_L1[7]
port 21 nsew signal input
rlabel metal1 s 0 31694 800 31750 6 bi_u1y0s_L1[8]
port 22 nsew signal input
rlabel metal1 s 0 35298 800 35354 6 bi_u1y0s_L1[9]
port 23 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 clk
port 24 nsew signal input
rlabel metal1 s 32320 890 33120 946 6 cu_x0y0n_L1[0]
port 25 nsew signal tristate
rlabel metal1 s 32320 37134 33120 37190 6 cu_x0y0n_L1[10]
port 26 nsew signal tristate
rlabel metal1 s 32320 40738 33120 40794 6 cu_x0y0n_L1[11]
port 27 nsew signal tristate
rlabel metal1 s 32320 4494 33120 4550 6 cu_x0y0n_L1[1]
port 28 nsew signal tristate
rlabel metal1 s 32320 8098 33120 8154 6 cu_x0y0n_L1[2]
port 29 nsew signal tristate
rlabel metal1 s 32320 11770 33120 11826 6 cu_x0y0n_L1[3]
port 30 nsew signal tristate
rlabel metal1 s 32320 15374 33120 15430 6 cu_x0y0n_L1[4]
port 31 nsew signal tristate
rlabel metal1 s 32320 18978 33120 19034 6 cu_x0y0n_L1[5]
port 32 nsew signal tristate
rlabel metal1 s 32320 22650 33120 22706 6 cu_x0y0n_L1[6]
port 33 nsew signal tristate
rlabel metal1 s 32320 26254 33120 26310 6 cu_x0y0n_L1[7]
port 34 nsew signal tristate
rlabel metal1 s 32320 29858 33120 29914 6 cu_x0y0n_L1[8]
port 35 nsew signal tristate
rlabel metal1 s 32320 33530 33120 33586 6 cu_x0y0n_L1[9]
port 36 nsew signal tristate
rlabel metal1 s 32320 2658 33120 2714 6 cu_x0y0s_L1[0]
port 37 nsew signal tristate
rlabel metal1 s 32320 38970 33120 39026 6 cu_x0y0s_L1[10]
port 38 nsew signal tristate
rlabel metal1 s 32320 42574 33120 42630 6 cu_x0y0s_L1[11]
port 39 nsew signal tristate
rlabel metal1 s 32320 6330 33120 6386 6 cu_x0y0s_L1[1]
port 40 nsew signal tristate
rlabel metal1 s 32320 9934 33120 9990 6 cu_x0y0s_L1[2]
port 41 nsew signal tristate
rlabel metal1 s 32320 13538 33120 13594 6 cu_x0y0s_L1[3]
port 42 nsew signal tristate
rlabel metal1 s 32320 17210 33120 17266 6 cu_x0y0s_L1[4]
port 43 nsew signal tristate
rlabel metal1 s 32320 20814 33120 20870 6 cu_x0y0s_L1[5]
port 44 nsew signal tristate
rlabel metal1 s 32320 24418 33120 24474 6 cu_x0y0s_L1[6]
port 45 nsew signal tristate
rlabel metal1 s 32320 28090 33120 28146 6 cu_x0y0s_L1[7]
port 46 nsew signal tristate
rlabel metal1 s 32320 31694 33120 31750 6 cu_x0y0s_L1[8]
port 47 nsew signal tristate
rlabel metal1 s 32320 35298 33120 35354 6 cu_x0y0s_L1[9]
port 48 nsew signal tristate
rlabel metal2 s 30378 0 30434 800 6 prog_clk
port 49 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 prog_din
port 50 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 prog_done
port 51 nsew signal input
rlabel metal2 s 8298 42720 8354 43520 6 prog_dout
port 52 nsew signal tristate
rlabel metal2 s 13818 0 13874 800 6 prog_rst
port 53 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 prog_we
port 54 nsew signal input
rlabel metal2 s 24858 42720 24914 43520 6 prog_we_o
port 55 nsew signal tristate
rlabel metal2 s 2134 1040 2190 42480 6 vccd1
port 56 nsew power input
rlabel metal2 s 12438 1040 12494 42480 6 vccd1
port 56 nsew power input
rlabel metal2 s 22742 1040 22798 42480 6 vccd1
port 56 nsew power input
rlabel metal2 s 7286 1040 7342 42480 6 vssd1
port 57 nsew ground input
rlabel metal2 s 17590 1040 17646 42480 6 vssd1
port 57 nsew ground input
rlabel metal2 s 27894 1040 27950 42480 6 vssd1
port 57 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 33120 43520
<< end >>
