VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top
  CLASS BLOCK ;
  FOREIGN top ;
  ORIGIN 0.000 0.000 ;
  SIZE 2600.000 BY 3200.000 ;
  PIN ipin_x0y1_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END ipin_x0y1_0
  PIN ipin_x0y1_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END ipin_x0y1_1
  PIN ipin_x0y2_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END ipin_x0y2_0
  PIN ipin_x0y2_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.280 4.000 233.880 ;
    END
  END ipin_x0y2_1
  PIN ipin_x0y3_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.920 4.000 300.520 ;
    END
  END ipin_x0y3_0
  PIN ipin_x0y3_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 366.560 4.000 367.160 ;
    END
  END ipin_x0y3_1
  PIN ipin_x0y4_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.200 4.000 433.800 ;
    END
  END ipin_x0y4_0
  PIN ipin_x0y4_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.840 4.000 500.440 ;
    END
  END ipin_x0y4_1
  PIN ipin_x0y5_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 566.480 4.000 567.080 ;
    END
  END ipin_x0y5_0
  PIN ipin_x0y5_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 633.120 4.000 633.720 ;
    END
  END ipin_x0y5_1
  PIN ipin_x0y6_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 699.760 4.000 700.360 ;
    END
  END ipin_x0y6_0
  PIN ipin_x0y6_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 766.400 4.000 767.000 ;
    END
  END ipin_x0y6_1
  PIN ipin_x0y7_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.040 4.000 833.640 ;
    END
  END ipin_x0y7_0
  PIN ipin_x0y7_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 899.680 4.000 900.280 ;
    END
  END ipin_x0y7_1
  PIN ipin_x0y8_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 966.320 4.000 966.920 ;
    END
  END ipin_x0y8_0
  PIN ipin_x0y8_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1032.960 4.000 1033.560 ;
    END
  END ipin_x0y8_1
  PIN ipin_x1y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 3196.000 27.050 3200.000 ;
    END
  END ipin_x1y9_0
  PIN ipin_x1y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 3196.000 80.870 3200.000 ;
    END
  END ipin_x1y9_1
  PIN ipin_x2y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 3196.000 135.150 3200.000 ;
    END
  END ipin_x2y9_0
  PIN ipin_x2y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 3196.000 189.430 3200.000 ;
    END
  END ipin_x2y9_1
  PIN ipin_x3y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 3196.000 243.710 3200.000 ;
    END
  END ipin_x3y9_0
  PIN ipin_x3y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 3196.000 297.530 3200.000 ;
    END
  END ipin_x3y9_1
  PIN ipin_x4y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 3196.000 351.810 3200.000 ;
    END
  END ipin_x4y9_0
  PIN ipin_x4y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 3196.000 406.090 3200.000 ;
    END
  END ipin_x4y9_1
  PIN ipin_x5y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 3196.000 460.370 3200.000 ;
    END
  END ipin_x5y9_0
  PIN ipin_x5y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 3196.000 514.190 3200.000 ;
    END
  END ipin_x5y9_1
  PIN ipin_x6y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.190 3196.000 568.470 3200.000 ;
    END
  END ipin_x6y9_0
  PIN ipin_x6y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.470 3196.000 622.750 3200.000 ;
    END
  END ipin_x6y9_1
  PIN ipin_x7y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 3196.000 677.030 3200.000 ;
    END
  END ipin_x7y9_0
  PIN ipin_x7y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.570 3196.000 730.850 3200.000 ;
    END
  END ipin_x7y9_1
  PIN ipin_x8y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.850 3196.000 785.130 3200.000 ;
    END
  END ipin_x8y9_0
  PIN ipin_x8y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.130 3196.000 839.410 3200.000 ;
    END
  END ipin_x8y9_1
  PIN ipin_x9y1_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 33.360 2600.000 33.960 ;
    END
  END ipin_x9y1_0
  PIN ipin_x9y1_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 100.000 2600.000 100.600 ;
    END
  END ipin_x9y1_1
  PIN ipin_x9y2_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 166.640 2600.000 167.240 ;
    END
  END ipin_x9y2_0
  PIN ipin_x9y2_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 233.280 2600.000 233.880 ;
    END
  END ipin_x9y2_1
  PIN ipin_x9y3_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 299.920 2600.000 300.520 ;
    END
  END ipin_x9y3_0
  PIN ipin_x9y3_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 366.560 2600.000 367.160 ;
    END
  END ipin_x9y3_1
  PIN ipin_x9y4_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 433.200 2600.000 433.800 ;
    END
  END ipin_x9y4_0
  PIN ipin_x9y4_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 499.840 2600.000 500.440 ;
    END
  END ipin_x9y4_1
  PIN ipin_x9y5_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 566.480 2600.000 567.080 ;
    END
  END ipin_x9y5_0
  PIN ipin_x9y5_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 633.120 2600.000 633.720 ;
    END
  END ipin_x9y5_1
  PIN ipin_x9y6_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 699.760 2600.000 700.360 ;
    END
  END ipin_x9y6_0
  PIN ipin_x9y6_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 766.400 2600.000 767.000 ;
    END
  END ipin_x9y6_1
  PIN ipin_x9y7_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 833.040 2600.000 833.640 ;
    END
  END ipin_x9y7_0
  PIN ipin_x9y7_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 899.680 2600.000 900.280 ;
    END
  END ipin_x9y7_1
  PIN ipin_x9y8_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 966.320 2600.000 966.920 ;
    END
  END ipin_x9y8_0
  PIN ipin_x9y8_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1032.960 2600.000 1033.560 ;
    END
  END ipin_x9y8_1
  PIN oe_x0y1_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2166.520 4.000 2167.120 ;
    END
  END oe_x0y1_0
  PIN oe_x0y1_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2233.160 4.000 2233.760 ;
    END
  END oe_x0y1_1
  PIN oe_x0y2_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2299.800 4.000 2300.400 ;
    END
  END oe_x0y2_0
  PIN oe_x0y2_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2366.440 4.000 2367.040 ;
    END
  END oe_x0y2_1
  PIN oe_x0y3_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2433.080 4.000 2433.680 ;
    END
  END oe_x0y3_0
  PIN oe_x0y3_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2499.720 4.000 2500.320 ;
    END
  END oe_x0y3_1
  PIN oe_x0y4_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2566.360 4.000 2566.960 ;
    END
  END oe_x0y4_0
  PIN oe_x0y4_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2633.000 4.000 2633.600 ;
    END
  END oe_x0y4_1
  PIN oe_x0y5_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2699.640 4.000 2700.240 ;
    END
  END oe_x0y5_0
  PIN oe_x0y5_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2766.280 4.000 2766.880 ;
    END
  END oe_x0y5_1
  PIN oe_x0y6_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2832.920 4.000 2833.520 ;
    END
  END oe_x0y6_0
  PIN oe_x0y6_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2899.560 4.000 2900.160 ;
    END
  END oe_x0y6_1
  PIN oe_x0y7_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2966.200 4.000 2966.800 ;
    END
  END oe_x0y7_0
  PIN oe_x0y7_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3032.840 4.000 3033.440 ;
    END
  END oe_x0y7_1
  PIN oe_x0y8_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3099.480 4.000 3100.080 ;
    END
  END oe_x0y8_0
  PIN oe_x0y8_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3166.120 4.000 3166.720 ;
    END
  END oe_x0y8_1
  PIN oe_x1y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.050 3196.000 1760.330 3200.000 ;
    END
  END oe_x1y9_0
  PIN oe_x1y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1813.870 3196.000 1814.150 3200.000 ;
    END
  END oe_x1y9_1
  PIN oe_x2y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1868.150 3196.000 1868.430 3200.000 ;
    END
  END oe_x2y9_0
  PIN oe_x2y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1922.430 3196.000 1922.710 3200.000 ;
    END
  END oe_x2y9_1
  PIN oe_x3y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.710 3196.000 1976.990 3200.000 ;
    END
  END oe_x3y9_0
  PIN oe_x3y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.530 3196.000 2030.810 3200.000 ;
    END
  END oe_x3y9_1
  PIN oe_x4y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2084.810 3196.000 2085.090 3200.000 ;
    END
  END oe_x4y9_0
  PIN oe_x4y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2139.090 3196.000 2139.370 3200.000 ;
    END
  END oe_x4y9_1
  PIN oe_x5y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2193.370 3196.000 2193.650 3200.000 ;
    END
  END oe_x5y9_0
  PIN oe_x5y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2247.190 3196.000 2247.470 3200.000 ;
    END
  END oe_x5y9_1
  PIN oe_x6y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.470 3196.000 2301.750 3200.000 ;
    END
  END oe_x6y9_0
  PIN oe_x6y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2355.750 3196.000 2356.030 3200.000 ;
    END
  END oe_x6y9_1
  PIN oe_x7y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2410.030 3196.000 2410.310 3200.000 ;
    END
  END oe_x7y9_0
  PIN oe_x7y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2463.850 3196.000 2464.130 3200.000 ;
    END
  END oe_x7y9_1
  PIN oe_x8y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2518.130 3196.000 2518.410 3200.000 ;
    END
  END oe_x8y9_0
  PIN oe_x8y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2572.410 3196.000 2572.690 3200.000 ;
    END
  END oe_x8y9_1
  PIN oe_x9y1_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2166.520 2600.000 2167.120 ;
    END
  END oe_x9y1_0
  PIN oe_x9y1_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2233.160 2600.000 2233.760 ;
    END
  END oe_x9y1_1
  PIN oe_x9y2_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2299.800 2600.000 2300.400 ;
    END
  END oe_x9y2_0
  PIN oe_x9y2_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2366.440 2600.000 2367.040 ;
    END
  END oe_x9y2_1
  PIN oe_x9y3_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2433.080 2600.000 2433.680 ;
    END
  END oe_x9y3_0
  PIN oe_x9y3_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2499.720 2600.000 2500.320 ;
    END
  END oe_x9y3_1
  PIN oe_x9y4_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2566.360 2600.000 2566.960 ;
    END
  END oe_x9y4_0
  PIN oe_x9y4_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2633.000 2600.000 2633.600 ;
    END
  END oe_x9y4_1
  PIN oe_x9y5_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2699.640 2600.000 2700.240 ;
    END
  END oe_x9y5_0
  PIN oe_x9y5_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2766.280 2600.000 2766.880 ;
    END
  END oe_x9y5_1
  PIN oe_x9y6_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2832.920 2600.000 2833.520 ;
    END
  END oe_x9y6_0
  PIN oe_x9y6_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2899.560 2600.000 2900.160 ;
    END
  END oe_x9y6_1
  PIN oe_x9y7_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2966.200 2600.000 2966.800 ;
    END
  END oe_x9y7_0
  PIN oe_x9y7_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 3032.840 2600.000 3033.440 ;
    END
  END oe_x9y7_1
  PIN oe_x9y8_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 3099.480 2600.000 3100.080 ;
    END
  END oe_x9y8_0
  PIN oe_x9y8_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 3166.120 2600.000 3166.720 ;
    END
  END oe_x9y8_1
  PIN opin_x0y1_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1099.600 4.000 1100.200 ;
    END
  END opin_x0y1_0
  PIN opin_x0y1_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1166.240 4.000 1166.840 ;
    END
  END opin_x0y1_1
  PIN opin_x0y2_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1232.880 4.000 1233.480 ;
    END
  END opin_x0y2_0
  PIN opin_x0y2_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1299.520 4.000 1300.120 ;
    END
  END opin_x0y2_1
  PIN opin_x0y3_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1366.160 4.000 1366.760 ;
    END
  END opin_x0y3_0
  PIN opin_x0y3_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1432.800 4.000 1433.400 ;
    END
  END opin_x0y3_1
  PIN opin_x0y4_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1499.440 4.000 1500.040 ;
    END
  END opin_x0y4_0
  PIN opin_x0y4_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1566.080 4.000 1566.680 ;
    END
  END opin_x0y4_1
  PIN opin_x0y5_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1633.400 4.000 1634.000 ;
    END
  END opin_x0y5_0
  PIN opin_x0y5_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1700.040 4.000 1700.640 ;
    END
  END opin_x0y5_1
  PIN opin_x0y6_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1766.680 4.000 1767.280 ;
    END
  END opin_x0y6_0
  PIN opin_x0y6_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1833.320 4.000 1833.920 ;
    END
  END opin_x0y6_1
  PIN opin_x0y7_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1899.960 4.000 1900.560 ;
    END
  END opin_x0y7_0
  PIN opin_x0y7_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1966.600 4.000 1967.200 ;
    END
  END opin_x0y7_1
  PIN opin_x0y8_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2033.240 4.000 2033.840 ;
    END
  END opin_x0y8_0
  PIN opin_x0y8_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2099.880 4.000 2100.480 ;
    END
  END opin_x0y8_1
  PIN opin_x1y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.410 3196.000 893.690 3200.000 ;
    END
  END opin_x1y9_0
  PIN opin_x1y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.230 3196.000 947.510 3200.000 ;
    END
  END opin_x1y9_1
  PIN opin_x2y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.510 3196.000 1001.790 3200.000 ;
    END
  END opin_x2y9_0
  PIN opin_x2y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1055.790 3196.000 1056.070 3200.000 ;
    END
  END opin_x2y9_1
  PIN opin_x3y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.070 3196.000 1110.350 3200.000 ;
    END
  END opin_x3y9_0
  PIN opin_x3y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1163.890 3196.000 1164.170 3200.000 ;
    END
  END opin_x3y9_1
  PIN opin_x4y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1218.170 3196.000 1218.450 3200.000 ;
    END
  END opin_x4y9_0
  PIN opin_x4y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1272.450 3196.000 1272.730 3200.000 ;
    END
  END opin_x4y9_1
  PIN opin_x5y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.730 3196.000 1327.010 3200.000 ;
    END
  END opin_x5y9_0
  PIN opin_x5y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1380.550 3196.000 1380.830 3200.000 ;
    END
  END opin_x5y9_1
  PIN opin_x6y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1434.830 3196.000 1435.110 3200.000 ;
    END
  END opin_x6y9_0
  PIN opin_x6y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.110 3196.000 1489.390 3200.000 ;
    END
  END opin_x6y9_1
  PIN opin_x7y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1543.390 3196.000 1543.670 3200.000 ;
    END
  END opin_x7y9_0
  PIN opin_x7y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.210 3196.000 1597.490 3200.000 ;
    END
  END opin_x7y9_1
  PIN opin_x8y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.490 3196.000 1651.770 3200.000 ;
    END
  END opin_x8y9_0
  PIN opin_x8y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1705.770 3196.000 1706.050 3200.000 ;
    END
  END opin_x8y9_1
  PIN opin_x9y1_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1099.600 2600.000 1100.200 ;
    END
  END opin_x9y1_0
  PIN opin_x9y1_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1166.240 2600.000 1166.840 ;
    END
  END opin_x9y1_1
  PIN opin_x9y2_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1232.880 2600.000 1233.480 ;
    END
  END opin_x9y2_0
  PIN opin_x9y2_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1299.520 2600.000 1300.120 ;
    END
  END opin_x9y2_1
  PIN opin_x9y3_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1366.160 2600.000 1366.760 ;
    END
  END opin_x9y3_0
  PIN opin_x9y3_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1432.800 2600.000 1433.400 ;
    END
  END opin_x9y3_1
  PIN opin_x9y4_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1499.440 2600.000 1500.040 ;
    END
  END opin_x9y4_0
  PIN opin_x9y4_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1566.080 2600.000 1566.680 ;
    END
  END opin_x9y4_1
  PIN opin_x9y5_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1633.400 2600.000 1634.000 ;
    END
  END opin_x9y5_0
  PIN opin_x9y5_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1700.040 2600.000 1700.640 ;
    END
  END opin_x9y5_1
  PIN opin_x9y6_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1766.680 2600.000 1767.280 ;
    END
  END opin_x9y6_0
  PIN opin_x9y6_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1833.320 2600.000 1833.920 ;
    END
  END opin_x9y6_1
  PIN opin_x9y7_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1899.960 2600.000 1900.560 ;
    END
  END opin_x9y7_0
  PIN opin_x9y7_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1966.600 2600.000 1967.200 ;
    END
  END opin_x9y7_1
  PIN opin_x9y8_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2033.240 2600.000 2033.840 ;
    END
  END opin_x9y8_0
  PIN opin_x9y8_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2099.880 2600.000 2100.480 ;
    END
  END opin_x9y8_1
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END prog_clk
  PIN prog_din
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 0.000 556.970 4.000 ;
    END
  END prog_din
  PIN prog_done
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.910 0.000 928.190 4.000 ;
    END
  END prog_done
  PIN prog_dout
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1299.590 0.000 1299.870 4.000 ;
    END
  END prog_dout
  PIN prog_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1670.810 0.000 1671.090 4.000 ;
    END
  END prog_rst
  PIN prog_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2042.490 0.000 2042.770 4.000 ;
    END
  END prog_we
  PIN prog_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2413.710 0.000 2413.990 4.000 ;
    END
  END prog_we_o
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 3188.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2555.440 10.640 2557.040 3188.080 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2594.400 3187.925 ;
      LAYER met1 ;
        RECT 5.520 10.640 2597.090 3188.080 ;
      LAYER met2 ;
        RECT 6.990 3195.720 26.490 3196.410 ;
        RECT 27.330 3195.720 80.310 3196.410 ;
        RECT 81.150 3195.720 134.590 3196.410 ;
        RECT 135.430 3195.720 188.870 3196.410 ;
        RECT 189.710 3195.720 243.150 3196.410 ;
        RECT 243.990 3195.720 296.970 3196.410 ;
        RECT 297.810 3195.720 351.250 3196.410 ;
        RECT 352.090 3195.720 405.530 3196.410 ;
        RECT 406.370 3195.720 459.810 3196.410 ;
        RECT 460.650 3195.720 513.630 3196.410 ;
        RECT 514.470 3195.720 567.910 3196.410 ;
        RECT 568.750 3195.720 622.190 3196.410 ;
        RECT 623.030 3195.720 676.470 3196.410 ;
        RECT 677.310 3195.720 730.290 3196.410 ;
        RECT 731.130 3195.720 784.570 3196.410 ;
        RECT 785.410 3195.720 838.850 3196.410 ;
        RECT 839.690 3195.720 893.130 3196.410 ;
        RECT 893.970 3195.720 946.950 3196.410 ;
        RECT 947.790 3195.720 1001.230 3196.410 ;
        RECT 1002.070 3195.720 1055.510 3196.410 ;
        RECT 1056.350 3195.720 1109.790 3196.410 ;
        RECT 1110.630 3195.720 1163.610 3196.410 ;
        RECT 1164.450 3195.720 1217.890 3196.410 ;
        RECT 1218.730 3195.720 1272.170 3196.410 ;
        RECT 1273.010 3195.720 1326.450 3196.410 ;
        RECT 1327.290 3195.720 1380.270 3196.410 ;
        RECT 1381.110 3195.720 1434.550 3196.410 ;
        RECT 1435.390 3195.720 1488.830 3196.410 ;
        RECT 1489.670 3195.720 1543.110 3196.410 ;
        RECT 1543.950 3195.720 1596.930 3196.410 ;
        RECT 1597.770 3195.720 1651.210 3196.410 ;
        RECT 1652.050 3195.720 1705.490 3196.410 ;
        RECT 1706.330 3195.720 1759.770 3196.410 ;
        RECT 1760.610 3195.720 1813.590 3196.410 ;
        RECT 1814.430 3195.720 1867.870 3196.410 ;
        RECT 1868.710 3195.720 1922.150 3196.410 ;
        RECT 1922.990 3195.720 1976.430 3196.410 ;
        RECT 1977.270 3195.720 2030.250 3196.410 ;
        RECT 2031.090 3195.720 2084.530 3196.410 ;
        RECT 2085.370 3195.720 2138.810 3196.410 ;
        RECT 2139.650 3195.720 2193.090 3196.410 ;
        RECT 2193.930 3195.720 2246.910 3196.410 ;
        RECT 2247.750 3195.720 2301.190 3196.410 ;
        RECT 2302.030 3195.720 2355.470 3196.410 ;
        RECT 2356.310 3195.720 2409.750 3196.410 ;
        RECT 2410.590 3195.720 2463.570 3196.410 ;
        RECT 2464.410 3195.720 2517.850 3196.410 ;
        RECT 2518.690 3195.720 2572.130 3196.410 ;
        RECT 2572.970 3195.720 2597.060 3196.410 ;
        RECT 6.990 4.280 2597.060 3195.720 ;
        RECT 6.990 3.670 185.190 4.280 ;
        RECT 186.030 3.670 556.410 4.280 ;
        RECT 557.250 3.670 927.630 4.280 ;
        RECT 928.470 3.670 1299.310 4.280 ;
        RECT 1300.150 3.670 1670.530 4.280 ;
        RECT 1671.370 3.670 2042.210 4.280 ;
        RECT 2043.050 3.670 2413.430 4.280 ;
        RECT 2414.270 3.670 2597.060 4.280 ;
      LAYER met3 ;
        RECT 4.000 3167.120 2596.000 3188.005 ;
        RECT 4.400 3165.720 2595.600 3167.120 ;
        RECT 4.000 3100.480 2596.000 3165.720 ;
        RECT 4.400 3099.080 2595.600 3100.480 ;
        RECT 4.000 3033.840 2596.000 3099.080 ;
        RECT 4.400 3032.440 2595.600 3033.840 ;
        RECT 4.000 2967.200 2596.000 3032.440 ;
        RECT 4.400 2965.800 2595.600 2967.200 ;
        RECT 4.000 2900.560 2596.000 2965.800 ;
        RECT 4.400 2899.160 2595.600 2900.560 ;
        RECT 4.000 2833.920 2596.000 2899.160 ;
        RECT 4.400 2832.520 2595.600 2833.920 ;
        RECT 4.000 2767.280 2596.000 2832.520 ;
        RECT 4.400 2765.880 2595.600 2767.280 ;
        RECT 4.000 2700.640 2596.000 2765.880 ;
        RECT 4.400 2699.240 2595.600 2700.640 ;
        RECT 4.000 2634.000 2596.000 2699.240 ;
        RECT 4.400 2632.600 2595.600 2634.000 ;
        RECT 4.000 2567.360 2596.000 2632.600 ;
        RECT 4.400 2565.960 2595.600 2567.360 ;
        RECT 4.000 2500.720 2596.000 2565.960 ;
        RECT 4.400 2499.320 2595.600 2500.720 ;
        RECT 4.000 2434.080 2596.000 2499.320 ;
        RECT 4.400 2432.680 2595.600 2434.080 ;
        RECT 4.000 2367.440 2596.000 2432.680 ;
        RECT 4.400 2366.040 2595.600 2367.440 ;
        RECT 4.000 2300.800 2596.000 2366.040 ;
        RECT 4.400 2299.400 2595.600 2300.800 ;
        RECT 4.000 2234.160 2596.000 2299.400 ;
        RECT 4.400 2232.760 2595.600 2234.160 ;
        RECT 4.000 2167.520 2596.000 2232.760 ;
        RECT 4.400 2166.120 2595.600 2167.520 ;
        RECT 4.000 2100.880 2596.000 2166.120 ;
        RECT 4.400 2099.480 2595.600 2100.880 ;
        RECT 4.000 2034.240 2596.000 2099.480 ;
        RECT 4.400 2032.840 2595.600 2034.240 ;
        RECT 4.000 1967.600 2596.000 2032.840 ;
        RECT 4.400 1966.200 2595.600 1967.600 ;
        RECT 4.000 1900.960 2596.000 1966.200 ;
        RECT 4.400 1899.560 2595.600 1900.960 ;
        RECT 4.000 1834.320 2596.000 1899.560 ;
        RECT 4.400 1832.920 2595.600 1834.320 ;
        RECT 4.000 1767.680 2596.000 1832.920 ;
        RECT 4.400 1766.280 2595.600 1767.680 ;
        RECT 4.000 1701.040 2596.000 1766.280 ;
        RECT 4.400 1699.640 2595.600 1701.040 ;
        RECT 4.000 1634.400 2596.000 1699.640 ;
        RECT 4.400 1633.000 2595.600 1634.400 ;
        RECT 4.000 1567.080 2596.000 1633.000 ;
        RECT 4.400 1565.680 2595.600 1567.080 ;
        RECT 4.000 1500.440 2596.000 1565.680 ;
        RECT 4.400 1499.040 2595.600 1500.440 ;
        RECT 4.000 1433.800 2596.000 1499.040 ;
        RECT 4.400 1432.400 2595.600 1433.800 ;
        RECT 4.000 1367.160 2596.000 1432.400 ;
        RECT 4.400 1365.760 2595.600 1367.160 ;
        RECT 4.000 1300.520 2596.000 1365.760 ;
        RECT 4.400 1299.120 2595.600 1300.520 ;
        RECT 4.000 1233.880 2596.000 1299.120 ;
        RECT 4.400 1232.480 2595.600 1233.880 ;
        RECT 4.000 1167.240 2596.000 1232.480 ;
        RECT 4.400 1165.840 2595.600 1167.240 ;
        RECT 4.000 1100.600 2596.000 1165.840 ;
        RECT 4.400 1099.200 2595.600 1100.600 ;
        RECT 4.000 1033.960 2596.000 1099.200 ;
        RECT 4.400 1032.560 2595.600 1033.960 ;
        RECT 4.000 967.320 2596.000 1032.560 ;
        RECT 4.400 965.920 2595.600 967.320 ;
        RECT 4.000 900.680 2596.000 965.920 ;
        RECT 4.400 899.280 2595.600 900.680 ;
        RECT 4.000 834.040 2596.000 899.280 ;
        RECT 4.400 832.640 2595.600 834.040 ;
        RECT 4.000 767.400 2596.000 832.640 ;
        RECT 4.400 766.000 2595.600 767.400 ;
        RECT 4.000 700.760 2596.000 766.000 ;
        RECT 4.400 699.360 2595.600 700.760 ;
        RECT 4.000 634.120 2596.000 699.360 ;
        RECT 4.400 632.720 2595.600 634.120 ;
        RECT 4.000 567.480 2596.000 632.720 ;
        RECT 4.400 566.080 2595.600 567.480 ;
        RECT 4.000 500.840 2596.000 566.080 ;
        RECT 4.400 499.440 2595.600 500.840 ;
        RECT 4.000 434.200 2596.000 499.440 ;
        RECT 4.400 432.800 2595.600 434.200 ;
        RECT 4.000 367.560 2596.000 432.800 ;
        RECT 4.400 366.160 2595.600 367.560 ;
        RECT 4.000 300.920 2596.000 366.160 ;
        RECT 4.400 299.520 2595.600 300.920 ;
        RECT 4.000 234.280 2596.000 299.520 ;
        RECT 4.400 232.880 2595.600 234.280 ;
        RECT 4.000 167.640 2596.000 232.880 ;
        RECT 4.400 166.240 2595.600 167.640 ;
        RECT 4.000 101.000 2596.000 166.240 ;
        RECT 4.400 99.600 2595.600 101.000 ;
        RECT 4.000 34.360 2596.000 99.600 ;
        RECT 4.400 32.960 2595.600 34.360 ;
        RECT 4.000 10.715 2596.000 32.960 ;
      LAYER met4 ;
        RECT 40.775 102.175 97.440 3128.505 ;
        RECT 99.840 102.175 174.240 3128.505 ;
        RECT 176.640 102.175 251.040 3128.505 ;
        RECT 253.440 102.175 327.840 3128.505 ;
        RECT 330.240 102.175 404.640 3128.505 ;
        RECT 407.040 102.175 481.440 3128.505 ;
        RECT 483.840 102.175 558.240 3128.505 ;
        RECT 560.640 102.175 635.040 3128.505 ;
        RECT 637.440 102.175 711.840 3128.505 ;
        RECT 714.240 102.175 788.640 3128.505 ;
        RECT 791.040 102.175 865.440 3128.505 ;
        RECT 867.840 102.175 942.240 3128.505 ;
        RECT 944.640 102.175 1019.040 3128.505 ;
        RECT 1021.440 102.175 1095.840 3128.505 ;
        RECT 1098.240 102.175 1172.640 3128.505 ;
        RECT 1175.040 102.175 1249.440 3128.505 ;
        RECT 1251.840 102.175 1326.240 3128.505 ;
        RECT 1328.640 102.175 1403.040 3128.505 ;
        RECT 1405.440 102.175 1479.840 3128.505 ;
        RECT 1482.240 102.175 1556.640 3128.505 ;
        RECT 1559.040 102.175 1633.440 3128.505 ;
        RECT 1635.840 102.175 1710.240 3128.505 ;
        RECT 1712.640 102.175 1787.040 3128.505 ;
        RECT 1789.440 102.175 1863.840 3128.505 ;
        RECT 1866.240 102.175 1940.640 3128.505 ;
        RECT 1943.040 102.175 2017.440 3128.505 ;
        RECT 2019.840 102.175 2094.240 3128.505 ;
        RECT 2096.640 102.175 2171.040 3128.505 ;
        RECT 2173.440 102.175 2247.840 3128.505 ;
        RECT 2250.240 102.175 2324.640 3128.505 ;
        RECT 2327.040 102.175 2401.440 3128.505 ;
        RECT 2403.840 102.175 2478.240 3128.505 ;
        RECT 2480.640 102.175 2481.865 3128.505 ;
  END
END top
END LIBRARY

