magic
tech sky130A
magscale 1 2
timestamp 1653678508
<< obsli1 >>
rect 1104 2159 518880 637585
<< obsm1 >>
rect 1104 2128 519970 637616
<< metal2 >>
rect 4802 639200 4858 640000
rect 14370 639200 14426 640000
rect 24030 639200 24086 640000
rect 33690 639200 33746 640000
rect 43258 639200 43314 640000
rect 52918 639200 52974 640000
rect 62578 639200 62634 640000
rect 72146 639200 72202 640000
rect 81806 639200 81862 640000
rect 91466 639200 91522 640000
rect 101034 639200 101090 640000
rect 110694 639200 110750 640000
rect 120354 639200 120410 640000
rect 129922 639200 129978 640000
rect 139582 639200 139638 640000
rect 149242 639200 149298 640000
rect 158810 639200 158866 640000
rect 168470 639200 168526 640000
rect 178130 639200 178186 640000
rect 187698 639200 187754 640000
rect 197358 639200 197414 640000
rect 207018 639200 207074 640000
rect 216586 639200 216642 640000
rect 226246 639200 226302 640000
rect 235906 639200 235962 640000
rect 245474 639200 245530 640000
rect 255134 639200 255190 640000
rect 264794 639200 264850 640000
rect 274362 639200 274418 640000
rect 284022 639200 284078 640000
rect 293682 639200 293738 640000
rect 303250 639200 303306 640000
rect 312910 639200 312966 640000
rect 322570 639200 322626 640000
rect 332138 639200 332194 640000
rect 341798 639200 341854 640000
rect 351458 639200 351514 640000
rect 361026 639200 361082 640000
rect 370686 639200 370742 640000
rect 380346 639200 380402 640000
rect 389914 639200 389970 640000
rect 399574 639200 399630 640000
rect 409234 639200 409290 640000
rect 418802 639200 418858 640000
rect 428462 639200 428518 640000
rect 438122 639200 438178 640000
rect 447690 639200 447746 640000
rect 457350 639200 457406 640000
rect 467010 639200 467066 640000
rect 476578 639200 476634 640000
rect 486238 639200 486294 640000
rect 495898 639200 495954 640000
rect 505466 639200 505522 640000
rect 515126 639200 515182 640000
rect 37094 0 37150 800
rect 111338 0 111394 800
rect 185582 0 185638 800
rect 259918 0 259974 800
rect 334162 0 334218 800
rect 408498 0 408554 800
rect 482742 0 482798 800
<< obsm2 >>
rect 1216 639144 4746 639282
rect 4914 639144 14314 639282
rect 14482 639144 23974 639282
rect 24142 639144 33634 639282
rect 33802 639144 43202 639282
rect 43370 639144 52862 639282
rect 53030 639144 62522 639282
rect 62690 639144 72090 639282
rect 72258 639144 81750 639282
rect 81918 639144 91410 639282
rect 91578 639144 100978 639282
rect 101146 639144 110638 639282
rect 110806 639144 120298 639282
rect 120466 639144 129866 639282
rect 130034 639144 139526 639282
rect 139694 639144 149186 639282
rect 149354 639144 158754 639282
rect 158922 639144 168414 639282
rect 168582 639144 178074 639282
rect 178242 639144 187642 639282
rect 187810 639144 197302 639282
rect 197470 639144 206962 639282
rect 207130 639144 216530 639282
rect 216698 639144 226190 639282
rect 226358 639144 235850 639282
rect 236018 639144 245418 639282
rect 245586 639144 255078 639282
rect 255246 639144 264738 639282
rect 264906 639144 274306 639282
rect 274474 639144 283966 639282
rect 284134 639144 293626 639282
rect 293794 639144 303194 639282
rect 303362 639144 312854 639282
rect 313022 639144 322514 639282
rect 322682 639144 332082 639282
rect 332250 639144 341742 639282
rect 341910 639144 351402 639282
rect 351570 639144 360970 639282
rect 361138 639144 370630 639282
rect 370798 639144 380290 639282
rect 380458 639144 389858 639282
rect 390026 639144 399518 639282
rect 399686 639144 409178 639282
rect 409346 639144 418746 639282
rect 418914 639144 428406 639282
rect 428574 639144 438066 639282
rect 438234 639144 447634 639282
rect 447802 639144 457294 639282
rect 457462 639144 466954 639282
rect 467122 639144 476522 639282
rect 476690 639144 486182 639282
rect 486350 639144 495842 639282
rect 496010 639144 505410 639282
rect 505578 639144 515070 639282
rect 515238 639144 519964 639282
rect 1216 856 519964 639144
rect 1216 800 37038 856
rect 37206 800 111282 856
rect 111450 800 185526 856
rect 185694 800 259862 856
rect 260030 800 334106 856
rect 334274 800 408442 856
rect 408610 800 482686 856
rect 482854 800 519964 856
<< metal3 >>
rect 0 633904 800 634024
rect 519200 633904 520000 634024
rect 0 622072 800 622192
rect 519200 622072 520000 622192
rect 0 610240 800 610360
rect 519200 610240 520000 610360
rect 0 598408 800 598528
rect 519200 598408 520000 598528
rect 0 586576 800 586696
rect 519200 586576 520000 586696
rect 0 574744 800 574864
rect 519200 574744 520000 574864
rect 0 562776 800 562896
rect 519200 562776 520000 562896
rect 0 550944 800 551064
rect 519200 550944 520000 551064
rect 0 539112 800 539232
rect 519200 539112 520000 539232
rect 0 527280 800 527400
rect 519200 527280 520000 527400
rect 0 515448 800 515568
rect 519200 515448 520000 515568
rect 0 503616 800 503736
rect 519200 503616 520000 503736
rect 0 491784 800 491904
rect 519200 491784 520000 491904
rect 0 479816 800 479936
rect 519200 479816 520000 479936
rect 0 467984 800 468104
rect 519200 467984 520000 468104
rect 0 456152 800 456272
rect 519200 456152 520000 456272
rect 0 444320 800 444440
rect 519200 444320 520000 444440
rect 0 432488 800 432608
rect 519200 432488 520000 432608
rect 0 420656 800 420776
rect 519200 420656 520000 420776
rect 0 408824 800 408944
rect 519200 408824 520000 408944
rect 0 396856 800 396976
rect 519200 396856 520000 396976
rect 0 385024 800 385144
rect 519200 385024 520000 385144
rect 0 373192 800 373312
rect 519200 373192 520000 373312
rect 0 361360 800 361480
rect 519200 361360 520000 361480
rect 0 349528 800 349648
rect 519200 349528 520000 349648
rect 0 337696 800 337816
rect 519200 337696 520000 337816
rect 0 325864 800 325984
rect 519200 325864 520000 325984
rect 0 313896 800 314016
rect 519200 313896 520000 314016
rect 0 302064 800 302184
rect 519200 302064 520000 302184
rect 0 290232 800 290352
rect 519200 290232 520000 290352
rect 0 278400 800 278520
rect 519200 278400 520000 278520
rect 0 266568 800 266688
rect 519200 266568 520000 266688
rect 0 254736 800 254856
rect 519200 254736 520000 254856
rect 0 242768 800 242888
rect 519200 242768 520000 242888
rect 0 230936 800 231056
rect 519200 230936 520000 231056
rect 0 219104 800 219224
rect 519200 219104 520000 219224
rect 0 207272 800 207392
rect 519200 207272 520000 207392
rect 0 195440 800 195560
rect 519200 195440 520000 195560
rect 0 183608 800 183728
rect 519200 183608 520000 183728
rect 0 171776 800 171896
rect 519200 171776 520000 171896
rect 0 159808 800 159928
rect 519200 159808 520000 159928
rect 0 147976 800 148096
rect 519200 147976 520000 148096
rect 0 136144 800 136264
rect 519200 136144 520000 136264
rect 0 124312 800 124432
rect 519200 124312 520000 124432
rect 0 112480 800 112600
rect 519200 112480 520000 112600
rect 0 100648 800 100768
rect 519200 100648 520000 100768
rect 0 88816 800 88936
rect 519200 88816 520000 88936
rect 0 76848 800 76968
rect 519200 76848 520000 76968
rect 0 65016 800 65136
rect 519200 65016 520000 65136
rect 0 53184 800 53304
rect 519200 53184 520000 53304
rect 0 41352 800 41472
rect 519200 41352 520000 41472
rect 0 29520 800 29640
rect 519200 29520 520000 29640
rect 0 17688 800 17808
rect 519200 17688 520000 17808
rect 0 5856 800 5976
rect 519200 5856 520000 5976
<< obsm3 >>
rect 800 634104 519200 637601
rect 880 633824 519120 634104
rect 800 622272 519200 633824
rect 880 621992 519120 622272
rect 800 610440 519200 621992
rect 880 610160 519120 610440
rect 800 598608 519200 610160
rect 880 598328 519120 598608
rect 800 586776 519200 598328
rect 880 586496 519120 586776
rect 800 574944 519200 586496
rect 880 574664 519120 574944
rect 800 562976 519200 574664
rect 880 562696 519120 562976
rect 800 551144 519200 562696
rect 880 550864 519120 551144
rect 800 539312 519200 550864
rect 880 539032 519120 539312
rect 800 527480 519200 539032
rect 880 527200 519120 527480
rect 800 515648 519200 527200
rect 880 515368 519120 515648
rect 800 503816 519200 515368
rect 880 503536 519120 503816
rect 800 491984 519200 503536
rect 880 491704 519120 491984
rect 800 480016 519200 491704
rect 880 479736 519120 480016
rect 800 468184 519200 479736
rect 880 467904 519120 468184
rect 800 456352 519200 467904
rect 880 456072 519120 456352
rect 800 444520 519200 456072
rect 880 444240 519120 444520
rect 800 432688 519200 444240
rect 880 432408 519120 432688
rect 800 420856 519200 432408
rect 880 420576 519120 420856
rect 800 409024 519200 420576
rect 880 408744 519120 409024
rect 800 397056 519200 408744
rect 880 396776 519120 397056
rect 800 385224 519200 396776
rect 880 384944 519120 385224
rect 800 373392 519200 384944
rect 880 373112 519120 373392
rect 800 361560 519200 373112
rect 880 361280 519120 361560
rect 800 349728 519200 361280
rect 880 349448 519120 349728
rect 800 337896 519200 349448
rect 880 337616 519120 337896
rect 800 326064 519200 337616
rect 880 325784 519120 326064
rect 800 314096 519200 325784
rect 880 313816 519120 314096
rect 800 302264 519200 313816
rect 880 301984 519120 302264
rect 800 290432 519200 301984
rect 880 290152 519120 290432
rect 800 278600 519200 290152
rect 880 278320 519120 278600
rect 800 266768 519200 278320
rect 880 266488 519120 266768
rect 800 254936 519200 266488
rect 880 254656 519120 254936
rect 800 242968 519200 254656
rect 880 242688 519120 242968
rect 800 231136 519200 242688
rect 880 230856 519120 231136
rect 800 219304 519200 230856
rect 880 219024 519120 219304
rect 800 207472 519200 219024
rect 880 207192 519120 207472
rect 800 195640 519200 207192
rect 880 195360 519120 195640
rect 800 183808 519200 195360
rect 880 183528 519120 183808
rect 800 171976 519200 183528
rect 880 171696 519120 171976
rect 800 160008 519200 171696
rect 880 159728 519120 160008
rect 800 148176 519200 159728
rect 880 147896 519120 148176
rect 800 136344 519200 147896
rect 880 136064 519120 136344
rect 800 124512 519200 136064
rect 880 124232 519120 124512
rect 800 112680 519200 124232
rect 880 112400 519120 112680
rect 800 100848 519200 112400
rect 880 100568 519120 100848
rect 800 89016 519200 100568
rect 880 88736 519120 89016
rect 800 77048 519200 88736
rect 880 76768 519120 77048
rect 800 65216 519200 76768
rect 880 64936 519120 65216
rect 800 53384 519200 64936
rect 880 53104 519120 53384
rect 800 41552 519200 53104
rect 880 41272 519120 41552
rect 800 29720 519200 41272
rect 880 29440 519120 29720
rect 800 17888 519200 29440
rect 880 17608 519120 17888
rect 800 6056 519200 17608
rect 880 5776 519120 6056
rect 800 2143 519200 5776
<< metal4 >>
rect 4208 2128 4528 637616
rect 9328 2128 9648 637616
rect 14448 2128 14768 637616
rect 19568 2128 19888 637616
rect 24688 2128 25008 637616
rect 29808 2128 30128 637616
rect 34928 2128 35248 637616
rect 40048 2128 40368 637616
rect 45168 2128 45488 637616
rect 50288 2128 50608 637616
rect 55408 2128 55728 637616
rect 60528 2128 60848 637616
rect 65648 2128 65968 637616
rect 70768 2128 71088 637616
rect 75888 2128 76208 637616
rect 81008 2128 81328 637616
rect 86128 2128 86448 637616
rect 91248 2128 91568 637616
rect 96368 2128 96688 637616
rect 101488 2128 101808 637616
rect 106608 2128 106928 637616
rect 111728 2128 112048 637616
rect 116848 2128 117168 637616
rect 121968 2128 122288 637616
rect 127088 2128 127408 637616
rect 132208 2128 132528 637616
rect 137328 2128 137648 637616
rect 142448 2128 142768 637616
rect 147568 2128 147888 637616
rect 152688 2128 153008 637616
rect 157808 2128 158128 637616
rect 162928 2128 163248 637616
rect 168048 2128 168368 637616
rect 173168 2128 173488 637616
rect 178288 2128 178608 637616
rect 183408 2128 183728 637616
rect 188528 2128 188848 637616
rect 193648 2128 193968 637616
rect 198768 2128 199088 637616
rect 203888 2128 204208 637616
rect 209008 2128 209328 637616
rect 214128 2128 214448 637616
rect 219248 2128 219568 637616
rect 224368 2128 224688 637616
rect 229488 2128 229808 637616
rect 234608 2128 234928 637616
rect 239728 2128 240048 637616
rect 244848 2128 245168 637616
rect 249968 2128 250288 637616
rect 255088 2128 255408 637616
rect 260208 2128 260528 637616
rect 265328 2128 265648 637616
rect 270448 2128 270768 637616
rect 275568 2128 275888 637616
rect 280688 2128 281008 637616
rect 285808 2128 286128 637616
rect 290928 2128 291248 637616
rect 296048 2128 296368 637616
rect 301168 2128 301488 637616
rect 306288 2128 306608 637616
rect 311408 2128 311728 637616
rect 316528 2128 316848 637616
rect 321648 2128 321968 637616
rect 326768 2128 327088 637616
rect 331888 2128 332208 637616
rect 337008 2128 337328 637616
rect 342128 2128 342448 637616
rect 347248 2128 347568 637616
rect 352368 2128 352688 637616
rect 357488 2128 357808 637616
rect 362608 2128 362928 637616
rect 367728 2128 368048 637616
rect 372848 2128 373168 637616
rect 377968 2128 378288 637616
rect 383088 2128 383408 637616
rect 388208 2128 388528 637616
rect 393328 2128 393648 637616
rect 398448 2128 398768 637616
rect 403568 2128 403888 637616
rect 408688 2128 409008 637616
rect 413808 2128 414128 637616
rect 418928 2128 419248 637616
rect 424048 2128 424368 637616
rect 429168 2128 429488 637616
rect 434288 2128 434608 637616
rect 439408 2128 439728 637616
rect 444528 2128 444848 637616
rect 449648 2128 449968 637616
rect 454768 2128 455088 637616
rect 459888 2128 460208 637616
rect 465008 2128 465328 637616
rect 470128 2128 470448 637616
rect 475248 2128 475568 637616
rect 480368 2128 480688 637616
rect 485488 2128 485808 637616
rect 490608 2128 490928 637616
rect 495728 2128 496048 637616
rect 500848 2128 501168 637616
rect 505968 2128 506288 637616
rect 511088 2128 511408 637616
rect 516208 2128 516528 637616
<< obsm4 >>
rect 3923 3435 4128 629645
rect 4608 3435 9248 629645
rect 9728 3435 14368 629645
rect 14848 3435 19488 629645
rect 19968 3435 24608 629645
rect 25088 3435 29728 629645
rect 30208 3435 34848 629645
rect 35328 3435 39968 629645
rect 40448 3435 45088 629645
rect 45568 3435 50208 629645
rect 50688 3435 55328 629645
rect 55808 3435 60448 629645
rect 60928 3435 65568 629645
rect 66048 3435 70688 629645
rect 71168 3435 75808 629645
rect 76288 3435 80928 629645
rect 81408 3435 86048 629645
rect 86528 3435 91168 629645
rect 91648 3435 96288 629645
rect 96768 3435 101408 629645
rect 101888 3435 106528 629645
rect 107008 3435 111648 629645
rect 112128 3435 116768 629645
rect 117248 3435 121888 629645
rect 122368 3435 127008 629645
rect 127488 3435 132128 629645
rect 132608 3435 137248 629645
rect 137728 3435 142368 629645
rect 142848 3435 147488 629645
rect 147968 3435 152608 629645
rect 153088 3435 157728 629645
rect 158208 3435 162848 629645
rect 163328 3435 167968 629645
rect 168448 3435 173088 629645
rect 173568 3435 178208 629645
rect 178688 3435 183328 629645
rect 183808 3435 188448 629645
rect 188928 3435 193568 629645
rect 194048 3435 198688 629645
rect 199168 3435 203808 629645
rect 204288 3435 208928 629645
rect 209408 3435 214048 629645
rect 214528 3435 219168 629645
rect 219648 3435 224288 629645
rect 224768 3435 229408 629645
rect 229888 3435 234528 629645
rect 235008 3435 239648 629645
rect 240128 3435 244768 629645
rect 245248 3435 249888 629645
rect 250368 3435 255008 629645
rect 255488 3435 260128 629645
rect 260608 3435 265248 629645
rect 265728 3435 270368 629645
rect 270848 3435 275488 629645
rect 275968 3435 280608 629645
rect 281088 3435 285728 629645
rect 286208 3435 290848 629645
rect 291328 3435 295968 629645
rect 296448 3435 301088 629645
rect 301568 3435 306208 629645
rect 306688 3435 311328 629645
rect 311808 3435 316448 629645
rect 316928 3435 321568 629645
rect 322048 3435 326688 629645
rect 327168 3435 331808 629645
rect 332288 3435 336928 629645
rect 337408 3435 342048 629645
rect 342528 3435 347168 629645
rect 347648 3435 352288 629645
rect 352768 3435 357408 629645
rect 357888 3435 362528 629645
rect 363008 3435 367648 629645
rect 368128 3435 372768 629645
rect 373248 3435 377888 629645
rect 378368 3435 383008 629645
rect 383488 3435 388128 629645
rect 388608 3435 393248 629645
rect 393728 3435 398368 629645
rect 398848 3435 403488 629645
rect 403968 3435 408608 629645
rect 409088 3435 413728 629645
rect 414208 3435 418848 629645
rect 419328 3435 423968 629645
rect 424448 3435 429088 629645
rect 429568 3435 434208 629645
rect 434688 3435 439328 629645
rect 439808 3435 444448 629645
rect 444928 3435 449568 629645
rect 450048 3435 454688 629645
rect 455168 3435 459808 629645
rect 460288 3435 464928 629645
rect 465408 3435 470048 629645
rect 470528 3435 475168 629645
rect 475648 3435 480288 629645
rect 480768 3435 485408 629645
rect 485888 3435 490528 629645
rect 491008 3435 495648 629645
rect 496128 3435 500768 629645
rect 501248 3435 505888 629645
rect 506368 3435 511008 629645
rect 511488 3435 516128 629645
rect 516608 3435 517349 629645
<< labels >>
rlabel metal3 s 0 5856 800 5976 6 ipin_x0y1_0
port 1 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 ipin_x0y1_1
port 2 nsew signal input
rlabel metal3 s 0 29520 800 29640 6 ipin_x0y2_0
port 3 nsew signal input
rlabel metal3 s 0 41352 800 41472 6 ipin_x0y2_1
port 4 nsew signal input
rlabel metal3 s 0 53184 800 53304 6 ipin_x0y3_0
port 5 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 ipin_x0y3_1
port 6 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 ipin_x0y4_0
port 7 nsew signal input
rlabel metal3 s 0 88816 800 88936 6 ipin_x0y4_1
port 8 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 ipin_x0y5_0
port 9 nsew signal input
rlabel metal3 s 0 112480 800 112600 6 ipin_x0y5_1
port 10 nsew signal input
rlabel metal3 s 0 124312 800 124432 6 ipin_x0y6_0
port 11 nsew signal input
rlabel metal3 s 0 136144 800 136264 6 ipin_x0y6_1
port 12 nsew signal input
rlabel metal3 s 0 147976 800 148096 6 ipin_x0y7_0
port 13 nsew signal input
rlabel metal3 s 0 159808 800 159928 6 ipin_x0y7_1
port 14 nsew signal input
rlabel metal3 s 0 171776 800 171896 6 ipin_x0y8_0
port 15 nsew signal input
rlabel metal3 s 0 183608 800 183728 6 ipin_x0y8_1
port 16 nsew signal input
rlabel metal3 s 0 195440 800 195560 6 ipin_x0y9_0
port 17 nsew signal input
rlabel metal3 s 0 207272 800 207392 6 ipin_x0y9_1
port 18 nsew signal input
rlabel metal3 s 519200 5856 520000 5976 6 ipin_x10y1_0
port 19 nsew signal input
rlabel metal3 s 519200 17688 520000 17808 6 ipin_x10y1_1
port 20 nsew signal input
rlabel metal3 s 519200 29520 520000 29640 6 ipin_x10y2_0
port 21 nsew signal input
rlabel metal3 s 519200 41352 520000 41472 6 ipin_x10y2_1
port 22 nsew signal input
rlabel metal3 s 519200 53184 520000 53304 6 ipin_x10y3_0
port 23 nsew signal input
rlabel metal3 s 519200 65016 520000 65136 6 ipin_x10y3_1
port 24 nsew signal input
rlabel metal3 s 519200 76848 520000 76968 6 ipin_x10y4_0
port 25 nsew signal input
rlabel metal3 s 519200 88816 520000 88936 6 ipin_x10y4_1
port 26 nsew signal input
rlabel metal3 s 519200 100648 520000 100768 6 ipin_x10y5_0
port 27 nsew signal input
rlabel metal3 s 519200 112480 520000 112600 6 ipin_x10y5_1
port 28 nsew signal input
rlabel metal3 s 519200 124312 520000 124432 6 ipin_x10y6_0
port 29 nsew signal input
rlabel metal3 s 519200 136144 520000 136264 6 ipin_x10y6_1
port 30 nsew signal input
rlabel metal3 s 519200 147976 520000 148096 6 ipin_x10y7_0
port 31 nsew signal input
rlabel metal3 s 519200 159808 520000 159928 6 ipin_x10y7_1
port 32 nsew signal input
rlabel metal3 s 519200 171776 520000 171896 6 ipin_x10y8_0
port 33 nsew signal input
rlabel metal3 s 519200 183608 520000 183728 6 ipin_x10y8_1
port 34 nsew signal input
rlabel metal3 s 519200 195440 520000 195560 6 ipin_x10y9_0
port 35 nsew signal input
rlabel metal3 s 519200 207272 520000 207392 6 ipin_x10y9_1
port 36 nsew signal input
rlabel metal2 s 4802 639200 4858 640000 6 ipin_x1y10_0
port 37 nsew signal input
rlabel metal2 s 14370 639200 14426 640000 6 ipin_x1y10_1
port 38 nsew signal input
rlabel metal2 s 24030 639200 24086 640000 6 ipin_x2y10_0
port 39 nsew signal input
rlabel metal2 s 33690 639200 33746 640000 6 ipin_x2y10_1
port 40 nsew signal input
rlabel metal2 s 43258 639200 43314 640000 6 ipin_x3y10_0
port 41 nsew signal input
rlabel metal2 s 52918 639200 52974 640000 6 ipin_x3y10_1
port 42 nsew signal input
rlabel metal2 s 62578 639200 62634 640000 6 ipin_x4y10_0
port 43 nsew signal input
rlabel metal2 s 72146 639200 72202 640000 6 ipin_x4y10_1
port 44 nsew signal input
rlabel metal2 s 81806 639200 81862 640000 6 ipin_x5y10_0
port 45 nsew signal input
rlabel metal2 s 91466 639200 91522 640000 6 ipin_x5y10_1
port 46 nsew signal input
rlabel metal2 s 101034 639200 101090 640000 6 ipin_x6y10_0
port 47 nsew signal input
rlabel metal2 s 110694 639200 110750 640000 6 ipin_x6y10_1
port 48 nsew signal input
rlabel metal2 s 120354 639200 120410 640000 6 ipin_x7y10_0
port 49 nsew signal input
rlabel metal2 s 129922 639200 129978 640000 6 ipin_x7y10_1
port 50 nsew signal input
rlabel metal2 s 139582 639200 139638 640000 6 ipin_x8y10_0
port 51 nsew signal input
rlabel metal2 s 149242 639200 149298 640000 6 ipin_x8y10_1
port 52 nsew signal input
rlabel metal2 s 158810 639200 158866 640000 6 ipin_x9y10_0
port 53 nsew signal input
rlabel metal2 s 168470 639200 168526 640000 6 ipin_x9y10_1
port 54 nsew signal input
rlabel metal3 s 0 432488 800 432608 6 oeb_x0y1_0
port 55 nsew signal output
rlabel metal3 s 0 444320 800 444440 6 oeb_x0y1_1
port 56 nsew signal output
rlabel metal3 s 0 456152 800 456272 6 oeb_x0y2_0
port 57 nsew signal output
rlabel metal3 s 0 467984 800 468104 6 oeb_x0y2_1
port 58 nsew signal output
rlabel metal3 s 0 479816 800 479936 6 oeb_x0y3_0
port 59 nsew signal output
rlabel metal3 s 0 491784 800 491904 6 oeb_x0y3_1
port 60 nsew signal output
rlabel metal3 s 0 503616 800 503736 6 oeb_x0y4_0
port 61 nsew signal output
rlabel metal3 s 0 515448 800 515568 6 oeb_x0y4_1
port 62 nsew signal output
rlabel metal3 s 0 527280 800 527400 6 oeb_x0y5_0
port 63 nsew signal output
rlabel metal3 s 0 539112 800 539232 6 oeb_x0y5_1
port 64 nsew signal output
rlabel metal3 s 0 550944 800 551064 6 oeb_x0y6_0
port 65 nsew signal output
rlabel metal3 s 0 562776 800 562896 6 oeb_x0y6_1
port 66 nsew signal output
rlabel metal3 s 0 574744 800 574864 6 oeb_x0y7_0
port 67 nsew signal output
rlabel metal3 s 0 586576 800 586696 6 oeb_x0y7_1
port 68 nsew signal output
rlabel metal3 s 0 598408 800 598528 6 oeb_x0y8_0
port 69 nsew signal output
rlabel metal3 s 0 610240 800 610360 6 oeb_x0y8_1
port 70 nsew signal output
rlabel metal3 s 0 622072 800 622192 6 oeb_x0y9_0
port 71 nsew signal output
rlabel metal3 s 0 633904 800 634024 6 oeb_x0y9_1
port 72 nsew signal output
rlabel metal3 s 519200 432488 520000 432608 6 oeb_x10y1_0
port 73 nsew signal output
rlabel metal3 s 519200 444320 520000 444440 6 oeb_x10y1_1
port 74 nsew signal output
rlabel metal3 s 519200 456152 520000 456272 6 oeb_x10y2_0
port 75 nsew signal output
rlabel metal3 s 519200 467984 520000 468104 6 oeb_x10y2_1
port 76 nsew signal output
rlabel metal3 s 519200 479816 520000 479936 6 oeb_x10y3_0
port 77 nsew signal output
rlabel metal3 s 519200 491784 520000 491904 6 oeb_x10y3_1
port 78 nsew signal output
rlabel metal3 s 519200 503616 520000 503736 6 oeb_x10y4_0
port 79 nsew signal output
rlabel metal3 s 519200 515448 520000 515568 6 oeb_x10y4_1
port 80 nsew signal output
rlabel metal3 s 519200 527280 520000 527400 6 oeb_x10y5_0
port 81 nsew signal output
rlabel metal3 s 519200 539112 520000 539232 6 oeb_x10y5_1
port 82 nsew signal output
rlabel metal3 s 519200 550944 520000 551064 6 oeb_x10y6_0
port 83 nsew signal output
rlabel metal3 s 519200 562776 520000 562896 6 oeb_x10y6_1
port 84 nsew signal output
rlabel metal3 s 519200 574744 520000 574864 6 oeb_x10y7_0
port 85 nsew signal output
rlabel metal3 s 519200 586576 520000 586696 6 oeb_x10y7_1
port 86 nsew signal output
rlabel metal3 s 519200 598408 520000 598528 6 oeb_x10y8_0
port 87 nsew signal output
rlabel metal3 s 519200 610240 520000 610360 6 oeb_x10y8_1
port 88 nsew signal output
rlabel metal3 s 519200 622072 520000 622192 6 oeb_x10y9_0
port 89 nsew signal output
rlabel metal3 s 519200 633904 520000 634024 6 oeb_x10y9_1
port 90 nsew signal output
rlabel metal2 s 351458 639200 351514 640000 6 oeb_x1y10_0
port 91 nsew signal output
rlabel metal2 s 361026 639200 361082 640000 6 oeb_x1y10_1
port 92 nsew signal output
rlabel metal2 s 370686 639200 370742 640000 6 oeb_x2y10_0
port 93 nsew signal output
rlabel metal2 s 380346 639200 380402 640000 6 oeb_x2y10_1
port 94 nsew signal output
rlabel metal2 s 389914 639200 389970 640000 6 oeb_x3y10_0
port 95 nsew signal output
rlabel metal2 s 399574 639200 399630 640000 6 oeb_x3y10_1
port 96 nsew signal output
rlabel metal2 s 409234 639200 409290 640000 6 oeb_x4y10_0
port 97 nsew signal output
rlabel metal2 s 418802 639200 418858 640000 6 oeb_x4y10_1
port 98 nsew signal output
rlabel metal2 s 428462 639200 428518 640000 6 oeb_x5y10_0
port 99 nsew signal output
rlabel metal2 s 438122 639200 438178 640000 6 oeb_x5y10_1
port 100 nsew signal output
rlabel metal2 s 447690 639200 447746 640000 6 oeb_x6y10_0
port 101 nsew signal output
rlabel metal2 s 457350 639200 457406 640000 6 oeb_x6y10_1
port 102 nsew signal output
rlabel metal2 s 467010 639200 467066 640000 6 oeb_x7y10_0
port 103 nsew signal output
rlabel metal2 s 476578 639200 476634 640000 6 oeb_x7y10_1
port 104 nsew signal output
rlabel metal2 s 486238 639200 486294 640000 6 oeb_x8y10_0
port 105 nsew signal output
rlabel metal2 s 495898 639200 495954 640000 6 oeb_x8y10_1
port 106 nsew signal output
rlabel metal2 s 505466 639200 505522 640000 6 oeb_x9y10_0
port 107 nsew signal output
rlabel metal2 s 515126 639200 515182 640000 6 oeb_x9y10_1
port 108 nsew signal output
rlabel metal3 s 0 219104 800 219224 6 opin_x0y1_0
port 109 nsew signal output
rlabel metal3 s 0 230936 800 231056 6 opin_x0y1_1
port 110 nsew signal output
rlabel metal3 s 0 242768 800 242888 6 opin_x0y2_0
port 111 nsew signal output
rlabel metal3 s 0 254736 800 254856 6 opin_x0y2_1
port 112 nsew signal output
rlabel metal3 s 0 266568 800 266688 6 opin_x0y3_0
port 113 nsew signal output
rlabel metal3 s 0 278400 800 278520 6 opin_x0y3_1
port 114 nsew signal output
rlabel metal3 s 0 290232 800 290352 6 opin_x0y4_0
port 115 nsew signal output
rlabel metal3 s 0 302064 800 302184 6 opin_x0y4_1
port 116 nsew signal output
rlabel metal3 s 0 313896 800 314016 6 opin_x0y5_0
port 117 nsew signal output
rlabel metal3 s 0 325864 800 325984 6 opin_x0y5_1
port 118 nsew signal output
rlabel metal3 s 0 337696 800 337816 6 opin_x0y6_0
port 119 nsew signal output
rlabel metal3 s 0 349528 800 349648 6 opin_x0y6_1
port 120 nsew signal output
rlabel metal3 s 0 361360 800 361480 6 opin_x0y7_0
port 121 nsew signal output
rlabel metal3 s 0 373192 800 373312 6 opin_x0y7_1
port 122 nsew signal output
rlabel metal3 s 0 385024 800 385144 6 opin_x0y8_0
port 123 nsew signal output
rlabel metal3 s 0 396856 800 396976 6 opin_x0y8_1
port 124 nsew signal output
rlabel metal3 s 0 408824 800 408944 6 opin_x0y9_0
port 125 nsew signal output
rlabel metal3 s 0 420656 800 420776 6 opin_x0y9_1
port 126 nsew signal output
rlabel metal3 s 519200 219104 520000 219224 6 opin_x10y1_0
port 127 nsew signal output
rlabel metal3 s 519200 230936 520000 231056 6 opin_x10y1_1
port 128 nsew signal output
rlabel metal3 s 519200 242768 520000 242888 6 opin_x10y2_0
port 129 nsew signal output
rlabel metal3 s 519200 254736 520000 254856 6 opin_x10y2_1
port 130 nsew signal output
rlabel metal3 s 519200 266568 520000 266688 6 opin_x10y3_0
port 131 nsew signal output
rlabel metal3 s 519200 278400 520000 278520 6 opin_x10y3_1
port 132 nsew signal output
rlabel metal3 s 519200 290232 520000 290352 6 opin_x10y4_0
port 133 nsew signal output
rlabel metal3 s 519200 302064 520000 302184 6 opin_x10y4_1
port 134 nsew signal output
rlabel metal3 s 519200 313896 520000 314016 6 opin_x10y5_0
port 135 nsew signal output
rlabel metal3 s 519200 325864 520000 325984 6 opin_x10y5_1
port 136 nsew signal output
rlabel metal3 s 519200 337696 520000 337816 6 opin_x10y6_0
port 137 nsew signal output
rlabel metal3 s 519200 349528 520000 349648 6 opin_x10y6_1
port 138 nsew signal output
rlabel metal3 s 519200 361360 520000 361480 6 opin_x10y7_0
port 139 nsew signal output
rlabel metal3 s 519200 373192 520000 373312 6 opin_x10y7_1
port 140 nsew signal output
rlabel metal3 s 519200 385024 520000 385144 6 opin_x10y8_0
port 141 nsew signal output
rlabel metal3 s 519200 396856 520000 396976 6 opin_x10y8_1
port 142 nsew signal output
rlabel metal3 s 519200 408824 520000 408944 6 opin_x10y9_0
port 143 nsew signal output
rlabel metal3 s 519200 420656 520000 420776 6 opin_x10y9_1
port 144 nsew signal output
rlabel metal2 s 178130 639200 178186 640000 6 opin_x1y10_0
port 145 nsew signal output
rlabel metal2 s 187698 639200 187754 640000 6 opin_x1y10_1
port 146 nsew signal output
rlabel metal2 s 197358 639200 197414 640000 6 opin_x2y10_0
port 147 nsew signal output
rlabel metal2 s 207018 639200 207074 640000 6 opin_x2y10_1
port 148 nsew signal output
rlabel metal2 s 216586 639200 216642 640000 6 opin_x3y10_0
port 149 nsew signal output
rlabel metal2 s 226246 639200 226302 640000 6 opin_x3y10_1
port 150 nsew signal output
rlabel metal2 s 235906 639200 235962 640000 6 opin_x4y10_0
port 151 nsew signal output
rlabel metal2 s 245474 639200 245530 640000 6 opin_x4y10_1
port 152 nsew signal output
rlabel metal2 s 255134 639200 255190 640000 6 opin_x5y10_0
port 153 nsew signal output
rlabel metal2 s 264794 639200 264850 640000 6 opin_x5y10_1
port 154 nsew signal output
rlabel metal2 s 274362 639200 274418 640000 6 opin_x6y10_0
port 155 nsew signal output
rlabel metal2 s 284022 639200 284078 640000 6 opin_x6y10_1
port 156 nsew signal output
rlabel metal2 s 293682 639200 293738 640000 6 opin_x7y10_0
port 157 nsew signal output
rlabel metal2 s 303250 639200 303306 640000 6 opin_x7y10_1
port 158 nsew signal output
rlabel metal2 s 312910 639200 312966 640000 6 opin_x8y10_0
port 159 nsew signal output
rlabel metal2 s 322570 639200 322626 640000 6 opin_x8y10_1
port 160 nsew signal output
rlabel metal2 s 332138 639200 332194 640000 6 opin_x9y10_0
port 161 nsew signal output
rlabel metal2 s 341798 639200 341854 640000 6 opin_x9y10_1
port 162 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 prog_clk
port 163 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 prog_din
port 164 nsew signal input
rlabel metal2 s 185582 0 185638 800 6 prog_done
port 165 nsew signal input
rlabel metal2 s 259918 0 259974 800 6 prog_dout
port 166 nsew signal output
rlabel metal2 s 334162 0 334218 800 6 prog_rst
port 167 nsew signal input
rlabel metal2 s 408498 0 408554 800 6 prog_we
port 168 nsew signal input
rlabel metal2 s 482742 0 482798 800 6 prog_we_o
port 169 nsew signal output
rlabel metal4 s 4208 2128 4528 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 14448 2128 14768 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 24688 2128 25008 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 34928 2128 35248 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 45168 2128 45488 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 55408 2128 55728 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 65648 2128 65968 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 75888 2128 76208 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 86128 2128 86448 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 96368 2128 96688 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 106608 2128 106928 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 116848 2128 117168 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 127088 2128 127408 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 137328 2128 137648 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 147568 2128 147888 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 157808 2128 158128 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 168048 2128 168368 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 178288 2128 178608 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 188528 2128 188848 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 198768 2128 199088 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 209008 2128 209328 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 219248 2128 219568 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 229488 2128 229808 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 239728 2128 240048 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 249968 2128 250288 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 260208 2128 260528 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 270448 2128 270768 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 280688 2128 281008 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 290928 2128 291248 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 301168 2128 301488 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 311408 2128 311728 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 321648 2128 321968 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 331888 2128 332208 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 342128 2128 342448 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 352368 2128 352688 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 362608 2128 362928 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 372848 2128 373168 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 383088 2128 383408 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 393328 2128 393648 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 403568 2128 403888 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 413808 2128 414128 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 424048 2128 424368 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 434288 2128 434608 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 444528 2128 444848 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 454768 2128 455088 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 465008 2128 465328 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 475248 2128 475568 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 485488 2128 485808 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 495728 2128 496048 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 505968 2128 506288 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 516208 2128 516528 637616 6 vccd1
port 170 nsew power input
rlabel metal4 s 9328 2128 9648 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 19568 2128 19888 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 29808 2128 30128 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 40048 2128 40368 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 50288 2128 50608 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 60528 2128 60848 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 70768 2128 71088 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 81008 2128 81328 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 91248 2128 91568 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 101488 2128 101808 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 111728 2128 112048 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 121968 2128 122288 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 132208 2128 132528 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 142448 2128 142768 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 152688 2128 153008 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 162928 2128 163248 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 173168 2128 173488 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 183408 2128 183728 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 193648 2128 193968 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 203888 2128 204208 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 214128 2128 214448 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 224368 2128 224688 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 234608 2128 234928 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 244848 2128 245168 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 255088 2128 255408 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 265328 2128 265648 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 275568 2128 275888 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 285808 2128 286128 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 296048 2128 296368 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 306288 2128 306608 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 316528 2128 316848 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 326768 2128 327088 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 337008 2128 337328 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 347248 2128 347568 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 357488 2128 357808 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 367728 2128 368048 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 377968 2128 378288 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 388208 2128 388528 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 398448 2128 398768 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 408688 2128 409008 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 418928 2128 419248 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 429168 2128 429488 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 439408 2128 439728 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 449648 2128 449968 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 459888 2128 460208 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 470128 2128 470448 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 480368 2128 480688 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 490608 2128 490928 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 500848 2128 501168 637616 6 vssd1
port 171 nsew ground input
rlabel metal4 s 511088 2128 511408 637616 6 vssd1
port 171 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 520000 640000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 402623354
string GDS_FILE /home/angl/mpw6-prga/caravel/openlane/prga/runs/prga/results/finishing/top.magic.gds
string GDS_START 6276588
<< end >>

