VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO top
  CLASS BLOCK ;
  FOREIGN top ;
  ORIGIN 0.000 0.000 ;
  SIZE 2600.000 BY 3200.000 ;
  PIN ipin_x0y1_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END ipin_x0y1_0
  PIN ipin_x0y1_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END ipin_x0y1_1
  PIN ipin_x0y2_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.600 4.000 148.200 ;
    END
  END ipin_x0y2_0
  PIN ipin_x0y2_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END ipin_x0y2_1
  PIN ipin_x0y3_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.920 4.000 266.520 ;
    END
  END ipin_x0y3_0
  PIN ipin_x0y3_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END ipin_x0y3_1
  PIN ipin_x0y4_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END ipin_x0y4_0
  PIN ipin_x0y4_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.080 4.000 444.680 ;
    END
  END ipin_x0y4_1
  PIN ipin_x0y5_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END ipin_x0y5_0
  PIN ipin_x0y5_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 562.400 4.000 563.000 ;
    END
  END ipin_x0y5_1
  PIN ipin_x0y6_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 621.560 4.000 622.160 ;
    END
  END ipin_x0y6_0
  PIN ipin_x0y6_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.720 4.000 681.320 ;
    END
  END ipin_x0y6_1
  PIN ipin_x0y7_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 739.880 4.000 740.480 ;
    END
  END ipin_x0y7_0
  PIN ipin_x0y7_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.040 4.000 799.640 ;
    END
  END ipin_x0y7_1
  PIN ipin_x0y8_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 858.880 4.000 859.480 ;
    END
  END ipin_x0y8_0
  PIN ipin_x0y8_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 918.040 4.000 918.640 ;
    END
  END ipin_x0y8_1
  PIN ipin_x0y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 977.200 4.000 977.800 ;
    END
  END ipin_x0y9_0
  PIN ipin_x0y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1036.360 4.000 1036.960 ;
    END
  END ipin_x0y9_1
  PIN ipin_x10y1_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 29.280 2600.000 29.880 ;
    END
  END ipin_x10y1_0
  PIN ipin_x10y1_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 88.440 2600.000 89.040 ;
    END
  END ipin_x10y1_1
  PIN ipin_x10y2_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 147.600 2600.000 148.200 ;
    END
  END ipin_x10y2_0
  PIN ipin_x10y2_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 206.760 2600.000 207.360 ;
    END
  END ipin_x10y2_1
  PIN ipin_x10y3_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 265.920 2600.000 266.520 ;
    END
  END ipin_x10y3_0
  PIN ipin_x10y3_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 325.080 2600.000 325.680 ;
    END
  END ipin_x10y3_1
  PIN ipin_x10y4_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 384.240 2600.000 384.840 ;
    END
  END ipin_x10y4_0
  PIN ipin_x10y4_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 444.080 2600.000 444.680 ;
    END
  END ipin_x10y4_1
  PIN ipin_x10y5_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 503.240 2600.000 503.840 ;
    END
  END ipin_x10y5_0
  PIN ipin_x10y5_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 562.400 2600.000 563.000 ;
    END
  END ipin_x10y5_1
  PIN ipin_x10y6_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 621.560 2600.000 622.160 ;
    END
  END ipin_x10y6_0
  PIN ipin_x10y6_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 680.720 2600.000 681.320 ;
    END
  END ipin_x10y6_1
  PIN ipin_x10y7_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 739.880 2600.000 740.480 ;
    END
  END ipin_x10y7_0
  PIN ipin_x10y7_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 799.040 2600.000 799.640 ;
    END
  END ipin_x10y7_1
  PIN ipin_x10y8_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 858.880 2600.000 859.480 ;
    END
  END ipin_x10y8_0
  PIN ipin_x10y8_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 918.040 2600.000 918.640 ;
    END
  END ipin_x10y8_1
  PIN ipin_x10y9_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 977.200 2600.000 977.800 ;
    END
  END ipin_x10y9_0
  PIN ipin_x10y9_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1036.360 2600.000 1036.960 ;
    END
  END ipin_x10y9_1
  PIN ipin_x1y10_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 3196.000 24.290 3200.000 ;
    END
  END ipin_x1y10_0
  PIN ipin_x1y10_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 3196.000 72.130 3200.000 ;
    END
  END ipin_x1y10_1
  PIN ipin_x2y10_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 3196.000 120.430 3200.000 ;
    END
  END ipin_x2y10_0
  PIN ipin_x2y10_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 3196.000 168.730 3200.000 ;
    END
  END ipin_x2y10_1
  PIN ipin_x3y10_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 3196.000 216.570 3200.000 ;
    END
  END ipin_x3y10_0
  PIN ipin_x3y10_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 3196.000 264.870 3200.000 ;
    END
  END ipin_x3y10_1
  PIN ipin_x4y10_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 3196.000 313.170 3200.000 ;
    END
  END ipin_x4y10_0
  PIN ipin_x4y10_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 3196.000 361.010 3200.000 ;
    END
  END ipin_x4y10_1
  PIN ipin_x5y10_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 3196.000 409.310 3200.000 ;
    END
  END ipin_x5y10_0
  PIN ipin_x5y10_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 3196.000 457.610 3200.000 ;
    END
  END ipin_x5y10_1
  PIN ipin_x6y10_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 3196.000 505.450 3200.000 ;
    END
  END ipin_x6y10_0
  PIN ipin_x6y10_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 3196.000 553.750 3200.000 ;
    END
  END ipin_x6y10_1
  PIN ipin_x7y10_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.770 3196.000 602.050 3200.000 ;
    END
  END ipin_x7y10_0
  PIN ipin_x7y10_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 3196.000 649.890 3200.000 ;
    END
  END ipin_x7y10_1
  PIN ipin_x8y10_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.910 3196.000 698.190 3200.000 ;
    END
  END ipin_x8y10_0
  PIN ipin_x8y10_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.210 3196.000 746.490 3200.000 ;
    END
  END ipin_x8y10_1
  PIN ipin_x9y10_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.050 3196.000 794.330 3200.000 ;
    END
  END ipin_x9y10_0
  PIN ipin_x9y10_1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.350 3196.000 842.630 3200.000 ;
    END
  END ipin_x9y10_1
  PIN oeb_x0y1_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2162.440 4.000 2163.040 ;
    END
  END oeb_x0y1_0
  PIN oeb_x0y1_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2221.600 4.000 2222.200 ;
    END
  END oeb_x0y1_1
  PIN oeb_x0y2_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2280.760 4.000 2281.360 ;
    END
  END oeb_x0y2_0
  PIN oeb_x0y2_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2339.920 4.000 2340.520 ;
    END
  END oeb_x0y2_1
  PIN oeb_x0y3_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2399.080 4.000 2399.680 ;
    END
  END oeb_x0y3_0
  PIN oeb_x0y3_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2458.920 4.000 2459.520 ;
    END
  END oeb_x0y3_1
  PIN oeb_x0y4_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2518.080 4.000 2518.680 ;
    END
  END oeb_x0y4_0
  PIN oeb_x0y4_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2577.240 4.000 2577.840 ;
    END
  END oeb_x0y4_1
  PIN oeb_x0y5_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2636.400 4.000 2637.000 ;
    END
  END oeb_x0y5_0
  PIN oeb_x0y5_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2695.560 4.000 2696.160 ;
    END
  END oeb_x0y5_1
  PIN oeb_x0y6_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2754.720 4.000 2755.320 ;
    END
  END oeb_x0y6_0
  PIN oeb_x0y6_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2813.880 4.000 2814.480 ;
    END
  END oeb_x0y6_1
  PIN oeb_x0y7_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2873.720 4.000 2874.320 ;
    END
  END oeb_x0y7_0
  PIN oeb_x0y7_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2932.880 4.000 2933.480 ;
    END
  END oeb_x0y7_1
  PIN oeb_x0y8_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2992.040 4.000 2992.640 ;
    END
  END oeb_x0y8_0
  PIN oeb_x0y8_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3051.200 4.000 3051.800 ;
    END
  END oeb_x0y8_1
  PIN oeb_x0y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3110.360 4.000 3110.960 ;
    END
  END oeb_x0y9_0
  PIN oeb_x0y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3169.520 4.000 3170.120 ;
    END
  END oeb_x0y9_1
  PIN oeb_x10y1_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2162.440 2600.000 2163.040 ;
    END
  END oeb_x10y1_0
  PIN oeb_x10y1_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2221.600 2600.000 2222.200 ;
    END
  END oeb_x10y1_1
  PIN oeb_x10y2_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2280.760 2600.000 2281.360 ;
    END
  END oeb_x10y2_0
  PIN oeb_x10y2_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2339.920 2600.000 2340.520 ;
    END
  END oeb_x10y2_1
  PIN oeb_x10y3_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2399.080 2600.000 2399.680 ;
    END
  END oeb_x10y3_0
  PIN oeb_x10y3_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2458.920 2600.000 2459.520 ;
    END
  END oeb_x10y3_1
  PIN oeb_x10y4_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2518.080 2600.000 2518.680 ;
    END
  END oeb_x10y4_0
  PIN oeb_x10y4_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2577.240 2600.000 2577.840 ;
    END
  END oeb_x10y4_1
  PIN oeb_x10y5_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2636.400 2600.000 2637.000 ;
    END
  END oeb_x10y5_0
  PIN oeb_x10y5_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2695.560 2600.000 2696.160 ;
    END
  END oeb_x10y5_1
  PIN oeb_x10y6_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2754.720 2600.000 2755.320 ;
    END
  END oeb_x10y6_0
  PIN oeb_x10y6_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2813.880 2600.000 2814.480 ;
    END
  END oeb_x10y6_1
  PIN oeb_x10y7_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2873.720 2600.000 2874.320 ;
    END
  END oeb_x10y7_0
  PIN oeb_x10y7_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2932.880 2600.000 2933.480 ;
    END
  END oeb_x10y7_1
  PIN oeb_x10y8_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2992.040 2600.000 2992.640 ;
    END
  END oeb_x10y8_0
  PIN oeb_x10y8_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 3051.200 2600.000 3051.800 ;
    END
  END oeb_x10y8_1
  PIN oeb_x10y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 3110.360 2600.000 3110.960 ;
    END
  END oeb_x10y9_0
  PIN oeb_x10y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 3169.520 2600.000 3170.120 ;
    END
  END oeb_x10y9_1
  PIN oeb_x1y10_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1757.290 3196.000 1757.570 3200.000 ;
    END
  END oeb_x1y10_0
  PIN oeb_x1y10_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.130 3196.000 1805.410 3200.000 ;
    END
  END oeb_x1y10_1
  PIN oeb_x2y10_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1853.430 3196.000 1853.710 3200.000 ;
    END
  END oeb_x2y10_0
  PIN oeb_x2y10_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1901.730 3196.000 1902.010 3200.000 ;
    END
  END oeb_x2y10_1
  PIN oeb_x3y10_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1949.570 3196.000 1949.850 3200.000 ;
    END
  END oeb_x3y10_0
  PIN oeb_x3y10_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1997.870 3196.000 1998.150 3200.000 ;
    END
  END oeb_x3y10_1
  PIN oeb_x4y10_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2046.170 3196.000 2046.450 3200.000 ;
    END
  END oeb_x4y10_0
  PIN oeb_x4y10_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2094.010 3196.000 2094.290 3200.000 ;
    END
  END oeb_x4y10_1
  PIN oeb_x5y10_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2142.310 3196.000 2142.590 3200.000 ;
    END
  END oeb_x5y10_0
  PIN oeb_x5y10_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2190.610 3196.000 2190.890 3200.000 ;
    END
  END oeb_x5y10_1
  PIN oeb_x6y10_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2238.450 3196.000 2238.730 3200.000 ;
    END
  END oeb_x6y10_0
  PIN oeb_x6y10_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2286.750 3196.000 2287.030 3200.000 ;
    END
  END oeb_x6y10_1
  PIN oeb_x7y10_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2335.050 3196.000 2335.330 3200.000 ;
    END
  END oeb_x7y10_0
  PIN oeb_x7y10_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2382.890 3196.000 2383.170 3200.000 ;
    END
  END oeb_x7y10_1
  PIN oeb_x8y10_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.190 3196.000 2431.470 3200.000 ;
    END
  END oeb_x8y10_0
  PIN oeb_x8y10_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2479.490 3196.000 2479.770 3200.000 ;
    END
  END oeb_x8y10_1
  PIN oeb_x9y10_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2527.330 3196.000 2527.610 3200.000 ;
    END
  END oeb_x9y10_0
  PIN oeb_x9y10_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2575.630 3196.000 2575.910 3200.000 ;
    END
  END oeb_x9y10_1
  PIN opin_x0y1_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1095.520 4.000 1096.120 ;
    END
  END opin_x0y1_0
  PIN opin_x0y1_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1154.680 4.000 1155.280 ;
    END
  END opin_x0y1_1
  PIN opin_x0y2_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1213.840 4.000 1214.440 ;
    END
  END opin_x0y2_0
  PIN opin_x0y2_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1273.680 4.000 1274.280 ;
    END
  END opin_x0y2_1
  PIN opin_x0y3_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1332.840 4.000 1333.440 ;
    END
  END opin_x0y3_0
  PIN opin_x0y3_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1392.000 4.000 1392.600 ;
    END
  END opin_x0y3_1
  PIN opin_x0y4_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1451.160 4.000 1451.760 ;
    END
  END opin_x0y4_0
  PIN opin_x0y4_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1510.320 4.000 1510.920 ;
    END
  END opin_x0y4_1
  PIN opin_x0y5_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1569.480 4.000 1570.080 ;
    END
  END opin_x0y5_0
  PIN opin_x0y5_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1629.320 4.000 1629.920 ;
    END
  END opin_x0y5_1
  PIN opin_x0y6_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1688.480 4.000 1689.080 ;
    END
  END opin_x0y6_0
  PIN opin_x0y6_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1747.640 4.000 1748.240 ;
    END
  END opin_x0y6_1
  PIN opin_x0y7_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1806.800 4.000 1807.400 ;
    END
  END opin_x0y7_0
  PIN opin_x0y7_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1865.960 4.000 1866.560 ;
    END
  END opin_x0y7_1
  PIN opin_x0y8_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1925.120 4.000 1925.720 ;
    END
  END opin_x0y8_0
  PIN opin_x0y8_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1984.280 4.000 1984.880 ;
    END
  END opin_x0y8_1
  PIN opin_x0y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2044.120 4.000 2044.720 ;
    END
  END opin_x0y9_0
  PIN opin_x0y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2103.280 4.000 2103.880 ;
    END
  END opin_x0y9_1
  PIN opin_x10y1_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1095.520 2600.000 1096.120 ;
    END
  END opin_x10y1_0
  PIN opin_x10y1_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1154.680 2600.000 1155.280 ;
    END
  END opin_x10y1_1
  PIN opin_x10y2_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1213.840 2600.000 1214.440 ;
    END
  END opin_x10y2_0
  PIN opin_x10y2_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1273.680 2600.000 1274.280 ;
    END
  END opin_x10y2_1
  PIN opin_x10y3_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1332.840 2600.000 1333.440 ;
    END
  END opin_x10y3_0
  PIN opin_x10y3_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1392.000 2600.000 1392.600 ;
    END
  END opin_x10y3_1
  PIN opin_x10y4_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1451.160 2600.000 1451.760 ;
    END
  END opin_x10y4_0
  PIN opin_x10y4_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1510.320 2600.000 1510.920 ;
    END
  END opin_x10y4_1
  PIN opin_x10y5_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1569.480 2600.000 1570.080 ;
    END
  END opin_x10y5_0
  PIN opin_x10y5_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1629.320 2600.000 1629.920 ;
    END
  END opin_x10y5_1
  PIN opin_x10y6_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1688.480 2600.000 1689.080 ;
    END
  END opin_x10y6_0
  PIN opin_x10y6_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1747.640 2600.000 1748.240 ;
    END
  END opin_x10y6_1
  PIN opin_x10y7_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1806.800 2600.000 1807.400 ;
    END
  END opin_x10y7_0
  PIN opin_x10y7_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1865.960 2600.000 1866.560 ;
    END
  END opin_x10y7_1
  PIN opin_x10y8_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1925.120 2600.000 1925.720 ;
    END
  END opin_x10y8_0
  PIN opin_x10y8_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 1984.280 2600.000 1984.880 ;
    END
  END opin_x10y8_1
  PIN opin_x10y9_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2044.120 2600.000 2044.720 ;
    END
  END opin_x10y9_0
  PIN opin_x10y9_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2596.000 2103.280 2600.000 2103.880 ;
    END
  END opin_x10y9_1
  PIN opin_x1y10_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.650 3196.000 890.930 3200.000 ;
    END
  END opin_x1y10_0
  PIN opin_x1y10_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.490 3196.000 938.770 3200.000 ;
    END
  END opin_x1y10_1
  PIN opin_x2y10_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.790 3196.000 987.070 3200.000 ;
    END
  END opin_x2y10_0
  PIN opin_x2y10_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1035.090 3196.000 1035.370 3200.000 ;
    END
  END opin_x2y10_1
  PIN opin_x3y10_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.930 3196.000 1083.210 3200.000 ;
    END
  END opin_x3y10_0
  PIN opin_x3y10_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.230 3196.000 1131.510 3200.000 ;
    END
  END opin_x3y10_1
  PIN opin_x4y10_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.530 3196.000 1179.810 3200.000 ;
    END
  END opin_x4y10_0
  PIN opin_x4y10_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.370 3196.000 1227.650 3200.000 ;
    END
  END opin_x4y10_1
  PIN opin_x5y10_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.670 3196.000 1275.950 3200.000 ;
    END
  END opin_x5y10_0
  PIN opin_x5y10_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.970 3196.000 1324.250 3200.000 ;
    END
  END opin_x5y10_1
  PIN opin_x6y10_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.810 3196.000 1372.090 3200.000 ;
    END
  END opin_x6y10_0
  PIN opin_x6y10_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.110 3196.000 1420.390 3200.000 ;
    END
  END opin_x6y10_1
  PIN opin_x7y10_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.410 3196.000 1468.690 3200.000 ;
    END
  END opin_x7y10_0
  PIN opin_x7y10_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1516.250 3196.000 1516.530 3200.000 ;
    END
  END opin_x7y10_1
  PIN opin_x8y10_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1564.550 3196.000 1564.830 3200.000 ;
    END
  END opin_x8y10_0
  PIN opin_x8y10_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1612.850 3196.000 1613.130 3200.000 ;
    END
  END opin_x8y10_1
  PIN opin_x9y10_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1660.690 3196.000 1660.970 3200.000 ;
    END
  END opin_x9y10_0
  PIN opin_x9y10_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1708.990 3196.000 1709.270 3200.000 ;
    END
  END opin_x9y10_1
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END prog_clk
  PIN prog_din
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 0.000 556.970 4.000 ;
    END
  END prog_din
  PIN prog_done
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.910 0.000 928.190 4.000 ;
    END
  END prog_done
  PIN prog_dout
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1299.590 0.000 1299.870 4.000 ;
    END
  END prog_dout
  PIN prog_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1670.810 0.000 1671.090 4.000 ;
    END
  END prog_rst
  PIN prog_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2042.490 0.000 2042.770 4.000 ;
    END
  END prog_we
  PIN prog_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2413.710 0.000 2413.990 4.000 ;
    END
  END prog_we_o
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 72.240 10.640 73.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 123.440 10.640 125.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 225.840 10.640 227.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 277.040 10.640 278.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 379.440 10.640 381.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 430.640 10.640 432.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 533.040 10.640 534.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 584.240 10.640 585.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 686.640 10.640 688.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 737.840 10.640 739.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 840.240 10.640 841.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 891.440 10.640 893.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 993.840 10.640 995.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1045.040 10.640 1046.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1147.440 10.640 1149.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1198.640 10.640 1200.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1301.040 10.640 1302.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1352.240 10.640 1353.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1454.640 10.640 1456.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1505.840 10.640 1507.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1608.240 10.640 1609.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1659.440 10.640 1661.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1761.840 10.640 1763.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1813.040 10.640 1814.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1915.440 10.640 1917.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1966.640 10.640 1968.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2069.040 10.640 2070.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2120.240 10.640 2121.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2222.640 10.640 2224.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2273.840 10.640 2275.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.240 10.640 2377.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2427.440 10.640 2429.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2529.840 10.640 2531.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2581.040 10.640 2582.640 3188.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 46.640 10.640 48.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 149.040 10.640 150.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 200.240 10.640 201.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 302.640 10.640 304.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 353.840 10.640 355.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 456.240 10.640 457.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 507.440 10.640 509.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 609.840 10.640 611.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 661.040 10.640 662.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 763.440 10.640 765.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 814.640 10.640 816.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 917.040 10.640 918.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 968.240 10.640 969.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1070.640 10.640 1072.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1121.840 10.640 1123.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1224.240 10.640 1225.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1275.440 10.640 1277.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1377.840 10.640 1379.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1429.040 10.640 1430.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1531.440 10.640 1533.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1582.640 10.640 1584.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1685.040 10.640 1686.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.240 10.640 1737.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1838.640 10.640 1840.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1889.840 10.640 1891.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1992.240 10.640 1993.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2043.440 10.640 2045.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2145.840 10.640 2147.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2197.040 10.640 2198.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2299.440 10.640 2301.040 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2350.640 10.640 2352.240 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2453.040 10.640 2454.640 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2504.240 10.640 2505.840 3188.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 2555.440 10.640 2557.040 3188.080 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2594.400 3187.925 ;
      LAYER met1 ;
        RECT 5.520 10.640 2599.850 3188.080 ;
      LAYER met2 ;
        RECT 6.080 3195.720 23.730 3196.410 ;
        RECT 24.570 3195.720 71.570 3196.410 ;
        RECT 72.410 3195.720 119.870 3196.410 ;
        RECT 120.710 3195.720 168.170 3196.410 ;
        RECT 169.010 3195.720 216.010 3196.410 ;
        RECT 216.850 3195.720 264.310 3196.410 ;
        RECT 265.150 3195.720 312.610 3196.410 ;
        RECT 313.450 3195.720 360.450 3196.410 ;
        RECT 361.290 3195.720 408.750 3196.410 ;
        RECT 409.590 3195.720 457.050 3196.410 ;
        RECT 457.890 3195.720 504.890 3196.410 ;
        RECT 505.730 3195.720 553.190 3196.410 ;
        RECT 554.030 3195.720 601.490 3196.410 ;
        RECT 602.330 3195.720 649.330 3196.410 ;
        RECT 650.170 3195.720 697.630 3196.410 ;
        RECT 698.470 3195.720 745.930 3196.410 ;
        RECT 746.770 3195.720 793.770 3196.410 ;
        RECT 794.610 3195.720 842.070 3196.410 ;
        RECT 842.910 3195.720 890.370 3196.410 ;
        RECT 891.210 3195.720 938.210 3196.410 ;
        RECT 939.050 3195.720 986.510 3196.410 ;
        RECT 987.350 3195.720 1034.810 3196.410 ;
        RECT 1035.650 3195.720 1082.650 3196.410 ;
        RECT 1083.490 3195.720 1130.950 3196.410 ;
        RECT 1131.790 3195.720 1179.250 3196.410 ;
        RECT 1180.090 3195.720 1227.090 3196.410 ;
        RECT 1227.930 3195.720 1275.390 3196.410 ;
        RECT 1276.230 3195.720 1323.690 3196.410 ;
        RECT 1324.530 3195.720 1371.530 3196.410 ;
        RECT 1372.370 3195.720 1419.830 3196.410 ;
        RECT 1420.670 3195.720 1468.130 3196.410 ;
        RECT 1468.970 3195.720 1515.970 3196.410 ;
        RECT 1516.810 3195.720 1564.270 3196.410 ;
        RECT 1565.110 3195.720 1612.570 3196.410 ;
        RECT 1613.410 3195.720 1660.410 3196.410 ;
        RECT 1661.250 3195.720 1708.710 3196.410 ;
        RECT 1709.550 3195.720 1757.010 3196.410 ;
        RECT 1757.850 3195.720 1804.850 3196.410 ;
        RECT 1805.690 3195.720 1853.150 3196.410 ;
        RECT 1853.990 3195.720 1901.450 3196.410 ;
        RECT 1902.290 3195.720 1949.290 3196.410 ;
        RECT 1950.130 3195.720 1997.590 3196.410 ;
        RECT 1998.430 3195.720 2045.890 3196.410 ;
        RECT 2046.730 3195.720 2093.730 3196.410 ;
        RECT 2094.570 3195.720 2142.030 3196.410 ;
        RECT 2142.870 3195.720 2190.330 3196.410 ;
        RECT 2191.170 3195.720 2238.170 3196.410 ;
        RECT 2239.010 3195.720 2286.470 3196.410 ;
        RECT 2287.310 3195.720 2334.770 3196.410 ;
        RECT 2335.610 3195.720 2382.610 3196.410 ;
        RECT 2383.450 3195.720 2430.910 3196.410 ;
        RECT 2431.750 3195.720 2479.210 3196.410 ;
        RECT 2480.050 3195.720 2527.050 3196.410 ;
        RECT 2527.890 3195.720 2575.350 3196.410 ;
        RECT 2576.190 3195.720 2599.820 3196.410 ;
        RECT 6.080 4.280 2599.820 3195.720 ;
        RECT 6.080 4.000 185.190 4.280 ;
        RECT 186.030 4.000 556.410 4.280 ;
        RECT 557.250 4.000 927.630 4.280 ;
        RECT 928.470 4.000 1299.310 4.280 ;
        RECT 1300.150 4.000 1670.530 4.280 ;
        RECT 1671.370 4.000 2042.210 4.280 ;
        RECT 2043.050 4.000 2413.430 4.280 ;
        RECT 2414.270 4.000 2599.820 4.280 ;
      LAYER met3 ;
        RECT 4.000 3170.520 2596.000 3188.005 ;
        RECT 4.400 3169.120 2595.600 3170.520 ;
        RECT 4.000 3111.360 2596.000 3169.120 ;
        RECT 4.400 3109.960 2595.600 3111.360 ;
        RECT 4.000 3052.200 2596.000 3109.960 ;
        RECT 4.400 3050.800 2595.600 3052.200 ;
        RECT 4.000 2993.040 2596.000 3050.800 ;
        RECT 4.400 2991.640 2595.600 2993.040 ;
        RECT 4.000 2933.880 2596.000 2991.640 ;
        RECT 4.400 2932.480 2595.600 2933.880 ;
        RECT 4.000 2874.720 2596.000 2932.480 ;
        RECT 4.400 2873.320 2595.600 2874.720 ;
        RECT 4.000 2814.880 2596.000 2873.320 ;
        RECT 4.400 2813.480 2595.600 2814.880 ;
        RECT 4.000 2755.720 2596.000 2813.480 ;
        RECT 4.400 2754.320 2595.600 2755.720 ;
        RECT 4.000 2696.560 2596.000 2754.320 ;
        RECT 4.400 2695.160 2595.600 2696.560 ;
        RECT 4.000 2637.400 2596.000 2695.160 ;
        RECT 4.400 2636.000 2595.600 2637.400 ;
        RECT 4.000 2578.240 2596.000 2636.000 ;
        RECT 4.400 2576.840 2595.600 2578.240 ;
        RECT 4.000 2519.080 2596.000 2576.840 ;
        RECT 4.400 2517.680 2595.600 2519.080 ;
        RECT 4.000 2459.920 2596.000 2517.680 ;
        RECT 4.400 2458.520 2595.600 2459.920 ;
        RECT 4.000 2400.080 2596.000 2458.520 ;
        RECT 4.400 2398.680 2595.600 2400.080 ;
        RECT 4.000 2340.920 2596.000 2398.680 ;
        RECT 4.400 2339.520 2595.600 2340.920 ;
        RECT 4.000 2281.760 2596.000 2339.520 ;
        RECT 4.400 2280.360 2595.600 2281.760 ;
        RECT 4.000 2222.600 2596.000 2280.360 ;
        RECT 4.400 2221.200 2595.600 2222.600 ;
        RECT 4.000 2163.440 2596.000 2221.200 ;
        RECT 4.400 2162.040 2595.600 2163.440 ;
        RECT 4.000 2104.280 2596.000 2162.040 ;
        RECT 4.400 2102.880 2595.600 2104.280 ;
        RECT 4.000 2045.120 2596.000 2102.880 ;
        RECT 4.400 2043.720 2595.600 2045.120 ;
        RECT 4.000 1985.280 2596.000 2043.720 ;
        RECT 4.400 1983.880 2595.600 1985.280 ;
        RECT 4.000 1926.120 2596.000 1983.880 ;
        RECT 4.400 1924.720 2595.600 1926.120 ;
        RECT 4.000 1866.960 2596.000 1924.720 ;
        RECT 4.400 1865.560 2595.600 1866.960 ;
        RECT 4.000 1807.800 2596.000 1865.560 ;
        RECT 4.400 1806.400 2595.600 1807.800 ;
        RECT 4.000 1748.640 2596.000 1806.400 ;
        RECT 4.400 1747.240 2595.600 1748.640 ;
        RECT 4.000 1689.480 2596.000 1747.240 ;
        RECT 4.400 1688.080 2595.600 1689.480 ;
        RECT 4.000 1630.320 2596.000 1688.080 ;
        RECT 4.400 1628.920 2595.600 1630.320 ;
        RECT 4.000 1570.480 2596.000 1628.920 ;
        RECT 4.400 1569.080 2595.600 1570.480 ;
        RECT 4.000 1511.320 2596.000 1569.080 ;
        RECT 4.400 1509.920 2595.600 1511.320 ;
        RECT 4.000 1452.160 2596.000 1509.920 ;
        RECT 4.400 1450.760 2595.600 1452.160 ;
        RECT 4.000 1393.000 2596.000 1450.760 ;
        RECT 4.400 1391.600 2595.600 1393.000 ;
        RECT 4.000 1333.840 2596.000 1391.600 ;
        RECT 4.400 1332.440 2595.600 1333.840 ;
        RECT 4.000 1274.680 2596.000 1332.440 ;
        RECT 4.400 1273.280 2595.600 1274.680 ;
        RECT 4.000 1214.840 2596.000 1273.280 ;
        RECT 4.400 1213.440 2595.600 1214.840 ;
        RECT 4.000 1155.680 2596.000 1213.440 ;
        RECT 4.400 1154.280 2595.600 1155.680 ;
        RECT 4.000 1096.520 2596.000 1154.280 ;
        RECT 4.400 1095.120 2595.600 1096.520 ;
        RECT 4.000 1037.360 2596.000 1095.120 ;
        RECT 4.400 1035.960 2595.600 1037.360 ;
        RECT 4.000 978.200 2596.000 1035.960 ;
        RECT 4.400 976.800 2595.600 978.200 ;
        RECT 4.000 919.040 2596.000 976.800 ;
        RECT 4.400 917.640 2595.600 919.040 ;
        RECT 4.000 859.880 2596.000 917.640 ;
        RECT 4.400 858.480 2595.600 859.880 ;
        RECT 4.000 800.040 2596.000 858.480 ;
        RECT 4.400 798.640 2595.600 800.040 ;
        RECT 4.000 740.880 2596.000 798.640 ;
        RECT 4.400 739.480 2595.600 740.880 ;
        RECT 4.000 681.720 2596.000 739.480 ;
        RECT 4.400 680.320 2595.600 681.720 ;
        RECT 4.000 622.560 2596.000 680.320 ;
        RECT 4.400 621.160 2595.600 622.560 ;
        RECT 4.000 563.400 2596.000 621.160 ;
        RECT 4.400 562.000 2595.600 563.400 ;
        RECT 4.000 504.240 2596.000 562.000 ;
        RECT 4.400 502.840 2595.600 504.240 ;
        RECT 4.000 445.080 2596.000 502.840 ;
        RECT 4.400 443.680 2595.600 445.080 ;
        RECT 4.000 385.240 2596.000 443.680 ;
        RECT 4.400 383.840 2595.600 385.240 ;
        RECT 4.000 326.080 2596.000 383.840 ;
        RECT 4.400 324.680 2595.600 326.080 ;
        RECT 4.000 266.920 2596.000 324.680 ;
        RECT 4.400 265.520 2595.600 266.920 ;
        RECT 4.000 207.760 2596.000 265.520 ;
        RECT 4.400 206.360 2595.600 207.760 ;
        RECT 4.000 148.600 2596.000 206.360 ;
        RECT 4.400 147.200 2595.600 148.600 ;
        RECT 4.000 89.440 2596.000 147.200 ;
        RECT 4.400 88.040 2595.600 89.440 ;
        RECT 4.000 30.280 2596.000 88.040 ;
        RECT 4.400 28.880 2595.600 30.280 ;
        RECT 4.000 10.715 2596.000 28.880 ;
      LAYER met4 ;
        RECT 19.615 17.175 20.640 3148.225 ;
        RECT 23.040 17.175 46.240 3148.225 ;
        RECT 48.640 17.175 71.840 3148.225 ;
        RECT 74.240 17.175 97.440 3148.225 ;
        RECT 99.840 17.175 123.040 3148.225 ;
        RECT 125.440 17.175 148.640 3148.225 ;
        RECT 151.040 17.175 174.240 3148.225 ;
        RECT 176.640 17.175 199.840 3148.225 ;
        RECT 202.240 17.175 225.440 3148.225 ;
        RECT 227.840 17.175 251.040 3148.225 ;
        RECT 253.440 17.175 276.640 3148.225 ;
        RECT 279.040 17.175 302.240 3148.225 ;
        RECT 304.640 17.175 327.840 3148.225 ;
        RECT 330.240 17.175 353.440 3148.225 ;
        RECT 355.840 17.175 379.040 3148.225 ;
        RECT 381.440 17.175 404.640 3148.225 ;
        RECT 407.040 17.175 430.240 3148.225 ;
        RECT 432.640 17.175 455.840 3148.225 ;
        RECT 458.240 17.175 481.440 3148.225 ;
        RECT 483.840 17.175 507.040 3148.225 ;
        RECT 509.440 17.175 532.640 3148.225 ;
        RECT 535.040 17.175 558.240 3148.225 ;
        RECT 560.640 17.175 583.840 3148.225 ;
        RECT 586.240 17.175 609.440 3148.225 ;
        RECT 611.840 17.175 635.040 3148.225 ;
        RECT 637.440 17.175 660.640 3148.225 ;
        RECT 663.040 17.175 686.240 3148.225 ;
        RECT 688.640 17.175 711.840 3148.225 ;
        RECT 714.240 17.175 737.440 3148.225 ;
        RECT 739.840 17.175 763.040 3148.225 ;
        RECT 765.440 17.175 788.640 3148.225 ;
        RECT 791.040 17.175 814.240 3148.225 ;
        RECT 816.640 17.175 839.840 3148.225 ;
        RECT 842.240 17.175 865.440 3148.225 ;
        RECT 867.840 17.175 891.040 3148.225 ;
        RECT 893.440 17.175 916.640 3148.225 ;
        RECT 919.040 17.175 942.240 3148.225 ;
        RECT 944.640 17.175 967.840 3148.225 ;
        RECT 970.240 17.175 993.440 3148.225 ;
        RECT 995.840 17.175 1019.040 3148.225 ;
        RECT 1021.440 17.175 1044.640 3148.225 ;
        RECT 1047.040 17.175 1070.240 3148.225 ;
        RECT 1072.640 17.175 1095.840 3148.225 ;
        RECT 1098.240 17.175 1121.440 3148.225 ;
        RECT 1123.840 17.175 1147.040 3148.225 ;
        RECT 1149.440 17.175 1172.640 3148.225 ;
        RECT 1175.040 17.175 1198.240 3148.225 ;
        RECT 1200.640 17.175 1223.840 3148.225 ;
        RECT 1226.240 17.175 1249.440 3148.225 ;
        RECT 1251.840 17.175 1275.040 3148.225 ;
        RECT 1277.440 17.175 1300.640 3148.225 ;
        RECT 1303.040 17.175 1326.240 3148.225 ;
        RECT 1328.640 17.175 1351.840 3148.225 ;
        RECT 1354.240 17.175 1377.440 3148.225 ;
        RECT 1379.840 17.175 1403.040 3148.225 ;
        RECT 1405.440 17.175 1428.640 3148.225 ;
        RECT 1431.040 17.175 1454.240 3148.225 ;
        RECT 1456.640 17.175 1479.840 3148.225 ;
        RECT 1482.240 17.175 1505.440 3148.225 ;
        RECT 1507.840 17.175 1531.040 3148.225 ;
        RECT 1533.440 17.175 1556.640 3148.225 ;
        RECT 1559.040 17.175 1582.240 3148.225 ;
        RECT 1584.640 17.175 1607.840 3148.225 ;
        RECT 1610.240 17.175 1633.440 3148.225 ;
        RECT 1635.840 17.175 1659.040 3148.225 ;
        RECT 1661.440 17.175 1684.640 3148.225 ;
        RECT 1687.040 17.175 1710.240 3148.225 ;
        RECT 1712.640 17.175 1735.840 3148.225 ;
        RECT 1738.240 17.175 1761.440 3148.225 ;
        RECT 1763.840 17.175 1787.040 3148.225 ;
        RECT 1789.440 17.175 1812.640 3148.225 ;
        RECT 1815.040 17.175 1838.240 3148.225 ;
        RECT 1840.640 17.175 1863.840 3148.225 ;
        RECT 1866.240 17.175 1889.440 3148.225 ;
        RECT 1891.840 17.175 1915.040 3148.225 ;
        RECT 1917.440 17.175 1940.640 3148.225 ;
        RECT 1943.040 17.175 1966.240 3148.225 ;
        RECT 1968.640 17.175 1991.840 3148.225 ;
        RECT 1994.240 17.175 2017.440 3148.225 ;
        RECT 2019.840 17.175 2043.040 3148.225 ;
        RECT 2045.440 17.175 2068.640 3148.225 ;
        RECT 2071.040 17.175 2094.240 3148.225 ;
        RECT 2096.640 17.175 2119.840 3148.225 ;
        RECT 2122.240 17.175 2145.440 3148.225 ;
        RECT 2147.840 17.175 2171.040 3148.225 ;
        RECT 2173.440 17.175 2196.640 3148.225 ;
        RECT 2199.040 17.175 2222.240 3148.225 ;
        RECT 2224.640 17.175 2247.840 3148.225 ;
        RECT 2250.240 17.175 2273.440 3148.225 ;
        RECT 2275.840 17.175 2299.040 3148.225 ;
        RECT 2301.440 17.175 2324.640 3148.225 ;
        RECT 2327.040 17.175 2350.240 3148.225 ;
        RECT 2352.640 17.175 2375.840 3148.225 ;
        RECT 2378.240 17.175 2401.440 3148.225 ;
        RECT 2403.840 17.175 2427.040 3148.225 ;
        RECT 2429.440 17.175 2452.640 3148.225 ;
        RECT 2455.040 17.175 2478.240 3148.225 ;
        RECT 2480.640 17.175 2503.840 3148.225 ;
        RECT 2506.240 17.175 2529.440 3148.225 ;
        RECT 2531.840 17.175 2555.040 3148.225 ;
        RECT 2557.440 17.175 2580.640 3148.225 ;
        RECT 2583.040 17.175 2586.745 3148.225 ;
  END
END top
END LIBRARY

