// SPDX-FileCopyrightText: 2022 Princeton University
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

// Automatically generated by PRGA's RTL generator
module top (
`ifdef USE_POWER_PINS
    inout vccd1,	// User area 1 1.8V supply
    inout vssd1,	// User area 1 digital ground
`endif
    input wire [0:0] ipin_x0y1_0
    , output wire [0:0] opin_x0y1_0
    , output wire [0:0] oe_x0y1_0
    , input wire [0:0] ipin_x0y1_1
    , output wire [0:0] opin_x0y1_1
    , output wire [0:0] oe_x0y1_1
    , input wire [0:0] ipin_x0y2_0
    , output wire [0:0] opin_x0y2_0
    , output wire [0:0] oe_x0y2_0
    , input wire [0:0] ipin_x0y2_1
    , output wire [0:0] opin_x0y2_1
    , output wire [0:0] oe_x0y2_1
    , input wire [0:0] ipin_x0y3_0
    , output wire [0:0] opin_x0y3_0
    , output wire [0:0] oe_x0y3_0
    , input wire [0:0] ipin_x0y3_1
    , output wire [0:0] opin_x0y3_1
    , output wire [0:0] oe_x0y3_1
    , input wire [0:0] ipin_x0y4_0
    , output wire [0:0] opin_x0y4_0
    , output wire [0:0] oe_x0y4_0
    , input wire [0:0] ipin_x0y4_1
    , output wire [0:0] opin_x0y4_1
    , output wire [0:0] oe_x0y4_1
    , input wire [0:0] ipin_x0y5_0
    , output wire [0:0] opin_x0y5_0
    , output wire [0:0] oe_x0y5_0
    , input wire [0:0] ipin_x0y5_1
    , output wire [0:0] opin_x0y5_1
    , output wire [0:0] oe_x0y5_1
    , input wire [0:0] ipin_x0y6_0
    , output wire [0:0] opin_x0y6_0
    , output wire [0:0] oe_x0y6_0
    , input wire [0:0] ipin_x0y6_1
    , output wire [0:0] opin_x0y6_1
    , output wire [0:0] oe_x0y6_1
    , input wire [0:0] ipin_x0y7_0
    , output wire [0:0] opin_x0y7_0
    , output wire [0:0] oe_x0y7_0
    , input wire [0:0] ipin_x0y7_1
    , output wire [0:0] opin_x0y7_1
    , output wire [0:0] oe_x0y7_1
    , input wire [0:0] ipin_x0y8_0
    , output wire [0:0] opin_x0y8_0
    , output wire [0:0] oe_x0y8_0
    , input wire [0:0] ipin_x0y8_1
    , output wire [0:0] opin_x0y8_1
    , output wire [0:0] oe_x0y8_1
    , input wire [0:0] ipin_x1y9_0
    , output wire [0:0] opin_x1y9_0
    , output wire [0:0] oe_x1y9_0
    , input wire [0:0] ipin_x1y9_1
    , output wire [0:0] opin_x1y9_1
    , output wire [0:0] oe_x1y9_1
    , input wire [0:0] ipin_x2y9_0
    , output wire [0:0] opin_x2y9_0
    , output wire [0:0] oe_x2y9_0
    , input wire [0:0] ipin_x2y9_1
    , output wire [0:0] opin_x2y9_1
    , output wire [0:0] oe_x2y9_1
    , input wire [0:0] ipin_x3y9_0
    , output wire [0:0] opin_x3y9_0
    , output wire [0:0] oe_x3y9_0
    , input wire [0:0] ipin_x3y9_1
    , output wire [0:0] opin_x3y9_1
    , output wire [0:0] oe_x3y9_1
    , input wire [0:0] ipin_x4y9_0
    , output wire [0:0] opin_x4y9_0
    , output wire [0:0] oe_x4y9_0
    , input wire [0:0] ipin_x4y9_1
    , output wire [0:0] opin_x4y9_1
    , output wire [0:0] oe_x4y9_1
    , input wire [0:0] ipin_x5y9_0
    , output wire [0:0] opin_x5y9_0
    , output wire [0:0] oe_x5y9_0
    , input wire [0:0] ipin_x5y9_1
    , output wire [0:0] opin_x5y9_1
    , output wire [0:0] oe_x5y9_1
    , input wire [0:0] ipin_x6y9_0
    , output wire [0:0] opin_x6y9_0
    , output wire [0:0] oe_x6y9_0
    , input wire [0:0] ipin_x6y9_1
    , output wire [0:0] opin_x6y9_1
    , output wire [0:0] oe_x6y9_1
    , input wire [0:0] ipin_x7y9_0
    , output wire [0:0] opin_x7y9_0
    , output wire [0:0] oe_x7y9_0
    , input wire [0:0] ipin_x7y9_1
    , output wire [0:0] opin_x7y9_1
    , output wire [0:0] oe_x7y9_1
    , input wire [0:0] ipin_x8y9_0
    , output wire [0:0] opin_x8y9_0
    , output wire [0:0] oe_x8y9_0
    , input wire [0:0] ipin_x8y9_1
    , output wire [0:0] opin_x8y9_1
    , output wire [0:0] oe_x8y9_1
    , input wire [0:0] ipin_x9y1_0
    , output wire [0:0] opin_x9y1_0
    , output wire [0:0] oe_x9y1_0
    , input wire [0:0] ipin_x9y1_1
    , output wire [0:0] opin_x9y1_1
    , output wire [0:0] oe_x9y1_1
    , input wire [0:0] ipin_x9y2_0
    , output wire [0:0] opin_x9y2_0
    , output wire [0:0] oe_x9y2_0
    , input wire [0:0] ipin_x9y2_1
    , output wire [0:0] opin_x9y2_1
    , output wire [0:0] oe_x9y2_1
    , input wire [0:0] ipin_x9y3_0
    , output wire [0:0] opin_x9y3_0
    , output wire [0:0] oe_x9y3_0
    , input wire [0:0] ipin_x9y3_1
    , output wire [0:0] opin_x9y3_1
    , output wire [0:0] oe_x9y3_1
    , input wire [0:0] ipin_x9y4_0
    , output wire [0:0] opin_x9y4_0
    , output wire [0:0] oe_x9y4_0
    , input wire [0:0] ipin_x9y4_1
    , output wire [0:0] opin_x9y4_1
    , output wire [0:0] oe_x9y4_1
    , input wire [0:0] ipin_x9y5_0
    , output wire [0:0] opin_x9y5_0
    , output wire [0:0] oe_x9y5_0
    , input wire [0:0] ipin_x9y5_1
    , output wire [0:0] opin_x9y5_1
    , output wire [0:0] oe_x9y5_1
    , input wire [0:0] ipin_x9y6_0
    , output wire [0:0] opin_x9y6_0
    , output wire [0:0] oe_x9y6_0
    , input wire [0:0] ipin_x9y6_1
    , output wire [0:0] opin_x9y6_1
    , output wire [0:0] oe_x9y6_1
    , input wire [0:0] ipin_x9y7_0
    , output wire [0:0] opin_x9y7_0
    , output wire [0:0] oe_x9y7_0
    , input wire [0:0] ipin_x9y7_1
    , output wire [0:0] opin_x9y7_1
    , output wire [0:0] oe_x9y7_1
    , input wire [0:0] ipin_x9y8_0
    , output wire [0:0] opin_x9y8_0
    , output wire [0:0] oe_x9y8_0
    , input wire [0:0] ipin_x9y8_1
    , output wire [0:0] opin_x9y8_1
    , output wire [0:0] oe_x9y8_1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [11:0] _i_tile_x0y1__cu_x0y0n_L1;
    wire [11:0] _i_tile_x0y1__cu_x0y0s_L1;
    wire [0:0] _i_tile_x0y1__opin_x0y0_0;
    wire [0:0] _i_tile_x0y1__oe_x0y0_0;
    wire [0:0] _i_tile_x0y1__opin_x0y0_1;
    wire [0:0] _i_tile_x0y1__oe_x0y0_1;
    wire [0:0] _i_tile_x0y1__prog_dout;
    wire [0:0] _i_tile_x0y1__prog_we_o;
    wire [11:0] _i_sbox_x0y1ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x0y1ne__prog_dout;
    wire [0:0] _i_sbox_x0y1ne__prog_we_o;
    wire [11:0] _i_tile_x0y2__cu_x0y0n_L1;
    wire [11:0] _i_tile_x0y2__cu_x0y0s_L1;
    wire [0:0] _i_tile_x0y2__opin_x0y0_0;
    wire [0:0] _i_tile_x0y2__oe_x0y0_0;
    wire [0:0] _i_tile_x0y2__opin_x0y0_1;
    wire [0:0] _i_tile_x0y2__oe_x0y0_1;
    wire [0:0] _i_tile_x0y2__prog_dout;
    wire [0:0] _i_tile_x0y2__prog_we_o;
    wire [11:0] _i_sbox_x0y2ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x0y2ne__prog_dout;
    wire [0:0] _i_sbox_x0y2ne__prog_we_o;
    wire [11:0] _i_tile_x0y3__cu_x0y0n_L1;
    wire [11:0] _i_tile_x0y3__cu_x0y0s_L1;
    wire [0:0] _i_tile_x0y3__opin_x0y0_0;
    wire [0:0] _i_tile_x0y3__oe_x0y0_0;
    wire [0:0] _i_tile_x0y3__opin_x0y0_1;
    wire [0:0] _i_tile_x0y3__oe_x0y0_1;
    wire [0:0] _i_tile_x0y3__prog_dout;
    wire [0:0] _i_tile_x0y3__prog_we_o;
    wire [11:0] _i_sbox_x0y3ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x0y3ne__prog_dout;
    wire [0:0] _i_sbox_x0y3ne__prog_we_o;
    wire [11:0] _i_tile_x0y4__cu_x0y0n_L1;
    wire [11:0] _i_tile_x0y4__cu_x0y0s_L1;
    wire [0:0] _i_tile_x0y4__opin_x0y0_0;
    wire [0:0] _i_tile_x0y4__oe_x0y0_0;
    wire [0:0] _i_tile_x0y4__opin_x0y0_1;
    wire [0:0] _i_tile_x0y4__oe_x0y0_1;
    wire [0:0] _i_tile_x0y4__prog_dout;
    wire [0:0] _i_tile_x0y4__prog_we_o;
    wire [11:0] _i_sbox_x0y4ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x0y4ne__prog_dout;
    wire [0:0] _i_sbox_x0y4ne__prog_we_o;
    wire [11:0] _i_tile_x0y5__cu_x0y0n_L1;
    wire [11:0] _i_tile_x0y5__cu_x0y0s_L1;
    wire [0:0] _i_tile_x0y5__opin_x0y0_0;
    wire [0:0] _i_tile_x0y5__oe_x0y0_0;
    wire [0:0] _i_tile_x0y5__opin_x0y0_1;
    wire [0:0] _i_tile_x0y5__oe_x0y0_1;
    wire [0:0] _i_tile_x0y5__prog_dout;
    wire [0:0] _i_tile_x0y5__prog_we_o;
    wire [11:0] _i_sbox_x0y5ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x0y5ne__prog_dout;
    wire [0:0] _i_sbox_x0y5ne__prog_we_o;
    wire [11:0] _i_tile_x0y6__cu_x0y0n_L1;
    wire [11:0] _i_tile_x0y6__cu_x0y0s_L1;
    wire [0:0] _i_tile_x0y6__opin_x0y0_0;
    wire [0:0] _i_tile_x0y6__oe_x0y0_0;
    wire [0:0] _i_tile_x0y6__opin_x0y0_1;
    wire [0:0] _i_tile_x0y6__oe_x0y0_1;
    wire [0:0] _i_tile_x0y6__prog_dout;
    wire [0:0] _i_tile_x0y6__prog_we_o;
    wire [11:0] _i_sbox_x0y6ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x0y6ne__prog_dout;
    wire [0:0] _i_sbox_x0y6ne__prog_we_o;
    wire [11:0] _i_tile_x0y7__cu_x0y0n_L1;
    wire [11:0] _i_tile_x0y7__cu_x0y0s_L1;
    wire [0:0] _i_tile_x0y7__opin_x0y0_0;
    wire [0:0] _i_tile_x0y7__oe_x0y0_0;
    wire [0:0] _i_tile_x0y7__opin_x0y0_1;
    wire [0:0] _i_tile_x0y7__oe_x0y0_1;
    wire [0:0] _i_tile_x0y7__prog_dout;
    wire [0:0] _i_tile_x0y7__prog_we_o;
    wire [11:0] _i_sbox_x0y7ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x0y7ne__prog_dout;
    wire [0:0] _i_sbox_x0y7ne__prog_we_o;
    wire [11:0] _i_tile_x0y8__cu_x0y0n_L1;
    wire [11:0] _i_tile_x0y8__cu_x0y0s_L1;
    wire [0:0] _i_tile_x0y8__opin_x0y0_0;
    wire [0:0] _i_tile_x0y8__oe_x0y0_0;
    wire [0:0] _i_tile_x0y8__opin_x0y0_1;
    wire [0:0] _i_tile_x0y8__oe_x0y0_1;
    wire [0:0] _i_tile_x0y8__prog_dout;
    wire [0:0] _i_tile_x0y8__prog_we_o;
    wire [11:0] _i_sbox_x0y8ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x0y8ne__prog_dout;
    wire [0:0] _i_sbox_x0y8ne__prog_we_o;
    wire [11:0] _i_sbox_x1y0nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x1y0nw__prog_dout;
    wire [0:0] _i_sbox_x1y0nw__prog_we_o;
    wire [11:0] _i_tile_x1y1__cu_x0y0n_L1;
    wire [11:0] _i_tile_x1y1__cu_x0y0s_L1;
    wire [0:0] _i_tile_x1y1__prog_dout;
    wire [0:0] _i_tile_x1y1__prog_we_o;
    wire [11:0] _i_sbox_x1y1ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x1y1ne__prog_dout;
    wire [0:0] _i_sbox_x1y1ne__prog_we_o;
    wire [11:0] _i_sbox_x1y1nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x1y1nw__prog_dout;
    wire [0:0] _i_sbox_x1y1nw__prog_we_o;
    wire [11:0] _i_sbox_x1y1se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x1y1se__prog_dout;
    wire [0:0] _i_sbox_x1y1se__prog_we_o;
    wire [11:0] _i_sbox_x1y1sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x1y1sw__prog_dout;
    wire [0:0] _i_sbox_x1y1sw__prog_we_o;
    wire [11:0] _i_tile_x1y2__cu_x0y0n_L1;
    wire [11:0] _i_tile_x1y2__cu_x0y0s_L1;
    wire [0:0] _i_tile_x1y2__prog_dout;
    wire [0:0] _i_tile_x1y2__prog_we_o;
    wire [11:0] _i_sbox_x1y2ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x1y2ne__prog_dout;
    wire [0:0] _i_sbox_x1y2ne__prog_we_o;
    wire [11:0] _i_sbox_x1y2nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x1y2nw__prog_dout;
    wire [0:0] _i_sbox_x1y2nw__prog_we_o;
    wire [11:0] _i_sbox_x1y2se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x1y2se__prog_dout;
    wire [0:0] _i_sbox_x1y2se__prog_we_o;
    wire [11:0] _i_sbox_x1y2sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x1y2sw__prog_dout;
    wire [0:0] _i_sbox_x1y2sw__prog_we_o;
    wire [11:0] _i_tile_x1y3__cu_x0y0n_L1;
    wire [11:0] _i_tile_x1y3__cu_x0y0s_L1;
    wire [0:0] _i_tile_x1y3__prog_dout;
    wire [0:0] _i_tile_x1y3__prog_we_o;
    wire [11:0] _i_sbox_x1y3ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x1y3ne__prog_dout;
    wire [0:0] _i_sbox_x1y3ne__prog_we_o;
    wire [11:0] _i_sbox_x1y3nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x1y3nw__prog_dout;
    wire [0:0] _i_sbox_x1y3nw__prog_we_o;
    wire [11:0] _i_sbox_x1y3se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x1y3se__prog_dout;
    wire [0:0] _i_sbox_x1y3se__prog_we_o;
    wire [11:0] _i_sbox_x1y3sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x1y3sw__prog_dout;
    wire [0:0] _i_sbox_x1y3sw__prog_we_o;
    wire [11:0] _i_tile_x1y4__cu_x0y0n_L1;
    wire [11:0] _i_tile_x1y4__cu_x0y0s_L1;
    wire [0:0] _i_tile_x1y4__prog_dout;
    wire [0:0] _i_tile_x1y4__prog_we_o;
    wire [11:0] _i_sbox_x1y4ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x1y4ne__prog_dout;
    wire [0:0] _i_sbox_x1y4ne__prog_we_o;
    wire [11:0] _i_sbox_x1y4nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x1y4nw__prog_dout;
    wire [0:0] _i_sbox_x1y4nw__prog_we_o;
    wire [11:0] _i_sbox_x1y4se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x1y4se__prog_dout;
    wire [0:0] _i_sbox_x1y4se__prog_we_o;
    wire [11:0] _i_sbox_x1y4sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x1y4sw__prog_dout;
    wire [0:0] _i_sbox_x1y4sw__prog_we_o;
    wire [11:0] _i_tile_x1y5__cu_x0y0n_L1;
    wire [11:0] _i_tile_x1y5__cu_x0y0s_L1;
    wire [0:0] _i_tile_x1y5__prog_dout;
    wire [0:0] _i_tile_x1y5__prog_we_o;
    wire [11:0] _i_sbox_x1y5ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x1y5ne__prog_dout;
    wire [0:0] _i_sbox_x1y5ne__prog_we_o;
    wire [11:0] _i_sbox_x1y5nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x1y5nw__prog_dout;
    wire [0:0] _i_sbox_x1y5nw__prog_we_o;
    wire [11:0] _i_sbox_x1y5se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x1y5se__prog_dout;
    wire [0:0] _i_sbox_x1y5se__prog_we_o;
    wire [11:0] _i_sbox_x1y5sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x1y5sw__prog_dout;
    wire [0:0] _i_sbox_x1y5sw__prog_we_o;
    wire [11:0] _i_tile_x1y6__cu_x0y0n_L1;
    wire [11:0] _i_tile_x1y6__cu_x0y0s_L1;
    wire [0:0] _i_tile_x1y6__prog_dout;
    wire [0:0] _i_tile_x1y6__prog_we_o;
    wire [11:0] _i_sbox_x1y6ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x1y6ne__prog_dout;
    wire [0:0] _i_sbox_x1y6ne__prog_we_o;
    wire [11:0] _i_sbox_x1y6nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x1y6nw__prog_dout;
    wire [0:0] _i_sbox_x1y6nw__prog_we_o;
    wire [11:0] _i_sbox_x1y6se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x1y6se__prog_dout;
    wire [0:0] _i_sbox_x1y6se__prog_we_o;
    wire [11:0] _i_sbox_x1y6sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x1y6sw__prog_dout;
    wire [0:0] _i_sbox_x1y6sw__prog_we_o;
    wire [11:0] _i_tile_x1y7__cu_x0y0n_L1;
    wire [11:0] _i_tile_x1y7__cu_x0y0s_L1;
    wire [0:0] _i_tile_x1y7__prog_dout;
    wire [0:0] _i_tile_x1y7__prog_we_o;
    wire [11:0] _i_sbox_x1y7ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x1y7ne__prog_dout;
    wire [0:0] _i_sbox_x1y7ne__prog_we_o;
    wire [11:0] _i_sbox_x1y7nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x1y7nw__prog_dout;
    wire [0:0] _i_sbox_x1y7nw__prog_we_o;
    wire [11:0] _i_sbox_x1y7se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x1y7se__prog_dout;
    wire [0:0] _i_sbox_x1y7se__prog_we_o;
    wire [11:0] _i_sbox_x1y7sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x1y7sw__prog_dout;
    wire [0:0] _i_sbox_x1y7sw__prog_we_o;
    wire [11:0] _i_tile_x1y8__cu_x0y0n_L1;
    wire [11:0] _i_tile_x1y8__cu_x0y0s_L1;
    wire [0:0] _i_tile_x1y8__prog_dout;
    wire [0:0] _i_tile_x1y8__prog_we_o;
    wire [11:0] _i_sbox_x1y8ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x1y8ne__prog_dout;
    wire [0:0] _i_sbox_x1y8ne__prog_we_o;
    wire [11:0] _i_sbox_x1y8nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x1y8nw__prog_dout;
    wire [0:0] _i_sbox_x1y8nw__prog_we_o;
    wire [11:0] _i_sbox_x1y8se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x1y8se__prog_dout;
    wire [0:0] _i_sbox_x1y8se__prog_we_o;
    wire [11:0] _i_sbox_x1y8sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x1y8sw__prog_dout;
    wire [0:0] _i_sbox_x1y8sw__prog_we_o;
    wire [11:0] _i_tile_x1y9__cu_x0v1e_L1;
    wire [11:0] _i_tile_x1y9__cu_x0v1w_L1;
    wire [0:0] _i_tile_x1y9__opin_x0y0_0;
    wire [0:0] _i_tile_x1y9__oe_x0y0_0;
    wire [0:0] _i_tile_x1y9__opin_x0y0_1;
    wire [0:0] _i_tile_x1y9__oe_x0y0_1;
    wire [0:0] _i_tile_x1y9__prog_dout;
    wire [0:0] _i_tile_x1y9__prog_we_o;
    wire [11:0] _i_sbox_x1y9se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x1y9se__prog_dout;
    wire [0:0] _i_sbox_x1y9se__prog_we_o;
    wire [11:0] _i_sbox_x2y0nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x2y0nw__prog_dout;
    wire [0:0] _i_sbox_x2y0nw__prog_we_o;
    wire [11:0] _i_tile_x2y1__cu_x0y0n_L1;
    wire [11:0] _i_tile_x2y1__cu_x0y0s_L1;
    wire [0:0] _i_tile_x2y1__prog_dout;
    wire [0:0] _i_tile_x2y1__prog_we_o;
    wire [11:0] _i_sbox_x2y1ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x2y1ne__prog_dout;
    wire [0:0] _i_sbox_x2y1ne__prog_we_o;
    wire [11:0] _i_sbox_x2y1nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x2y1nw__prog_dout;
    wire [0:0] _i_sbox_x2y1nw__prog_we_o;
    wire [11:0] _i_sbox_x2y1se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x2y1se__prog_dout;
    wire [0:0] _i_sbox_x2y1se__prog_we_o;
    wire [11:0] _i_sbox_x2y1sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x2y1sw__prog_dout;
    wire [0:0] _i_sbox_x2y1sw__prog_we_o;
    wire [11:0] _i_tile_x2y2__cu_x0y0n_L1;
    wire [11:0] _i_tile_x2y2__cu_x0y0s_L1;
    wire [0:0] _i_tile_x2y2__prog_dout;
    wire [0:0] _i_tile_x2y2__prog_we_o;
    wire [11:0] _i_sbox_x2y2ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x2y2ne__prog_dout;
    wire [0:0] _i_sbox_x2y2ne__prog_we_o;
    wire [11:0] _i_sbox_x2y2nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x2y2nw__prog_dout;
    wire [0:0] _i_sbox_x2y2nw__prog_we_o;
    wire [11:0] _i_sbox_x2y2se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x2y2se__prog_dout;
    wire [0:0] _i_sbox_x2y2se__prog_we_o;
    wire [11:0] _i_sbox_x2y2sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x2y2sw__prog_dout;
    wire [0:0] _i_sbox_x2y2sw__prog_we_o;
    wire [11:0] _i_tile_x2y3__cu_x0y0n_L1;
    wire [11:0] _i_tile_x2y3__cu_x0y0s_L1;
    wire [0:0] _i_tile_x2y3__prog_dout;
    wire [0:0] _i_tile_x2y3__prog_we_o;
    wire [11:0] _i_sbox_x2y3ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x2y3ne__prog_dout;
    wire [0:0] _i_sbox_x2y3ne__prog_we_o;
    wire [11:0] _i_sbox_x2y3nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x2y3nw__prog_dout;
    wire [0:0] _i_sbox_x2y3nw__prog_we_o;
    wire [11:0] _i_sbox_x2y3se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x2y3se__prog_dout;
    wire [0:0] _i_sbox_x2y3se__prog_we_o;
    wire [11:0] _i_sbox_x2y3sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x2y3sw__prog_dout;
    wire [0:0] _i_sbox_x2y3sw__prog_we_o;
    wire [11:0] _i_tile_x2y4__cu_x0y0n_L1;
    wire [11:0] _i_tile_x2y4__cu_x0y0s_L1;
    wire [0:0] _i_tile_x2y4__prog_dout;
    wire [0:0] _i_tile_x2y4__prog_we_o;
    wire [11:0] _i_sbox_x2y4ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x2y4ne__prog_dout;
    wire [0:0] _i_sbox_x2y4ne__prog_we_o;
    wire [11:0] _i_sbox_x2y4nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x2y4nw__prog_dout;
    wire [0:0] _i_sbox_x2y4nw__prog_we_o;
    wire [11:0] _i_sbox_x2y4se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x2y4se__prog_dout;
    wire [0:0] _i_sbox_x2y4se__prog_we_o;
    wire [11:0] _i_sbox_x2y4sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x2y4sw__prog_dout;
    wire [0:0] _i_sbox_x2y4sw__prog_we_o;
    wire [11:0] _i_tile_x2y5__cu_x0y0n_L1;
    wire [11:0] _i_tile_x2y5__cu_x0y0s_L1;
    wire [0:0] _i_tile_x2y5__prog_dout;
    wire [0:0] _i_tile_x2y5__prog_we_o;
    wire [11:0] _i_sbox_x2y5ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x2y5ne__prog_dout;
    wire [0:0] _i_sbox_x2y5ne__prog_we_o;
    wire [11:0] _i_sbox_x2y5nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x2y5nw__prog_dout;
    wire [0:0] _i_sbox_x2y5nw__prog_we_o;
    wire [11:0] _i_sbox_x2y5se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x2y5se__prog_dout;
    wire [0:0] _i_sbox_x2y5se__prog_we_o;
    wire [11:0] _i_sbox_x2y5sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x2y5sw__prog_dout;
    wire [0:0] _i_sbox_x2y5sw__prog_we_o;
    wire [11:0] _i_tile_x2y6__cu_x0y0n_L1;
    wire [11:0] _i_tile_x2y6__cu_x0y0s_L1;
    wire [0:0] _i_tile_x2y6__prog_dout;
    wire [0:0] _i_tile_x2y6__prog_we_o;
    wire [11:0] _i_sbox_x2y6ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x2y6ne__prog_dout;
    wire [0:0] _i_sbox_x2y6ne__prog_we_o;
    wire [11:0] _i_sbox_x2y6nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x2y6nw__prog_dout;
    wire [0:0] _i_sbox_x2y6nw__prog_we_o;
    wire [11:0] _i_sbox_x2y6se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x2y6se__prog_dout;
    wire [0:0] _i_sbox_x2y6se__prog_we_o;
    wire [11:0] _i_sbox_x2y6sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x2y6sw__prog_dout;
    wire [0:0] _i_sbox_x2y6sw__prog_we_o;
    wire [11:0] _i_tile_x2y7__cu_x0y0n_L1;
    wire [11:0] _i_tile_x2y7__cu_x0y0s_L1;
    wire [0:0] _i_tile_x2y7__prog_dout;
    wire [0:0] _i_tile_x2y7__prog_we_o;
    wire [11:0] _i_sbox_x2y7ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x2y7ne__prog_dout;
    wire [0:0] _i_sbox_x2y7ne__prog_we_o;
    wire [11:0] _i_sbox_x2y7nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x2y7nw__prog_dout;
    wire [0:0] _i_sbox_x2y7nw__prog_we_o;
    wire [11:0] _i_sbox_x2y7se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x2y7se__prog_dout;
    wire [0:0] _i_sbox_x2y7se__prog_we_o;
    wire [11:0] _i_sbox_x2y7sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x2y7sw__prog_dout;
    wire [0:0] _i_sbox_x2y7sw__prog_we_o;
    wire [11:0] _i_tile_x2y8__cu_x0y0n_L1;
    wire [11:0] _i_tile_x2y8__cu_x0y0s_L1;
    wire [0:0] _i_tile_x2y8__prog_dout;
    wire [0:0] _i_tile_x2y8__prog_we_o;
    wire [11:0] _i_sbox_x2y8ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x2y8ne__prog_dout;
    wire [0:0] _i_sbox_x2y8ne__prog_we_o;
    wire [11:0] _i_sbox_x2y8nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x2y8nw__prog_dout;
    wire [0:0] _i_sbox_x2y8nw__prog_we_o;
    wire [11:0] _i_sbox_x2y8se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x2y8se__prog_dout;
    wire [0:0] _i_sbox_x2y8se__prog_we_o;
    wire [11:0] _i_sbox_x2y8sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x2y8sw__prog_dout;
    wire [0:0] _i_sbox_x2y8sw__prog_we_o;
    wire [11:0] _i_tile_x2y9__cu_x0v1e_L1;
    wire [11:0] _i_tile_x2y9__cu_x0v1w_L1;
    wire [0:0] _i_tile_x2y9__opin_x0y0_0;
    wire [0:0] _i_tile_x2y9__oe_x0y0_0;
    wire [0:0] _i_tile_x2y9__opin_x0y0_1;
    wire [0:0] _i_tile_x2y9__oe_x0y0_1;
    wire [0:0] _i_tile_x2y9__prog_dout;
    wire [0:0] _i_tile_x2y9__prog_we_o;
    wire [11:0] _i_sbox_x2y9se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x2y9se__prog_dout;
    wire [0:0] _i_sbox_x2y9se__prog_we_o;
    wire [11:0] _i_sbox_x3y0nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x3y0nw__prog_dout;
    wire [0:0] _i_sbox_x3y0nw__prog_we_o;
    wire [11:0] _i_tile_x3y1__cu_x0y0n_L1;
    wire [11:0] _i_tile_x3y1__cu_x0y0s_L1;
    wire [0:0] _i_tile_x3y1__prog_dout;
    wire [0:0] _i_tile_x3y1__prog_we_o;
    wire [11:0] _i_sbox_x3y1ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x3y1ne__prog_dout;
    wire [0:0] _i_sbox_x3y1ne__prog_we_o;
    wire [11:0] _i_sbox_x3y1nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x3y1nw__prog_dout;
    wire [0:0] _i_sbox_x3y1nw__prog_we_o;
    wire [11:0] _i_sbox_x3y1se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x3y1se__prog_dout;
    wire [0:0] _i_sbox_x3y1se__prog_we_o;
    wire [11:0] _i_sbox_x3y1sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x3y1sw__prog_dout;
    wire [0:0] _i_sbox_x3y1sw__prog_we_o;
    wire [11:0] _i_tile_x3y2__cu_x0y0n_L1;
    wire [11:0] _i_tile_x3y2__cu_x0y0s_L1;
    wire [0:0] _i_tile_x3y2__prog_dout;
    wire [0:0] _i_tile_x3y2__prog_we_o;
    wire [11:0] _i_sbox_x3y2ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x3y2ne__prog_dout;
    wire [0:0] _i_sbox_x3y2ne__prog_we_o;
    wire [11:0] _i_sbox_x3y2nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x3y2nw__prog_dout;
    wire [0:0] _i_sbox_x3y2nw__prog_we_o;
    wire [11:0] _i_sbox_x3y2se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x3y2se__prog_dout;
    wire [0:0] _i_sbox_x3y2se__prog_we_o;
    wire [11:0] _i_sbox_x3y2sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x3y2sw__prog_dout;
    wire [0:0] _i_sbox_x3y2sw__prog_we_o;
    wire [11:0] _i_tile_x3y3__cu_x0y0n_L1;
    wire [11:0] _i_tile_x3y3__cu_x0y0s_L1;
    wire [0:0] _i_tile_x3y3__prog_dout;
    wire [0:0] _i_tile_x3y3__prog_we_o;
    wire [11:0] _i_sbox_x3y3ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x3y3ne__prog_dout;
    wire [0:0] _i_sbox_x3y3ne__prog_we_o;
    wire [11:0] _i_sbox_x3y3nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x3y3nw__prog_dout;
    wire [0:0] _i_sbox_x3y3nw__prog_we_o;
    wire [11:0] _i_sbox_x3y3se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x3y3se__prog_dout;
    wire [0:0] _i_sbox_x3y3se__prog_we_o;
    wire [11:0] _i_sbox_x3y3sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x3y3sw__prog_dout;
    wire [0:0] _i_sbox_x3y3sw__prog_we_o;
    wire [11:0] _i_tile_x3y4__cu_x0y0n_L1;
    wire [11:0] _i_tile_x3y4__cu_x0y0s_L1;
    wire [0:0] _i_tile_x3y4__prog_dout;
    wire [0:0] _i_tile_x3y4__prog_we_o;
    wire [11:0] _i_sbox_x3y4ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x3y4ne__prog_dout;
    wire [0:0] _i_sbox_x3y4ne__prog_we_o;
    wire [11:0] _i_sbox_x3y4nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x3y4nw__prog_dout;
    wire [0:0] _i_sbox_x3y4nw__prog_we_o;
    wire [11:0] _i_sbox_x3y4se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x3y4se__prog_dout;
    wire [0:0] _i_sbox_x3y4se__prog_we_o;
    wire [11:0] _i_sbox_x3y4sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x3y4sw__prog_dout;
    wire [0:0] _i_sbox_x3y4sw__prog_we_o;
    wire [11:0] _i_tile_x3y5__cu_x0y0n_L1;
    wire [11:0] _i_tile_x3y5__cu_x0y0s_L1;
    wire [0:0] _i_tile_x3y5__prog_dout;
    wire [0:0] _i_tile_x3y5__prog_we_o;
    wire [11:0] _i_sbox_x3y5ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x3y5ne__prog_dout;
    wire [0:0] _i_sbox_x3y5ne__prog_we_o;
    wire [11:0] _i_sbox_x3y5nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x3y5nw__prog_dout;
    wire [0:0] _i_sbox_x3y5nw__prog_we_o;
    wire [11:0] _i_sbox_x3y5se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x3y5se__prog_dout;
    wire [0:0] _i_sbox_x3y5se__prog_we_o;
    wire [11:0] _i_sbox_x3y5sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x3y5sw__prog_dout;
    wire [0:0] _i_sbox_x3y5sw__prog_we_o;
    wire [11:0] _i_tile_x3y6__cu_x0y0n_L1;
    wire [11:0] _i_tile_x3y6__cu_x0y0s_L1;
    wire [0:0] _i_tile_x3y6__prog_dout;
    wire [0:0] _i_tile_x3y6__prog_we_o;
    wire [11:0] _i_sbox_x3y6ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x3y6ne__prog_dout;
    wire [0:0] _i_sbox_x3y6ne__prog_we_o;
    wire [11:0] _i_sbox_x3y6nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x3y6nw__prog_dout;
    wire [0:0] _i_sbox_x3y6nw__prog_we_o;
    wire [11:0] _i_sbox_x3y6se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x3y6se__prog_dout;
    wire [0:0] _i_sbox_x3y6se__prog_we_o;
    wire [11:0] _i_sbox_x3y6sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x3y6sw__prog_dout;
    wire [0:0] _i_sbox_x3y6sw__prog_we_o;
    wire [11:0] _i_tile_x3y7__cu_x0y0n_L1;
    wire [11:0] _i_tile_x3y7__cu_x0y0s_L1;
    wire [0:0] _i_tile_x3y7__prog_dout;
    wire [0:0] _i_tile_x3y7__prog_we_o;
    wire [11:0] _i_sbox_x3y7ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x3y7ne__prog_dout;
    wire [0:0] _i_sbox_x3y7ne__prog_we_o;
    wire [11:0] _i_sbox_x3y7nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x3y7nw__prog_dout;
    wire [0:0] _i_sbox_x3y7nw__prog_we_o;
    wire [11:0] _i_sbox_x3y7se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x3y7se__prog_dout;
    wire [0:0] _i_sbox_x3y7se__prog_we_o;
    wire [11:0] _i_sbox_x3y7sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x3y7sw__prog_dout;
    wire [0:0] _i_sbox_x3y7sw__prog_we_o;
    wire [11:0] _i_tile_x3y8__cu_x0y0n_L1;
    wire [11:0] _i_tile_x3y8__cu_x0y0s_L1;
    wire [0:0] _i_tile_x3y8__prog_dout;
    wire [0:0] _i_tile_x3y8__prog_we_o;
    wire [11:0] _i_sbox_x3y8ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x3y8ne__prog_dout;
    wire [0:0] _i_sbox_x3y8ne__prog_we_o;
    wire [11:0] _i_sbox_x3y8nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x3y8nw__prog_dout;
    wire [0:0] _i_sbox_x3y8nw__prog_we_o;
    wire [11:0] _i_sbox_x3y8se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x3y8se__prog_dout;
    wire [0:0] _i_sbox_x3y8se__prog_we_o;
    wire [11:0] _i_sbox_x3y8sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x3y8sw__prog_dout;
    wire [0:0] _i_sbox_x3y8sw__prog_we_o;
    wire [11:0] _i_tile_x3y9__cu_x0v1e_L1;
    wire [11:0] _i_tile_x3y9__cu_x0v1w_L1;
    wire [0:0] _i_tile_x3y9__opin_x0y0_0;
    wire [0:0] _i_tile_x3y9__oe_x0y0_0;
    wire [0:0] _i_tile_x3y9__opin_x0y0_1;
    wire [0:0] _i_tile_x3y9__oe_x0y0_1;
    wire [0:0] _i_tile_x3y9__prog_dout;
    wire [0:0] _i_tile_x3y9__prog_we_o;
    wire [11:0] _i_sbox_x3y9se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x3y9se__prog_dout;
    wire [0:0] _i_sbox_x3y9se__prog_we_o;
    wire [11:0] _i_sbox_x4y0nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x4y0nw__prog_dout;
    wire [0:0] _i_sbox_x4y0nw__prog_we_o;
    wire [11:0] _i_tile_x4y1__cu_x0y0n_L1;
    wire [11:0] _i_tile_x4y1__cu_x0y0s_L1;
    wire [0:0] _i_tile_x4y1__prog_dout;
    wire [0:0] _i_tile_x4y1__prog_we_o;
    wire [11:0] _i_sbox_x4y1ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x4y1ne__prog_dout;
    wire [0:0] _i_sbox_x4y1ne__prog_we_o;
    wire [11:0] _i_sbox_x4y1nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x4y1nw__prog_dout;
    wire [0:0] _i_sbox_x4y1nw__prog_we_o;
    wire [11:0] _i_sbox_x4y1se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x4y1se__prog_dout;
    wire [0:0] _i_sbox_x4y1se__prog_we_o;
    wire [11:0] _i_sbox_x4y1sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x4y1sw__prog_dout;
    wire [0:0] _i_sbox_x4y1sw__prog_we_o;
    wire [11:0] _i_tile_x4y2__cu_x0y0n_L1;
    wire [11:0] _i_tile_x4y2__cu_x0y0s_L1;
    wire [0:0] _i_tile_x4y2__prog_dout;
    wire [0:0] _i_tile_x4y2__prog_we_o;
    wire [11:0] _i_sbox_x4y2ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x4y2ne__prog_dout;
    wire [0:0] _i_sbox_x4y2ne__prog_we_o;
    wire [11:0] _i_sbox_x4y2nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x4y2nw__prog_dout;
    wire [0:0] _i_sbox_x4y2nw__prog_we_o;
    wire [11:0] _i_sbox_x4y2se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x4y2se__prog_dout;
    wire [0:0] _i_sbox_x4y2se__prog_we_o;
    wire [11:0] _i_sbox_x4y2sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x4y2sw__prog_dout;
    wire [0:0] _i_sbox_x4y2sw__prog_we_o;
    wire [11:0] _i_tile_x4y3__cu_x0y0n_L1;
    wire [11:0] _i_tile_x4y3__cu_x0y0s_L1;
    wire [0:0] _i_tile_x4y3__prog_dout;
    wire [0:0] _i_tile_x4y3__prog_we_o;
    wire [11:0] _i_sbox_x4y3ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x4y3ne__prog_dout;
    wire [0:0] _i_sbox_x4y3ne__prog_we_o;
    wire [11:0] _i_sbox_x4y3nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x4y3nw__prog_dout;
    wire [0:0] _i_sbox_x4y3nw__prog_we_o;
    wire [11:0] _i_sbox_x4y3se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x4y3se__prog_dout;
    wire [0:0] _i_sbox_x4y3se__prog_we_o;
    wire [11:0] _i_sbox_x4y3sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x4y3sw__prog_dout;
    wire [0:0] _i_sbox_x4y3sw__prog_we_o;
    wire [11:0] _i_tile_x4y4__cu_x0y0n_L1;
    wire [11:0] _i_tile_x4y4__cu_x0y0s_L1;
    wire [0:0] _i_tile_x4y4__prog_dout;
    wire [0:0] _i_tile_x4y4__prog_we_o;
    wire [11:0] _i_sbox_x4y4ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x4y4ne__prog_dout;
    wire [0:0] _i_sbox_x4y4ne__prog_we_o;
    wire [11:0] _i_sbox_x4y4nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x4y4nw__prog_dout;
    wire [0:0] _i_sbox_x4y4nw__prog_we_o;
    wire [11:0] _i_sbox_x4y4se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x4y4se__prog_dout;
    wire [0:0] _i_sbox_x4y4se__prog_we_o;
    wire [11:0] _i_sbox_x4y4sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x4y4sw__prog_dout;
    wire [0:0] _i_sbox_x4y4sw__prog_we_o;
    wire [11:0] _i_tile_x4y5__cu_x0y0n_L1;
    wire [11:0] _i_tile_x4y5__cu_x0y0s_L1;
    wire [0:0] _i_tile_x4y5__prog_dout;
    wire [0:0] _i_tile_x4y5__prog_we_o;
    wire [11:0] _i_sbox_x4y5ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x4y5ne__prog_dout;
    wire [0:0] _i_sbox_x4y5ne__prog_we_o;
    wire [11:0] _i_sbox_x4y5nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x4y5nw__prog_dout;
    wire [0:0] _i_sbox_x4y5nw__prog_we_o;
    wire [11:0] _i_sbox_x4y5se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x4y5se__prog_dout;
    wire [0:0] _i_sbox_x4y5se__prog_we_o;
    wire [11:0] _i_sbox_x4y5sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x4y5sw__prog_dout;
    wire [0:0] _i_sbox_x4y5sw__prog_we_o;
    wire [11:0] _i_tile_x4y6__cu_x0y0n_L1;
    wire [11:0] _i_tile_x4y6__cu_x0y0s_L1;
    wire [0:0] _i_tile_x4y6__prog_dout;
    wire [0:0] _i_tile_x4y6__prog_we_o;
    wire [11:0] _i_sbox_x4y6ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x4y6ne__prog_dout;
    wire [0:0] _i_sbox_x4y6ne__prog_we_o;
    wire [11:0] _i_sbox_x4y6nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x4y6nw__prog_dout;
    wire [0:0] _i_sbox_x4y6nw__prog_we_o;
    wire [11:0] _i_sbox_x4y6se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x4y6se__prog_dout;
    wire [0:0] _i_sbox_x4y6se__prog_we_o;
    wire [11:0] _i_sbox_x4y6sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x4y6sw__prog_dout;
    wire [0:0] _i_sbox_x4y6sw__prog_we_o;
    wire [11:0] _i_tile_x4y7__cu_x0y0n_L1;
    wire [11:0] _i_tile_x4y7__cu_x0y0s_L1;
    wire [0:0] _i_tile_x4y7__prog_dout;
    wire [0:0] _i_tile_x4y7__prog_we_o;
    wire [11:0] _i_sbox_x4y7ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x4y7ne__prog_dout;
    wire [0:0] _i_sbox_x4y7ne__prog_we_o;
    wire [11:0] _i_sbox_x4y7nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x4y7nw__prog_dout;
    wire [0:0] _i_sbox_x4y7nw__prog_we_o;
    wire [11:0] _i_sbox_x4y7se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x4y7se__prog_dout;
    wire [0:0] _i_sbox_x4y7se__prog_we_o;
    wire [11:0] _i_sbox_x4y7sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x4y7sw__prog_dout;
    wire [0:0] _i_sbox_x4y7sw__prog_we_o;
    wire [11:0] _i_tile_x4y8__cu_x0y0n_L1;
    wire [11:0] _i_tile_x4y8__cu_x0y0s_L1;
    wire [0:0] _i_tile_x4y8__prog_dout;
    wire [0:0] _i_tile_x4y8__prog_we_o;
    wire [11:0] _i_sbox_x4y8ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x4y8ne__prog_dout;
    wire [0:0] _i_sbox_x4y8ne__prog_we_o;
    wire [11:0] _i_sbox_x4y8nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x4y8nw__prog_dout;
    wire [0:0] _i_sbox_x4y8nw__prog_we_o;
    wire [11:0] _i_sbox_x4y8se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x4y8se__prog_dout;
    wire [0:0] _i_sbox_x4y8se__prog_we_o;
    wire [11:0] _i_sbox_x4y8sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x4y8sw__prog_dout;
    wire [0:0] _i_sbox_x4y8sw__prog_we_o;
    wire [11:0] _i_tile_x4y9__cu_x0v1e_L1;
    wire [11:0] _i_tile_x4y9__cu_x0v1w_L1;
    wire [0:0] _i_tile_x4y9__opin_x0y0_0;
    wire [0:0] _i_tile_x4y9__oe_x0y0_0;
    wire [0:0] _i_tile_x4y9__opin_x0y0_1;
    wire [0:0] _i_tile_x4y9__oe_x0y0_1;
    wire [0:0] _i_tile_x4y9__prog_dout;
    wire [0:0] _i_tile_x4y9__prog_we_o;
    wire [11:0] _i_sbox_x4y9se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x4y9se__prog_dout;
    wire [0:0] _i_sbox_x4y9se__prog_we_o;
    wire [11:0] _i_sbox_x5y0nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x5y0nw__prog_dout;
    wire [0:0] _i_sbox_x5y0nw__prog_we_o;
    wire [11:0] _i_tile_x5y1__cu_x0y0n_L1;
    wire [11:0] _i_tile_x5y1__cu_x0y0s_L1;
    wire [0:0] _i_tile_x5y1__prog_dout;
    wire [0:0] _i_tile_x5y1__prog_we_o;
    wire [11:0] _i_sbox_x5y1ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x5y1ne__prog_dout;
    wire [0:0] _i_sbox_x5y1ne__prog_we_o;
    wire [11:0] _i_sbox_x5y1nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x5y1nw__prog_dout;
    wire [0:0] _i_sbox_x5y1nw__prog_we_o;
    wire [11:0] _i_sbox_x5y1se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x5y1se__prog_dout;
    wire [0:0] _i_sbox_x5y1se__prog_we_o;
    wire [11:0] _i_sbox_x5y1sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x5y1sw__prog_dout;
    wire [0:0] _i_sbox_x5y1sw__prog_we_o;
    wire [11:0] _i_tile_x5y2__cu_x0y0n_L1;
    wire [11:0] _i_tile_x5y2__cu_x0y0s_L1;
    wire [0:0] _i_tile_x5y2__prog_dout;
    wire [0:0] _i_tile_x5y2__prog_we_o;
    wire [11:0] _i_sbox_x5y2ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x5y2ne__prog_dout;
    wire [0:0] _i_sbox_x5y2ne__prog_we_o;
    wire [11:0] _i_sbox_x5y2nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x5y2nw__prog_dout;
    wire [0:0] _i_sbox_x5y2nw__prog_we_o;
    wire [11:0] _i_sbox_x5y2se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x5y2se__prog_dout;
    wire [0:0] _i_sbox_x5y2se__prog_we_o;
    wire [11:0] _i_sbox_x5y2sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x5y2sw__prog_dout;
    wire [0:0] _i_sbox_x5y2sw__prog_we_o;
    wire [11:0] _i_tile_x5y3__cu_x0y0n_L1;
    wire [11:0] _i_tile_x5y3__cu_x0y0s_L1;
    wire [0:0] _i_tile_x5y3__prog_dout;
    wire [0:0] _i_tile_x5y3__prog_we_o;
    wire [11:0] _i_sbox_x5y3ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x5y3ne__prog_dout;
    wire [0:0] _i_sbox_x5y3ne__prog_we_o;
    wire [11:0] _i_sbox_x5y3nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x5y3nw__prog_dout;
    wire [0:0] _i_sbox_x5y3nw__prog_we_o;
    wire [11:0] _i_sbox_x5y3se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x5y3se__prog_dout;
    wire [0:0] _i_sbox_x5y3se__prog_we_o;
    wire [11:0] _i_sbox_x5y3sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x5y3sw__prog_dout;
    wire [0:0] _i_sbox_x5y3sw__prog_we_o;
    wire [11:0] _i_tile_x5y4__cu_x0y0n_L1;
    wire [11:0] _i_tile_x5y4__cu_x0y0s_L1;
    wire [0:0] _i_tile_x5y4__prog_dout;
    wire [0:0] _i_tile_x5y4__prog_we_o;
    wire [11:0] _i_sbox_x5y4ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x5y4ne__prog_dout;
    wire [0:0] _i_sbox_x5y4ne__prog_we_o;
    wire [11:0] _i_sbox_x5y4nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x5y4nw__prog_dout;
    wire [0:0] _i_sbox_x5y4nw__prog_we_o;
    wire [11:0] _i_sbox_x5y4se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x5y4se__prog_dout;
    wire [0:0] _i_sbox_x5y4se__prog_we_o;
    wire [11:0] _i_sbox_x5y4sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x5y4sw__prog_dout;
    wire [0:0] _i_sbox_x5y4sw__prog_we_o;
    wire [11:0] _i_tile_x5y5__cu_x0y0n_L1;
    wire [11:0] _i_tile_x5y5__cu_x0y0s_L1;
    wire [0:0] _i_tile_x5y5__prog_dout;
    wire [0:0] _i_tile_x5y5__prog_we_o;
    wire [11:0] _i_sbox_x5y5ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x5y5ne__prog_dout;
    wire [0:0] _i_sbox_x5y5ne__prog_we_o;
    wire [11:0] _i_sbox_x5y5nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x5y5nw__prog_dout;
    wire [0:0] _i_sbox_x5y5nw__prog_we_o;
    wire [11:0] _i_sbox_x5y5se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x5y5se__prog_dout;
    wire [0:0] _i_sbox_x5y5se__prog_we_o;
    wire [11:0] _i_sbox_x5y5sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x5y5sw__prog_dout;
    wire [0:0] _i_sbox_x5y5sw__prog_we_o;
    wire [11:0] _i_tile_x5y6__cu_x0y0n_L1;
    wire [11:0] _i_tile_x5y6__cu_x0y0s_L1;
    wire [0:0] _i_tile_x5y6__prog_dout;
    wire [0:0] _i_tile_x5y6__prog_we_o;
    wire [11:0] _i_sbox_x5y6ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x5y6ne__prog_dout;
    wire [0:0] _i_sbox_x5y6ne__prog_we_o;
    wire [11:0] _i_sbox_x5y6nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x5y6nw__prog_dout;
    wire [0:0] _i_sbox_x5y6nw__prog_we_o;
    wire [11:0] _i_sbox_x5y6se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x5y6se__prog_dout;
    wire [0:0] _i_sbox_x5y6se__prog_we_o;
    wire [11:0] _i_sbox_x5y6sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x5y6sw__prog_dout;
    wire [0:0] _i_sbox_x5y6sw__prog_we_o;
    wire [11:0] _i_tile_x5y7__cu_x0y0n_L1;
    wire [11:0] _i_tile_x5y7__cu_x0y0s_L1;
    wire [0:0] _i_tile_x5y7__prog_dout;
    wire [0:0] _i_tile_x5y7__prog_we_o;
    wire [11:0] _i_sbox_x5y7ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x5y7ne__prog_dout;
    wire [0:0] _i_sbox_x5y7ne__prog_we_o;
    wire [11:0] _i_sbox_x5y7nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x5y7nw__prog_dout;
    wire [0:0] _i_sbox_x5y7nw__prog_we_o;
    wire [11:0] _i_sbox_x5y7se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x5y7se__prog_dout;
    wire [0:0] _i_sbox_x5y7se__prog_we_o;
    wire [11:0] _i_sbox_x5y7sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x5y7sw__prog_dout;
    wire [0:0] _i_sbox_x5y7sw__prog_we_o;
    wire [11:0] _i_tile_x5y8__cu_x0y0n_L1;
    wire [11:0] _i_tile_x5y8__cu_x0y0s_L1;
    wire [0:0] _i_tile_x5y8__prog_dout;
    wire [0:0] _i_tile_x5y8__prog_we_o;
    wire [11:0] _i_sbox_x5y8ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x5y8ne__prog_dout;
    wire [0:0] _i_sbox_x5y8ne__prog_we_o;
    wire [11:0] _i_sbox_x5y8nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x5y8nw__prog_dout;
    wire [0:0] _i_sbox_x5y8nw__prog_we_o;
    wire [11:0] _i_sbox_x5y8se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x5y8se__prog_dout;
    wire [0:0] _i_sbox_x5y8se__prog_we_o;
    wire [11:0] _i_sbox_x5y8sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x5y8sw__prog_dout;
    wire [0:0] _i_sbox_x5y8sw__prog_we_o;
    wire [11:0] _i_tile_x5y9__cu_x0v1e_L1;
    wire [11:0] _i_tile_x5y9__cu_x0v1w_L1;
    wire [0:0] _i_tile_x5y9__opin_x0y0_0;
    wire [0:0] _i_tile_x5y9__oe_x0y0_0;
    wire [0:0] _i_tile_x5y9__opin_x0y0_1;
    wire [0:0] _i_tile_x5y9__oe_x0y0_1;
    wire [0:0] _i_tile_x5y9__prog_dout;
    wire [0:0] _i_tile_x5y9__prog_we_o;
    wire [11:0] _i_sbox_x5y9se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x5y9se__prog_dout;
    wire [0:0] _i_sbox_x5y9se__prog_we_o;
    wire [11:0] _i_sbox_x6y0nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x6y0nw__prog_dout;
    wire [0:0] _i_sbox_x6y0nw__prog_we_o;
    wire [11:0] _i_tile_x6y1__cu_x0y0n_L1;
    wire [11:0] _i_tile_x6y1__cu_x0y0s_L1;
    wire [0:0] _i_tile_x6y1__prog_dout;
    wire [0:0] _i_tile_x6y1__prog_we_o;
    wire [11:0] _i_sbox_x6y1ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x6y1ne__prog_dout;
    wire [0:0] _i_sbox_x6y1ne__prog_we_o;
    wire [11:0] _i_sbox_x6y1nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x6y1nw__prog_dout;
    wire [0:0] _i_sbox_x6y1nw__prog_we_o;
    wire [11:0] _i_sbox_x6y1se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x6y1se__prog_dout;
    wire [0:0] _i_sbox_x6y1se__prog_we_o;
    wire [11:0] _i_sbox_x6y1sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x6y1sw__prog_dout;
    wire [0:0] _i_sbox_x6y1sw__prog_we_o;
    wire [11:0] _i_tile_x6y2__cu_x0y0n_L1;
    wire [11:0] _i_tile_x6y2__cu_x0y0s_L1;
    wire [0:0] _i_tile_x6y2__prog_dout;
    wire [0:0] _i_tile_x6y2__prog_we_o;
    wire [11:0] _i_sbox_x6y2ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x6y2ne__prog_dout;
    wire [0:0] _i_sbox_x6y2ne__prog_we_o;
    wire [11:0] _i_sbox_x6y2nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x6y2nw__prog_dout;
    wire [0:0] _i_sbox_x6y2nw__prog_we_o;
    wire [11:0] _i_sbox_x6y2se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x6y2se__prog_dout;
    wire [0:0] _i_sbox_x6y2se__prog_we_o;
    wire [11:0] _i_sbox_x6y2sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x6y2sw__prog_dout;
    wire [0:0] _i_sbox_x6y2sw__prog_we_o;
    wire [11:0] _i_tile_x6y3__cu_x0y0n_L1;
    wire [11:0] _i_tile_x6y3__cu_x0y0s_L1;
    wire [0:0] _i_tile_x6y3__prog_dout;
    wire [0:0] _i_tile_x6y3__prog_we_o;
    wire [11:0] _i_sbox_x6y3ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x6y3ne__prog_dout;
    wire [0:0] _i_sbox_x6y3ne__prog_we_o;
    wire [11:0] _i_sbox_x6y3nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x6y3nw__prog_dout;
    wire [0:0] _i_sbox_x6y3nw__prog_we_o;
    wire [11:0] _i_sbox_x6y3se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x6y3se__prog_dout;
    wire [0:0] _i_sbox_x6y3se__prog_we_o;
    wire [11:0] _i_sbox_x6y3sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x6y3sw__prog_dout;
    wire [0:0] _i_sbox_x6y3sw__prog_we_o;
    wire [11:0] _i_tile_x6y4__cu_x0y0n_L1;
    wire [11:0] _i_tile_x6y4__cu_x0y0s_L1;
    wire [0:0] _i_tile_x6y4__prog_dout;
    wire [0:0] _i_tile_x6y4__prog_we_o;
    wire [11:0] _i_sbox_x6y4ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x6y4ne__prog_dout;
    wire [0:0] _i_sbox_x6y4ne__prog_we_o;
    wire [11:0] _i_sbox_x6y4nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x6y4nw__prog_dout;
    wire [0:0] _i_sbox_x6y4nw__prog_we_o;
    wire [11:0] _i_sbox_x6y4se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x6y4se__prog_dout;
    wire [0:0] _i_sbox_x6y4se__prog_we_o;
    wire [11:0] _i_sbox_x6y4sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x6y4sw__prog_dout;
    wire [0:0] _i_sbox_x6y4sw__prog_we_o;
    wire [11:0] _i_tile_x6y5__cu_x0y0n_L1;
    wire [11:0] _i_tile_x6y5__cu_x0y0s_L1;
    wire [0:0] _i_tile_x6y5__prog_dout;
    wire [0:0] _i_tile_x6y5__prog_we_o;
    wire [11:0] _i_sbox_x6y5ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x6y5ne__prog_dout;
    wire [0:0] _i_sbox_x6y5ne__prog_we_o;
    wire [11:0] _i_sbox_x6y5nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x6y5nw__prog_dout;
    wire [0:0] _i_sbox_x6y5nw__prog_we_o;
    wire [11:0] _i_sbox_x6y5se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x6y5se__prog_dout;
    wire [0:0] _i_sbox_x6y5se__prog_we_o;
    wire [11:0] _i_sbox_x6y5sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x6y5sw__prog_dout;
    wire [0:0] _i_sbox_x6y5sw__prog_we_o;
    wire [11:0] _i_tile_x6y6__cu_x0y0n_L1;
    wire [11:0] _i_tile_x6y6__cu_x0y0s_L1;
    wire [0:0] _i_tile_x6y6__prog_dout;
    wire [0:0] _i_tile_x6y6__prog_we_o;
    wire [11:0] _i_sbox_x6y6ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x6y6ne__prog_dout;
    wire [0:0] _i_sbox_x6y6ne__prog_we_o;
    wire [11:0] _i_sbox_x6y6nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x6y6nw__prog_dout;
    wire [0:0] _i_sbox_x6y6nw__prog_we_o;
    wire [11:0] _i_sbox_x6y6se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x6y6se__prog_dout;
    wire [0:0] _i_sbox_x6y6se__prog_we_o;
    wire [11:0] _i_sbox_x6y6sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x6y6sw__prog_dout;
    wire [0:0] _i_sbox_x6y6sw__prog_we_o;
    wire [11:0] _i_tile_x6y7__cu_x0y0n_L1;
    wire [11:0] _i_tile_x6y7__cu_x0y0s_L1;
    wire [0:0] _i_tile_x6y7__prog_dout;
    wire [0:0] _i_tile_x6y7__prog_we_o;
    wire [11:0] _i_sbox_x6y7ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x6y7ne__prog_dout;
    wire [0:0] _i_sbox_x6y7ne__prog_we_o;
    wire [11:0] _i_sbox_x6y7nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x6y7nw__prog_dout;
    wire [0:0] _i_sbox_x6y7nw__prog_we_o;
    wire [11:0] _i_sbox_x6y7se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x6y7se__prog_dout;
    wire [0:0] _i_sbox_x6y7se__prog_we_o;
    wire [11:0] _i_sbox_x6y7sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x6y7sw__prog_dout;
    wire [0:0] _i_sbox_x6y7sw__prog_we_o;
    wire [11:0] _i_tile_x6y8__cu_x0y0n_L1;
    wire [11:0] _i_tile_x6y8__cu_x0y0s_L1;
    wire [0:0] _i_tile_x6y8__prog_dout;
    wire [0:0] _i_tile_x6y8__prog_we_o;
    wire [11:0] _i_sbox_x6y8ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x6y8ne__prog_dout;
    wire [0:0] _i_sbox_x6y8ne__prog_we_o;
    wire [11:0] _i_sbox_x6y8nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x6y8nw__prog_dout;
    wire [0:0] _i_sbox_x6y8nw__prog_we_o;
    wire [11:0] _i_sbox_x6y8se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x6y8se__prog_dout;
    wire [0:0] _i_sbox_x6y8se__prog_we_o;
    wire [11:0] _i_sbox_x6y8sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x6y8sw__prog_dout;
    wire [0:0] _i_sbox_x6y8sw__prog_we_o;
    wire [11:0] _i_tile_x6y9__cu_x0v1e_L1;
    wire [11:0] _i_tile_x6y9__cu_x0v1w_L1;
    wire [0:0] _i_tile_x6y9__opin_x0y0_0;
    wire [0:0] _i_tile_x6y9__oe_x0y0_0;
    wire [0:0] _i_tile_x6y9__opin_x0y0_1;
    wire [0:0] _i_tile_x6y9__oe_x0y0_1;
    wire [0:0] _i_tile_x6y9__prog_dout;
    wire [0:0] _i_tile_x6y9__prog_we_o;
    wire [11:0] _i_sbox_x6y9se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x6y9se__prog_dout;
    wire [0:0] _i_sbox_x6y9se__prog_we_o;
    wire [11:0] _i_sbox_x7y0nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x7y0nw__prog_dout;
    wire [0:0] _i_sbox_x7y0nw__prog_we_o;
    wire [11:0] _i_tile_x7y1__cu_x0y0n_L1;
    wire [11:0] _i_tile_x7y1__cu_x0y0s_L1;
    wire [0:0] _i_tile_x7y1__prog_dout;
    wire [0:0] _i_tile_x7y1__prog_we_o;
    wire [11:0] _i_sbox_x7y1ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x7y1ne__prog_dout;
    wire [0:0] _i_sbox_x7y1ne__prog_we_o;
    wire [11:0] _i_sbox_x7y1nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x7y1nw__prog_dout;
    wire [0:0] _i_sbox_x7y1nw__prog_we_o;
    wire [11:0] _i_sbox_x7y1se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x7y1se__prog_dout;
    wire [0:0] _i_sbox_x7y1se__prog_we_o;
    wire [11:0] _i_sbox_x7y1sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x7y1sw__prog_dout;
    wire [0:0] _i_sbox_x7y1sw__prog_we_o;
    wire [11:0] _i_tile_x7y2__cu_x0y0n_L1;
    wire [11:0] _i_tile_x7y2__cu_x0y0s_L1;
    wire [0:0] _i_tile_x7y2__prog_dout;
    wire [0:0] _i_tile_x7y2__prog_we_o;
    wire [11:0] _i_sbox_x7y2ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x7y2ne__prog_dout;
    wire [0:0] _i_sbox_x7y2ne__prog_we_o;
    wire [11:0] _i_sbox_x7y2nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x7y2nw__prog_dout;
    wire [0:0] _i_sbox_x7y2nw__prog_we_o;
    wire [11:0] _i_sbox_x7y2se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x7y2se__prog_dout;
    wire [0:0] _i_sbox_x7y2se__prog_we_o;
    wire [11:0] _i_sbox_x7y2sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x7y2sw__prog_dout;
    wire [0:0] _i_sbox_x7y2sw__prog_we_o;
    wire [11:0] _i_tile_x7y3__cu_x0y0n_L1;
    wire [11:0] _i_tile_x7y3__cu_x0y0s_L1;
    wire [0:0] _i_tile_x7y3__prog_dout;
    wire [0:0] _i_tile_x7y3__prog_we_o;
    wire [11:0] _i_sbox_x7y3ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x7y3ne__prog_dout;
    wire [0:0] _i_sbox_x7y3ne__prog_we_o;
    wire [11:0] _i_sbox_x7y3nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x7y3nw__prog_dout;
    wire [0:0] _i_sbox_x7y3nw__prog_we_o;
    wire [11:0] _i_sbox_x7y3se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x7y3se__prog_dout;
    wire [0:0] _i_sbox_x7y3se__prog_we_o;
    wire [11:0] _i_sbox_x7y3sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x7y3sw__prog_dout;
    wire [0:0] _i_sbox_x7y3sw__prog_we_o;
    wire [11:0] _i_tile_x7y4__cu_x0y0n_L1;
    wire [11:0] _i_tile_x7y4__cu_x0y0s_L1;
    wire [0:0] _i_tile_x7y4__prog_dout;
    wire [0:0] _i_tile_x7y4__prog_we_o;
    wire [11:0] _i_sbox_x7y4ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x7y4ne__prog_dout;
    wire [0:0] _i_sbox_x7y4ne__prog_we_o;
    wire [11:0] _i_sbox_x7y4nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x7y4nw__prog_dout;
    wire [0:0] _i_sbox_x7y4nw__prog_we_o;
    wire [11:0] _i_sbox_x7y4se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x7y4se__prog_dout;
    wire [0:0] _i_sbox_x7y4se__prog_we_o;
    wire [11:0] _i_sbox_x7y4sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x7y4sw__prog_dout;
    wire [0:0] _i_sbox_x7y4sw__prog_we_o;
    wire [11:0] _i_tile_x7y5__cu_x0y0n_L1;
    wire [11:0] _i_tile_x7y5__cu_x0y0s_L1;
    wire [0:0] _i_tile_x7y5__prog_dout;
    wire [0:0] _i_tile_x7y5__prog_we_o;
    wire [11:0] _i_sbox_x7y5ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x7y5ne__prog_dout;
    wire [0:0] _i_sbox_x7y5ne__prog_we_o;
    wire [11:0] _i_sbox_x7y5nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x7y5nw__prog_dout;
    wire [0:0] _i_sbox_x7y5nw__prog_we_o;
    wire [11:0] _i_sbox_x7y5se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x7y5se__prog_dout;
    wire [0:0] _i_sbox_x7y5se__prog_we_o;
    wire [11:0] _i_sbox_x7y5sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x7y5sw__prog_dout;
    wire [0:0] _i_sbox_x7y5sw__prog_we_o;
    wire [11:0] _i_tile_x7y6__cu_x0y0n_L1;
    wire [11:0] _i_tile_x7y6__cu_x0y0s_L1;
    wire [0:0] _i_tile_x7y6__prog_dout;
    wire [0:0] _i_tile_x7y6__prog_we_o;
    wire [11:0] _i_sbox_x7y6ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x7y6ne__prog_dout;
    wire [0:0] _i_sbox_x7y6ne__prog_we_o;
    wire [11:0] _i_sbox_x7y6nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x7y6nw__prog_dout;
    wire [0:0] _i_sbox_x7y6nw__prog_we_o;
    wire [11:0] _i_sbox_x7y6se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x7y6se__prog_dout;
    wire [0:0] _i_sbox_x7y6se__prog_we_o;
    wire [11:0] _i_sbox_x7y6sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x7y6sw__prog_dout;
    wire [0:0] _i_sbox_x7y6sw__prog_we_o;
    wire [11:0] _i_tile_x7y7__cu_x0y0n_L1;
    wire [11:0] _i_tile_x7y7__cu_x0y0s_L1;
    wire [0:0] _i_tile_x7y7__prog_dout;
    wire [0:0] _i_tile_x7y7__prog_we_o;
    wire [11:0] _i_sbox_x7y7ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x7y7ne__prog_dout;
    wire [0:0] _i_sbox_x7y7ne__prog_we_o;
    wire [11:0] _i_sbox_x7y7nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x7y7nw__prog_dout;
    wire [0:0] _i_sbox_x7y7nw__prog_we_o;
    wire [11:0] _i_sbox_x7y7se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x7y7se__prog_dout;
    wire [0:0] _i_sbox_x7y7se__prog_we_o;
    wire [11:0] _i_sbox_x7y7sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x7y7sw__prog_dout;
    wire [0:0] _i_sbox_x7y7sw__prog_we_o;
    wire [11:0] _i_tile_x7y8__cu_x0y0n_L1;
    wire [11:0] _i_tile_x7y8__cu_x0y0s_L1;
    wire [0:0] _i_tile_x7y8__prog_dout;
    wire [0:0] _i_tile_x7y8__prog_we_o;
    wire [11:0] _i_sbox_x7y8ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x7y8ne__prog_dout;
    wire [0:0] _i_sbox_x7y8ne__prog_we_o;
    wire [11:0] _i_sbox_x7y8nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x7y8nw__prog_dout;
    wire [0:0] _i_sbox_x7y8nw__prog_we_o;
    wire [11:0] _i_sbox_x7y8se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x7y8se__prog_dout;
    wire [0:0] _i_sbox_x7y8se__prog_we_o;
    wire [11:0] _i_sbox_x7y8sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x7y8sw__prog_dout;
    wire [0:0] _i_sbox_x7y8sw__prog_we_o;
    wire [11:0] _i_tile_x7y9__cu_x0v1e_L1;
    wire [11:0] _i_tile_x7y9__cu_x0v1w_L1;
    wire [0:0] _i_tile_x7y9__opin_x0y0_0;
    wire [0:0] _i_tile_x7y9__oe_x0y0_0;
    wire [0:0] _i_tile_x7y9__opin_x0y0_1;
    wire [0:0] _i_tile_x7y9__oe_x0y0_1;
    wire [0:0] _i_tile_x7y9__prog_dout;
    wire [0:0] _i_tile_x7y9__prog_we_o;
    wire [11:0] _i_sbox_x7y9se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x7y9se__prog_dout;
    wire [0:0] _i_sbox_x7y9se__prog_we_o;
    wire [11:0] _i_sbox_x8y0nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x8y0nw__prog_dout;
    wire [0:0] _i_sbox_x8y0nw__prog_we_o;
    wire [11:0] _i_tile_x8y1__cu_x0y0n_L1;
    wire [11:0] _i_tile_x8y1__cu_x0y0s_L1;
    wire [0:0] _i_tile_x8y1__prog_dout;
    wire [0:0] _i_tile_x8y1__prog_we_o;
    wire [11:0] _i_sbox_x8y1ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x8y1ne__prog_dout;
    wire [0:0] _i_sbox_x8y1ne__prog_we_o;
    wire [11:0] _i_sbox_x8y1nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x8y1nw__prog_dout;
    wire [0:0] _i_sbox_x8y1nw__prog_we_o;
    wire [11:0] _i_sbox_x8y1se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x8y1se__prog_dout;
    wire [0:0] _i_sbox_x8y1se__prog_we_o;
    wire [11:0] _i_sbox_x8y1sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x8y1sw__prog_dout;
    wire [0:0] _i_sbox_x8y1sw__prog_we_o;
    wire [11:0] _i_tile_x8y2__cu_x0y0n_L1;
    wire [11:0] _i_tile_x8y2__cu_x0y0s_L1;
    wire [0:0] _i_tile_x8y2__prog_dout;
    wire [0:0] _i_tile_x8y2__prog_we_o;
    wire [11:0] _i_sbox_x8y2ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x8y2ne__prog_dout;
    wire [0:0] _i_sbox_x8y2ne__prog_we_o;
    wire [11:0] _i_sbox_x8y2nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x8y2nw__prog_dout;
    wire [0:0] _i_sbox_x8y2nw__prog_we_o;
    wire [11:0] _i_sbox_x8y2se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x8y2se__prog_dout;
    wire [0:0] _i_sbox_x8y2se__prog_we_o;
    wire [11:0] _i_sbox_x8y2sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x8y2sw__prog_dout;
    wire [0:0] _i_sbox_x8y2sw__prog_we_o;
    wire [11:0] _i_tile_x8y3__cu_x0y0n_L1;
    wire [11:0] _i_tile_x8y3__cu_x0y0s_L1;
    wire [0:0] _i_tile_x8y3__prog_dout;
    wire [0:0] _i_tile_x8y3__prog_we_o;
    wire [11:0] _i_sbox_x8y3ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x8y3ne__prog_dout;
    wire [0:0] _i_sbox_x8y3ne__prog_we_o;
    wire [11:0] _i_sbox_x8y3nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x8y3nw__prog_dout;
    wire [0:0] _i_sbox_x8y3nw__prog_we_o;
    wire [11:0] _i_sbox_x8y3se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x8y3se__prog_dout;
    wire [0:0] _i_sbox_x8y3se__prog_we_o;
    wire [11:0] _i_sbox_x8y3sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x8y3sw__prog_dout;
    wire [0:0] _i_sbox_x8y3sw__prog_we_o;
    wire [11:0] _i_tile_x8y4__cu_x0y0n_L1;
    wire [11:0] _i_tile_x8y4__cu_x0y0s_L1;
    wire [0:0] _i_tile_x8y4__prog_dout;
    wire [0:0] _i_tile_x8y4__prog_we_o;
    wire [11:0] _i_sbox_x8y4ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x8y4ne__prog_dout;
    wire [0:0] _i_sbox_x8y4ne__prog_we_o;
    wire [11:0] _i_sbox_x8y4nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x8y4nw__prog_dout;
    wire [0:0] _i_sbox_x8y4nw__prog_we_o;
    wire [11:0] _i_sbox_x8y4se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x8y4se__prog_dout;
    wire [0:0] _i_sbox_x8y4se__prog_we_o;
    wire [11:0] _i_sbox_x8y4sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x8y4sw__prog_dout;
    wire [0:0] _i_sbox_x8y4sw__prog_we_o;
    wire [11:0] _i_tile_x8y5__cu_x0y0n_L1;
    wire [11:0] _i_tile_x8y5__cu_x0y0s_L1;
    wire [0:0] _i_tile_x8y5__prog_dout;
    wire [0:0] _i_tile_x8y5__prog_we_o;
    wire [11:0] _i_sbox_x8y5ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x8y5ne__prog_dout;
    wire [0:0] _i_sbox_x8y5ne__prog_we_o;
    wire [11:0] _i_sbox_x8y5nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x8y5nw__prog_dout;
    wire [0:0] _i_sbox_x8y5nw__prog_we_o;
    wire [11:0] _i_sbox_x8y5se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x8y5se__prog_dout;
    wire [0:0] _i_sbox_x8y5se__prog_we_o;
    wire [11:0] _i_sbox_x8y5sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x8y5sw__prog_dout;
    wire [0:0] _i_sbox_x8y5sw__prog_we_o;
    wire [11:0] _i_tile_x8y6__cu_x0y0n_L1;
    wire [11:0] _i_tile_x8y6__cu_x0y0s_L1;
    wire [0:0] _i_tile_x8y6__prog_dout;
    wire [0:0] _i_tile_x8y6__prog_we_o;
    wire [11:0] _i_sbox_x8y6ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x8y6ne__prog_dout;
    wire [0:0] _i_sbox_x8y6ne__prog_we_o;
    wire [11:0] _i_sbox_x8y6nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x8y6nw__prog_dout;
    wire [0:0] _i_sbox_x8y6nw__prog_we_o;
    wire [11:0] _i_sbox_x8y6se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x8y6se__prog_dout;
    wire [0:0] _i_sbox_x8y6se__prog_we_o;
    wire [11:0] _i_sbox_x8y6sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x8y6sw__prog_dout;
    wire [0:0] _i_sbox_x8y6sw__prog_we_o;
    wire [11:0] _i_tile_x8y7__cu_x0y0n_L1;
    wire [11:0] _i_tile_x8y7__cu_x0y0s_L1;
    wire [0:0] _i_tile_x8y7__prog_dout;
    wire [0:0] _i_tile_x8y7__prog_we_o;
    wire [11:0] _i_sbox_x8y7ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x8y7ne__prog_dout;
    wire [0:0] _i_sbox_x8y7ne__prog_we_o;
    wire [11:0] _i_sbox_x8y7nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x8y7nw__prog_dout;
    wire [0:0] _i_sbox_x8y7nw__prog_we_o;
    wire [11:0] _i_sbox_x8y7se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x8y7se__prog_dout;
    wire [0:0] _i_sbox_x8y7se__prog_we_o;
    wire [11:0] _i_sbox_x8y7sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x8y7sw__prog_dout;
    wire [0:0] _i_sbox_x8y7sw__prog_we_o;
    wire [11:0] _i_tile_x8y8__cu_x0y0n_L1;
    wire [11:0] _i_tile_x8y8__cu_x0y0s_L1;
    wire [0:0] _i_tile_x8y8__prog_dout;
    wire [0:0] _i_tile_x8y8__prog_we_o;
    wire [11:0] _i_sbox_x8y8ne__so_x0y0s_L1;
    wire [0:0] _i_sbox_x8y8ne__prog_dout;
    wire [0:0] _i_sbox_x8y8ne__prog_we_o;
    wire [11:0] _i_sbox_x8y8nw__so_x0y0e_L1;
    wire [0:0] _i_sbox_x8y8nw__prog_dout;
    wire [0:0] _i_sbox_x8y8nw__prog_we_o;
    wire [11:0] _i_sbox_x8y8se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x8y8se__prog_dout;
    wire [0:0] _i_sbox_x8y8se__prog_we_o;
    wire [11:0] _i_sbox_x8y8sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x8y8sw__prog_dout;
    wire [0:0] _i_sbox_x8y8sw__prog_we_o;
    wire [11:0] _i_tile_x8y9__cu_x0v1e_L1;
    wire [11:0] _i_tile_x8y9__cu_x0v1w_L1;
    wire [0:0] _i_tile_x8y9__opin_x0y0_0;
    wire [0:0] _i_tile_x8y9__oe_x0y0_0;
    wire [0:0] _i_tile_x8y9__opin_x0y0_1;
    wire [0:0] _i_tile_x8y9__oe_x0y0_1;
    wire [0:0] _i_tile_x8y9__prog_dout;
    wire [0:0] _i_tile_x8y9__prog_we_o;
    wire [11:0] _i_sbox_x8y9se__so_x0v1w_L1;
    wire [0:0] _i_sbox_x8y9se__prog_dout;
    wire [0:0] _i_sbox_x8y9se__prog_we_o;
    wire [11:0] _i_tile_x9y1__cu_u1y0n_L1;
    wire [11:0] _i_tile_x9y1__cu_u1y0s_L1;
    wire [0:0] _i_tile_x9y1__opin_x0y0_0;
    wire [0:0] _i_tile_x9y1__oe_x0y0_0;
    wire [0:0] _i_tile_x9y1__opin_x0y0_1;
    wire [0:0] _i_tile_x9y1__oe_x0y0_1;
    wire [0:0] _i_tile_x9y1__prog_dout;
    wire [0:0] _i_tile_x9y1__prog_we_o;
    wire [11:0] _i_sbox_x9y1sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x9y1sw__prog_dout;
    wire [0:0] _i_sbox_x9y1sw__prog_we_o;
    wire [11:0] _i_tile_x9y2__cu_u1y0n_L1;
    wire [11:0] _i_tile_x9y2__cu_u1y0s_L1;
    wire [0:0] _i_tile_x9y2__opin_x0y0_0;
    wire [0:0] _i_tile_x9y2__oe_x0y0_0;
    wire [0:0] _i_tile_x9y2__opin_x0y0_1;
    wire [0:0] _i_tile_x9y2__oe_x0y0_1;
    wire [0:0] _i_tile_x9y2__prog_dout;
    wire [0:0] _i_tile_x9y2__prog_we_o;
    wire [11:0] _i_sbox_x9y2sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x9y2sw__prog_dout;
    wire [0:0] _i_sbox_x9y2sw__prog_we_o;
    wire [11:0] _i_tile_x9y3__cu_u1y0n_L1;
    wire [11:0] _i_tile_x9y3__cu_u1y0s_L1;
    wire [0:0] _i_tile_x9y3__opin_x0y0_0;
    wire [0:0] _i_tile_x9y3__oe_x0y0_0;
    wire [0:0] _i_tile_x9y3__opin_x0y0_1;
    wire [0:0] _i_tile_x9y3__oe_x0y0_1;
    wire [0:0] _i_tile_x9y3__prog_dout;
    wire [0:0] _i_tile_x9y3__prog_we_o;
    wire [11:0] _i_sbox_x9y3sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x9y3sw__prog_dout;
    wire [0:0] _i_sbox_x9y3sw__prog_we_o;
    wire [11:0] _i_tile_x9y4__cu_u1y0n_L1;
    wire [11:0] _i_tile_x9y4__cu_u1y0s_L1;
    wire [0:0] _i_tile_x9y4__opin_x0y0_0;
    wire [0:0] _i_tile_x9y4__oe_x0y0_0;
    wire [0:0] _i_tile_x9y4__opin_x0y0_1;
    wire [0:0] _i_tile_x9y4__oe_x0y0_1;
    wire [0:0] _i_tile_x9y4__prog_dout;
    wire [0:0] _i_tile_x9y4__prog_we_o;
    wire [11:0] _i_sbox_x9y4sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x9y4sw__prog_dout;
    wire [0:0] _i_sbox_x9y4sw__prog_we_o;
    wire [11:0] _i_tile_x9y5__cu_u1y0n_L1;
    wire [11:0] _i_tile_x9y5__cu_u1y0s_L1;
    wire [0:0] _i_tile_x9y5__opin_x0y0_0;
    wire [0:0] _i_tile_x9y5__oe_x0y0_0;
    wire [0:0] _i_tile_x9y5__opin_x0y0_1;
    wire [0:0] _i_tile_x9y5__oe_x0y0_1;
    wire [0:0] _i_tile_x9y5__prog_dout;
    wire [0:0] _i_tile_x9y5__prog_we_o;
    wire [11:0] _i_sbox_x9y5sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x9y5sw__prog_dout;
    wire [0:0] _i_sbox_x9y5sw__prog_we_o;
    wire [11:0] _i_tile_x9y6__cu_u1y0n_L1;
    wire [11:0] _i_tile_x9y6__cu_u1y0s_L1;
    wire [0:0] _i_tile_x9y6__opin_x0y0_0;
    wire [0:0] _i_tile_x9y6__oe_x0y0_0;
    wire [0:0] _i_tile_x9y6__opin_x0y0_1;
    wire [0:0] _i_tile_x9y6__oe_x0y0_1;
    wire [0:0] _i_tile_x9y6__prog_dout;
    wire [0:0] _i_tile_x9y6__prog_we_o;
    wire [11:0] _i_sbox_x9y6sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x9y6sw__prog_dout;
    wire [0:0] _i_sbox_x9y6sw__prog_we_o;
    wire [11:0] _i_tile_x9y7__cu_u1y0n_L1;
    wire [11:0] _i_tile_x9y7__cu_u1y0s_L1;
    wire [0:0] _i_tile_x9y7__opin_x0y0_0;
    wire [0:0] _i_tile_x9y7__oe_x0y0_0;
    wire [0:0] _i_tile_x9y7__opin_x0y0_1;
    wire [0:0] _i_tile_x9y7__oe_x0y0_1;
    wire [0:0] _i_tile_x9y7__prog_dout;
    wire [0:0] _i_tile_x9y7__prog_we_o;
    wire [11:0] _i_sbox_x9y7sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x9y7sw__prog_dout;
    wire [0:0] _i_sbox_x9y7sw__prog_we_o;
    wire [11:0] _i_tile_x9y8__cu_u1y0n_L1;
    wire [11:0] _i_tile_x9y8__cu_u1y0s_L1;
    wire [0:0] _i_tile_x9y8__opin_x0y0_0;
    wire [0:0] _i_tile_x9y8__oe_x0y0_0;
    wire [0:0] _i_tile_x9y8__opin_x0y0_1;
    wire [0:0] _i_tile_x9y8__oe_x0y0_1;
    wire [0:0] _i_tile_x9y8__prog_dout;
    wire [0:0] _i_tile_x9y8__prog_we_o;
    wire [11:0] _i_sbox_x9y8sw__so_u1y0n_L1;
    wire [0:0] _i_sbox_x9y8sw__prog_dout;
    wire [0:0] _i_sbox_x9y8sw__prog_we_o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_buf_prog_rst_l1__Q;
    wire [0:0] _i_buf_prog_done_l1__Q;
    wire [0:0] _i_buf_prog_rst_l2__Q;
    wire [0:0] _i_buf_prog_done_l2__Q;
        
    sbox_ne_n_ex_ne i_sbox_x0y0ne (
        .bi_x1y0w_L1(_i_sbox_x1y1se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    t_io_w i_tile_x0y1 (
        .bi_x0y0n_L1(_i_sbox_x1y1sw__so_u1y0n_L1)
        ,.bi_x0y0s_L1(_i_sbox_x0y1ne__so_x0y0s_L1)
        ,.cu_x0y0n_L1(_i_tile_x0y1__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x0y1__cu_x0y0s_L1)
        ,.ipin_x0y0_0(ipin_x0y1_0)
        ,.opin_x0y0_0(_i_tile_x0y1__opin_x0y0_0)
        ,.oe_x0y0_0(_i_tile_x0y1__oe_x0y0_0)
        ,.ipin_x0y0_1(ipin_x0y1_1)
        ,.opin_x0y0_1(_i_tile_x0y1__opin_x0y0_1)
        ,.oe_x0y0_1(_i_tile_x0y1__oe_x0y0_1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_tile_x0y1__prog_dout)
        ,.prog_we_o(_i_tile_x0y1__prog_we_o)
        );
    sbox_ne_S_ex_e i_sbox_x0y1ne (
        .bi_x0y1s_L1(_i_sbox_x0y2ne__so_x0y0s_L1)
        ,.so_x0y0s_L1(_i_sbox_x0y1ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x1y2se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x0y1__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x0y2ne__prog_we_o)
        ,.prog_din(_i_sbox_x0y2ne__prog_dout)
        ,.prog_dout(_i_sbox_x0y1ne__prog_dout)
        ,.prog_we_o(_i_sbox_x0y1ne__prog_we_o)
        );
    sbox_se_e_ex_ne i_sbox_x0y1se (
        .bi_x0y0s_L1(_i_sbox_x0y1ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    t_io_w i_tile_x0y2 (
        .bi_x0y0n_L1(_i_sbox_x1y2sw__so_u1y0n_L1)
        ,.bi_x0y0s_L1(_i_sbox_x0y2ne__so_x0y0s_L1)
        ,.cu_x0y0n_L1(_i_tile_x0y2__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x0y2__cu_x0y0s_L1)
        ,.ipin_x0y0_0(ipin_x0y2_0)
        ,.opin_x0y0_0(_i_tile_x0y2__opin_x0y0_0)
        ,.oe_x0y0_0(_i_tile_x0y2__oe_x0y0_0)
        ,.ipin_x0y0_1(ipin_x0y2_1)
        ,.opin_x0y0_1(_i_tile_x0y2__opin_x0y0_1)
        ,.oe_x0y0_1(_i_tile_x0y2__oe_x0y0_1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_tile_x0y1__prog_we_o)
        ,.prog_din(_i_tile_x0y1__prog_dout)
        ,.prog_dout(_i_tile_x0y2__prog_dout)
        ,.prog_we_o(_i_tile_x0y2__prog_we_o)
        );
    sbox_ne_S_ex_e i_sbox_x0y2ne (
        .bi_x0y1s_L1(_i_sbox_x0y3ne__so_x0y0s_L1)
        ,.so_x0y0s_L1(_i_sbox_x0y2ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x1y3se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x0y2__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x0y3ne__prog_we_o)
        ,.prog_din(_i_sbox_x0y3ne__prog_dout)
        ,.prog_dout(_i_sbox_x0y2ne__prog_dout)
        ,.prog_we_o(_i_sbox_x0y2ne__prog_we_o)
        );
    sbox_se_e_ex_e i_sbox_x0y2se (
        .bi_x0v1n_L1(_i_sbox_x1y1sw__so_u1y0n_L1)
        ,.bi_x0y0s_L1(_i_sbox_x0y2ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    t_io_w i_tile_x0y3 (
        .bi_x0y0n_L1(_i_sbox_x1y3sw__so_u1y0n_L1)
        ,.bi_x0y0s_L1(_i_sbox_x0y3ne__so_x0y0s_L1)
        ,.cu_x0y0n_L1(_i_tile_x0y3__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x0y3__cu_x0y0s_L1)
        ,.ipin_x0y0_0(ipin_x0y3_0)
        ,.opin_x0y0_0(_i_tile_x0y3__opin_x0y0_0)
        ,.oe_x0y0_0(_i_tile_x0y3__oe_x0y0_0)
        ,.ipin_x0y0_1(ipin_x0y3_1)
        ,.opin_x0y0_1(_i_tile_x0y3__opin_x0y0_1)
        ,.oe_x0y0_1(_i_tile_x0y3__oe_x0y0_1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_tile_x0y2__prog_we_o)
        ,.prog_din(_i_tile_x0y2__prog_dout)
        ,.prog_dout(_i_tile_x0y3__prog_dout)
        ,.prog_we_o(_i_tile_x0y3__prog_we_o)
        );
    sbox_ne_S_ex_e i_sbox_x0y3ne (
        .bi_x0y1s_L1(_i_sbox_x0y4ne__so_x0y0s_L1)
        ,.so_x0y0s_L1(_i_sbox_x0y3ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x1y4se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x0y3__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x0y4ne__prog_we_o)
        ,.prog_din(_i_sbox_x0y4ne__prog_dout)
        ,.prog_dout(_i_sbox_x0y3ne__prog_dout)
        ,.prog_we_o(_i_sbox_x0y3ne__prog_we_o)
        );
    sbox_se_e_ex_e i_sbox_x0y3se (
        .bi_x0v1n_L1(_i_sbox_x1y2sw__so_u1y0n_L1)
        ,.bi_x0y0s_L1(_i_sbox_x0y3ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    t_io_w i_tile_x0y4 (
        .bi_x0y0n_L1(_i_sbox_x1y4sw__so_u1y0n_L1)
        ,.bi_x0y0s_L1(_i_sbox_x0y4ne__so_x0y0s_L1)
        ,.cu_x0y0n_L1(_i_tile_x0y4__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x0y4__cu_x0y0s_L1)
        ,.ipin_x0y0_0(ipin_x0y4_0)
        ,.opin_x0y0_0(_i_tile_x0y4__opin_x0y0_0)
        ,.oe_x0y0_0(_i_tile_x0y4__oe_x0y0_0)
        ,.ipin_x0y0_1(ipin_x0y4_1)
        ,.opin_x0y0_1(_i_tile_x0y4__opin_x0y0_1)
        ,.oe_x0y0_1(_i_tile_x0y4__oe_x0y0_1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_tile_x0y3__prog_we_o)
        ,.prog_din(_i_tile_x0y3__prog_dout)
        ,.prog_dout(_i_tile_x0y4__prog_dout)
        ,.prog_we_o(_i_tile_x0y4__prog_we_o)
        );
    sbox_ne_S_ex_e i_sbox_x0y4ne (
        .bi_x0y1s_L1(_i_sbox_x0y5ne__so_x0y0s_L1)
        ,.so_x0y0s_L1(_i_sbox_x0y4ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x1y5se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x0y4__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x0y5ne__prog_we_o)
        ,.prog_din(_i_sbox_x0y5ne__prog_dout)
        ,.prog_dout(_i_sbox_x0y4ne__prog_dout)
        ,.prog_we_o(_i_sbox_x0y4ne__prog_we_o)
        );
    sbox_se_e_ex_e i_sbox_x0y4se (
        .bi_x0v1n_L1(_i_sbox_x1y3sw__so_u1y0n_L1)
        ,.bi_x0y0s_L1(_i_sbox_x0y4ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    t_io_w i_tile_x0y5 (
        .bi_x0y0n_L1(_i_sbox_x1y5sw__so_u1y0n_L1)
        ,.bi_x0y0s_L1(_i_sbox_x0y5ne__so_x0y0s_L1)
        ,.cu_x0y0n_L1(_i_tile_x0y5__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x0y5__cu_x0y0s_L1)
        ,.ipin_x0y0_0(ipin_x0y5_0)
        ,.opin_x0y0_0(_i_tile_x0y5__opin_x0y0_0)
        ,.oe_x0y0_0(_i_tile_x0y5__oe_x0y0_0)
        ,.ipin_x0y0_1(ipin_x0y5_1)
        ,.opin_x0y0_1(_i_tile_x0y5__opin_x0y0_1)
        ,.oe_x0y0_1(_i_tile_x0y5__oe_x0y0_1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_tile_x0y4__prog_we_o)
        ,.prog_din(_i_tile_x0y4__prog_dout)
        ,.prog_dout(_i_tile_x0y5__prog_dout)
        ,.prog_we_o(_i_tile_x0y5__prog_we_o)
        );
    sbox_ne_S_ex_e i_sbox_x0y5ne (
        .bi_x0y1s_L1(_i_sbox_x0y6ne__so_x0y0s_L1)
        ,.so_x0y0s_L1(_i_sbox_x0y5ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x1y6se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x0y5__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x0y6ne__prog_we_o)
        ,.prog_din(_i_sbox_x0y6ne__prog_dout)
        ,.prog_dout(_i_sbox_x0y5ne__prog_dout)
        ,.prog_we_o(_i_sbox_x0y5ne__prog_we_o)
        );
    sbox_se_e_ex_e i_sbox_x0y5se (
        .bi_x0v1n_L1(_i_sbox_x1y4sw__so_u1y0n_L1)
        ,.bi_x0y0s_L1(_i_sbox_x0y5ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    t_io_w i_tile_x0y6 (
        .bi_x0y0n_L1(_i_sbox_x1y6sw__so_u1y0n_L1)
        ,.bi_x0y0s_L1(_i_sbox_x0y6ne__so_x0y0s_L1)
        ,.cu_x0y0n_L1(_i_tile_x0y6__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x0y6__cu_x0y0s_L1)
        ,.ipin_x0y0_0(ipin_x0y6_0)
        ,.opin_x0y0_0(_i_tile_x0y6__opin_x0y0_0)
        ,.oe_x0y0_0(_i_tile_x0y6__oe_x0y0_0)
        ,.ipin_x0y0_1(ipin_x0y6_1)
        ,.opin_x0y0_1(_i_tile_x0y6__opin_x0y0_1)
        ,.oe_x0y0_1(_i_tile_x0y6__oe_x0y0_1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_tile_x0y5__prog_we_o)
        ,.prog_din(_i_tile_x0y5__prog_dout)
        ,.prog_dout(_i_tile_x0y6__prog_dout)
        ,.prog_we_o(_i_tile_x0y6__prog_we_o)
        );
    sbox_ne_S_ex_e i_sbox_x0y6ne (
        .bi_x0y1s_L1(_i_sbox_x0y7ne__so_x0y0s_L1)
        ,.so_x0y0s_L1(_i_sbox_x0y6ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x1y7se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x0y6__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x0y7ne__prog_we_o)
        ,.prog_din(_i_sbox_x0y7ne__prog_dout)
        ,.prog_dout(_i_sbox_x0y6ne__prog_dout)
        ,.prog_we_o(_i_sbox_x0y6ne__prog_we_o)
        );
    sbox_se_e_ex_e i_sbox_x0y6se (
        .bi_x0v1n_L1(_i_sbox_x1y5sw__so_u1y0n_L1)
        ,.bi_x0y0s_L1(_i_sbox_x0y6ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    t_io_w i_tile_x0y7 (
        .bi_x0y0n_L1(_i_sbox_x1y7sw__so_u1y0n_L1)
        ,.bi_x0y0s_L1(_i_sbox_x0y7ne__so_x0y0s_L1)
        ,.cu_x0y0n_L1(_i_tile_x0y7__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x0y7__cu_x0y0s_L1)
        ,.ipin_x0y0_0(ipin_x0y7_0)
        ,.opin_x0y0_0(_i_tile_x0y7__opin_x0y0_0)
        ,.oe_x0y0_0(_i_tile_x0y7__oe_x0y0_0)
        ,.ipin_x0y0_1(ipin_x0y7_1)
        ,.opin_x0y0_1(_i_tile_x0y7__opin_x0y0_1)
        ,.oe_x0y0_1(_i_tile_x0y7__oe_x0y0_1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_tile_x0y6__prog_we_o)
        ,.prog_din(_i_tile_x0y6__prog_dout)
        ,.prog_dout(_i_tile_x0y7__prog_dout)
        ,.prog_we_o(_i_tile_x0y7__prog_we_o)
        );
    sbox_ne_S_ex_e i_sbox_x0y7ne (
        .bi_x0y1s_L1(_i_sbox_x0y8ne__so_x0y0s_L1)
        ,.so_x0y0s_L1(_i_sbox_x0y7ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x1y8se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x0y7__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x0y8ne__prog_we_o)
        ,.prog_din(_i_sbox_x0y8ne__prog_dout)
        ,.prog_dout(_i_sbox_x0y7ne__prog_dout)
        ,.prog_we_o(_i_sbox_x0y7ne__prog_we_o)
        );
    sbox_se_e_ex_e i_sbox_x0y7se (
        .bi_x0v1n_L1(_i_sbox_x1y6sw__so_u1y0n_L1)
        ,.bi_x0y0s_L1(_i_sbox_x0y7ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    t_io_w i_tile_x0y8 (
        .bi_x0y0n_L1(_i_sbox_x1y8sw__so_u1y0n_L1)
        ,.bi_x0y0s_L1(_i_sbox_x0y8ne__so_x0y0s_L1)
        ,.cu_x0y0n_L1(_i_tile_x0y8__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x0y8__cu_x0y0s_L1)
        ,.ipin_x0y0_0(ipin_x0y8_0)
        ,.opin_x0y0_0(_i_tile_x0y8__opin_x0y0_0)
        ,.oe_x0y0_0(_i_tile_x0y8__oe_x0y0_0)
        ,.ipin_x0y0_1(ipin_x0y8_1)
        ,.opin_x0y0_1(_i_tile_x0y8__opin_x0y0_1)
        ,.oe_x0y0_1(_i_tile_x0y8__oe_x0y0_1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_tile_x0y7__prog_we_o)
        ,.prog_din(_i_tile_x0y7__prog_dout)
        ,.prog_dout(_i_tile_x0y8__prog_dout)
        ,.prog_we_o(_i_tile_x0y8__prog_we_o)
        );
    sbox_ne_S_ex_es i_sbox_x0y8ne (
        .bi_x1y0w_L1(_i_sbox_x1y9se__so_x0v1w_L1)
        ,.so_x0y0s_L1(_i_sbox_x0y8ne__so_x0y0s_L1)
        ,.cu_x0y0s_L1(_i_tile_x0y8__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x0y8__prog_we_o)
        ,.prog_din(_i_tile_x0y8__prog_dout)
        ,.prog_dout(_i_sbox_x0y8ne__prog_dout)
        ,.prog_we_o(_i_sbox_x0y8ne__prog_we_o)
        );
    sbox_se_e_ex_e i_sbox_x0y8se (
        .bi_x0v1n_L1(_i_sbox_x1y7sw__so_u1y0n_L1)
        ,.bi_x0y0s_L1(_i_sbox_x0y8ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_se_e_ex_es i_sbox_x0y9se (
        .bi_x0v1n_L1(_i_sbox_x1y8sw__so_u1y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_ne_n_ex_n i_sbox_x1y0ne (
        .bi_x0y0e_L1(_i_sbox_x1y0nw__so_x0y0e_L1)
        ,.bi_x1y0w_L1(_i_sbox_x2y1se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_nw_E_ex_ne i_sbox_x1y0nw (
        .bi_u1y1s_L1(_i_sbox_x0y1ne__so_x0y0s_L1)
        ,.so_x0y0e_L1(_i_sbox_x1y0nw__so_x0y0e_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x0y1ne__prog_we_o)
        ,.prog_din(_i_sbox_x0y1ne__prog_dout)
        ,.prog_dout(_i_sbox_x1y0nw__prog_dout)
        ,.prog_we_o(_i_sbox_x1y0nw__prog_we_o)
        );
    tile_clb i_tile_x1y1 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x1y1__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x1y1__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x1y1sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x0y1ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x1y1sw__prog_we_o)
        ,.prog_din(_i_sbox_x1y1sw__prog_dout)
        ,.prog_dout(_i_tile_x1y1__prog_dout)
        ,.prog_we_o(_i_tile_x1y1__prog_we_o)
        );
    sbox_ne_S i_sbox_x1y1ne (
        .bi_x0y0e_L1(_i_sbox_x1y1nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x1y1ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x1y2ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x2y2se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x1y1__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x1y2se__prog_we_o)
        ,.prog_din(_i_sbox_x1y2se__prog_dout)
        ,.prog_dout(_i_sbox_x1y1ne__prog_dout)
        ,.prog_we_o(_i_sbox_x1y1ne__prog_we_o)
        );
    sbox_nw_E_ex_e i_sbox_x1y1nw (
        .bi_u1y0n_L1(_i_sbox_x1y1sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x1y1nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x0y2ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x1y1__prog_we_o)
        ,.prog_din(_i_tile_x1y1__prog_dout)
        ,.prog_dout(_i_sbox_x1y1nw__prog_dout)
        ,.prog_we_o(_i_sbox_x1y1nw__prog_we_o)
        );
    sbox_se_W_ex_n i_sbox_x1y1se (
        .bi_x0y0s_L1(_i_sbox_x1y1ne__so_x0y0s_L1)
        ,.so_x0v1w_L1(_i_sbox_x1y1se__so_x0v1w_L1)
        ,.bi_x1v1w_L1(_i_sbox_x2y1se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x1y1ne__prog_we_o)
        ,.prog_din(_i_sbox_x1y1ne__prog_dout)
        ,.prog_dout(_i_sbox_x1y1se__prog_dout)
        ,.prog_we_o(_i_sbox_x1y1se__prog_we_o)
        );
    sbox_sw_N_ex_ne i_sbox_x1y1sw (
        .bi_x0v1w_L1(_i_sbox_x1y1se__so_x0v1w_L1)
        ,.so_u1y0n_L1(_i_sbox_x1y1sw__so_u1y0n_L1)
        ,.cu_u1y0n_L1(_i_tile_x0y1__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x1y0nw__prog_we_o)
        ,.prog_din(_i_sbox_x1y0nw__prog_dout)
        ,.prog_dout(_i_sbox_x1y1sw__prog_dout)
        ,.prog_we_o(_i_sbox_x1y1sw__prog_we_o)
        );
    tile_clb i_tile_x1y2 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x1y2__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x1y2__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x1y2sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x0y2ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x1y2sw__prog_we_o)
        ,.prog_din(_i_sbox_x1y2sw__prog_dout)
        ,.prog_dout(_i_tile_x1y2__prog_dout)
        ,.prog_we_o(_i_tile_x1y2__prog_we_o)
        );
    sbox_ne_S i_sbox_x1y2ne (
        .bi_x0y0e_L1(_i_sbox_x1y2nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x1y2ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x1y3ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x2y3se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x1y2__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x1y3se__prog_we_o)
        ,.prog_din(_i_sbox_x1y3se__prog_dout)
        ,.prog_dout(_i_sbox_x1y2ne__prog_dout)
        ,.prog_we_o(_i_sbox_x1y2ne__prog_we_o)
        );
    sbox_nw_E_ex_e i_sbox_x1y2nw (
        .bi_u1y0n_L1(_i_sbox_x1y2sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x1y2nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x0y3ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x1y2__prog_we_o)
        ,.prog_din(_i_tile_x1y2__prog_dout)
        ,.prog_dout(_i_sbox_x1y2nw__prog_dout)
        ,.prog_we_o(_i_sbox_x1y2nw__prog_we_o)
        );
    sbox_se_W i_sbox_x1y2se (
        .bi_x0v1n_L1(_i_sbox_x2y1sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x1y2se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x1y2ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x2y2se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x1y2ne__prog_we_o)
        ,.prog_din(_i_sbox_x1y2ne__prog_dout)
        ,.prog_dout(_i_sbox_x1y2se__prog_dout)
        ,.prog_we_o(_i_sbox_x1y2se__prog_we_o)
        );
    sbox_sw_N_ex_e i_sbox_x1y2sw (
        .bi_u1v1n_L1(_i_sbox_x1y1sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x1y2sw__so_u1y0n_L1)
        ,.bi_x0v1w_L1(_i_sbox_x1y2se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x0y2__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x1y1nw__prog_we_o)
        ,.prog_din(_i_sbox_x1y1nw__prog_dout)
        ,.prog_dout(_i_sbox_x1y2sw__prog_dout)
        ,.prog_we_o(_i_sbox_x1y2sw__prog_we_o)
        );
    tile_clb i_tile_x1y3 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x1y3__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x1y3__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x1y3sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x0y3ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x1y3sw__prog_we_o)
        ,.prog_din(_i_sbox_x1y3sw__prog_dout)
        ,.prog_dout(_i_tile_x1y3__prog_dout)
        ,.prog_we_o(_i_tile_x1y3__prog_we_o)
        );
    sbox_ne_S i_sbox_x1y3ne (
        .bi_x0y0e_L1(_i_sbox_x1y3nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x1y3ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x1y4ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x2y4se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x1y3__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x1y4se__prog_we_o)
        ,.prog_din(_i_sbox_x1y4se__prog_dout)
        ,.prog_dout(_i_sbox_x1y3ne__prog_dout)
        ,.prog_we_o(_i_sbox_x1y3ne__prog_we_o)
        );
    sbox_nw_E_ex_e i_sbox_x1y3nw (
        .bi_u1y0n_L1(_i_sbox_x1y3sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x1y3nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x0y4ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x1y3__prog_we_o)
        ,.prog_din(_i_tile_x1y3__prog_dout)
        ,.prog_dout(_i_sbox_x1y3nw__prog_dout)
        ,.prog_we_o(_i_sbox_x1y3nw__prog_we_o)
        );
    sbox_se_W i_sbox_x1y3se (
        .bi_x0v1n_L1(_i_sbox_x2y2sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x1y3se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x1y3ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x2y3se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x1y3ne__prog_we_o)
        ,.prog_din(_i_sbox_x1y3ne__prog_dout)
        ,.prog_dout(_i_sbox_x1y3se__prog_dout)
        ,.prog_we_o(_i_sbox_x1y3se__prog_we_o)
        );
    sbox_sw_N_ex_e i_sbox_x1y3sw (
        .bi_u1v1n_L1(_i_sbox_x1y2sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x1y3sw__so_u1y0n_L1)
        ,.bi_x0v1w_L1(_i_sbox_x1y3se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x0y3__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x1y2nw__prog_we_o)
        ,.prog_din(_i_sbox_x1y2nw__prog_dout)
        ,.prog_dout(_i_sbox_x1y3sw__prog_dout)
        ,.prog_we_o(_i_sbox_x1y3sw__prog_we_o)
        );
    tile_clb i_tile_x1y4 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x1y4__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x1y4__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x1y4sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x0y4ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x1y4sw__prog_we_o)
        ,.prog_din(_i_sbox_x1y4sw__prog_dout)
        ,.prog_dout(_i_tile_x1y4__prog_dout)
        ,.prog_we_o(_i_tile_x1y4__prog_we_o)
        );
    sbox_ne_S i_sbox_x1y4ne (
        .bi_x0y0e_L1(_i_sbox_x1y4nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x1y4ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x1y5ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x2y5se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x1y4__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x1y5se__prog_we_o)
        ,.prog_din(_i_sbox_x1y5se__prog_dout)
        ,.prog_dout(_i_sbox_x1y4ne__prog_dout)
        ,.prog_we_o(_i_sbox_x1y4ne__prog_we_o)
        );
    sbox_nw_E_ex_e i_sbox_x1y4nw (
        .bi_u1y0n_L1(_i_sbox_x1y4sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x1y4nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x0y5ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x1y4__prog_we_o)
        ,.prog_din(_i_tile_x1y4__prog_dout)
        ,.prog_dout(_i_sbox_x1y4nw__prog_dout)
        ,.prog_we_o(_i_sbox_x1y4nw__prog_we_o)
        );
    sbox_se_W i_sbox_x1y4se (
        .bi_x0v1n_L1(_i_sbox_x2y3sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x1y4se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x1y4ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x2y4se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x1y4ne__prog_we_o)
        ,.prog_din(_i_sbox_x1y4ne__prog_dout)
        ,.prog_dout(_i_sbox_x1y4se__prog_dout)
        ,.prog_we_o(_i_sbox_x1y4se__prog_we_o)
        );
    sbox_sw_N_ex_e i_sbox_x1y4sw (
        .bi_u1v1n_L1(_i_sbox_x1y3sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x1y4sw__so_u1y0n_L1)
        ,.bi_x0v1w_L1(_i_sbox_x1y4se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x0y4__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x1y3nw__prog_we_o)
        ,.prog_din(_i_sbox_x1y3nw__prog_dout)
        ,.prog_dout(_i_sbox_x1y4sw__prog_dout)
        ,.prog_we_o(_i_sbox_x1y4sw__prog_we_o)
        );
    tile_clb i_tile_x1y5 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x1y5__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x1y5__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x1y5sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x0y5ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x1y5sw__prog_we_o)
        ,.prog_din(_i_sbox_x1y5sw__prog_dout)
        ,.prog_dout(_i_tile_x1y5__prog_dout)
        ,.prog_we_o(_i_tile_x1y5__prog_we_o)
        );
    sbox_ne_S i_sbox_x1y5ne (
        .bi_x0y0e_L1(_i_sbox_x1y5nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x1y5ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x1y6ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x2y6se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x1y5__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x1y6se__prog_we_o)
        ,.prog_din(_i_sbox_x1y6se__prog_dout)
        ,.prog_dout(_i_sbox_x1y5ne__prog_dout)
        ,.prog_we_o(_i_sbox_x1y5ne__prog_we_o)
        );
    sbox_nw_E_ex_e i_sbox_x1y5nw (
        .bi_u1y0n_L1(_i_sbox_x1y5sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x1y5nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x0y6ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x1y5__prog_we_o)
        ,.prog_din(_i_tile_x1y5__prog_dout)
        ,.prog_dout(_i_sbox_x1y5nw__prog_dout)
        ,.prog_we_o(_i_sbox_x1y5nw__prog_we_o)
        );
    sbox_se_W i_sbox_x1y5se (
        .bi_x0v1n_L1(_i_sbox_x2y4sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x1y5se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x1y5ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x2y5se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x1y5ne__prog_we_o)
        ,.prog_din(_i_sbox_x1y5ne__prog_dout)
        ,.prog_dout(_i_sbox_x1y5se__prog_dout)
        ,.prog_we_o(_i_sbox_x1y5se__prog_we_o)
        );
    sbox_sw_N_ex_e i_sbox_x1y5sw (
        .bi_u1v1n_L1(_i_sbox_x1y4sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x1y5sw__so_u1y0n_L1)
        ,.bi_x0v1w_L1(_i_sbox_x1y5se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x0y5__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x1y4nw__prog_we_o)
        ,.prog_din(_i_sbox_x1y4nw__prog_dout)
        ,.prog_dout(_i_sbox_x1y5sw__prog_dout)
        ,.prog_we_o(_i_sbox_x1y5sw__prog_we_o)
        );
    tile_clb i_tile_x1y6 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x1y6__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x1y6__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x1y6sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x0y6ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x1y6sw__prog_we_o)
        ,.prog_din(_i_sbox_x1y6sw__prog_dout)
        ,.prog_dout(_i_tile_x1y6__prog_dout)
        ,.prog_we_o(_i_tile_x1y6__prog_we_o)
        );
    sbox_ne_S i_sbox_x1y6ne (
        .bi_x0y0e_L1(_i_sbox_x1y6nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x1y6ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x1y7ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x2y7se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x1y6__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x1y7se__prog_we_o)
        ,.prog_din(_i_sbox_x1y7se__prog_dout)
        ,.prog_dout(_i_sbox_x1y6ne__prog_dout)
        ,.prog_we_o(_i_sbox_x1y6ne__prog_we_o)
        );
    sbox_nw_E_ex_e i_sbox_x1y6nw (
        .bi_u1y0n_L1(_i_sbox_x1y6sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x1y6nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x0y7ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x1y6__prog_we_o)
        ,.prog_din(_i_tile_x1y6__prog_dout)
        ,.prog_dout(_i_sbox_x1y6nw__prog_dout)
        ,.prog_we_o(_i_sbox_x1y6nw__prog_we_o)
        );
    sbox_se_W i_sbox_x1y6se (
        .bi_x0v1n_L1(_i_sbox_x2y5sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x1y6se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x1y6ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x2y6se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x1y6ne__prog_we_o)
        ,.prog_din(_i_sbox_x1y6ne__prog_dout)
        ,.prog_dout(_i_sbox_x1y6se__prog_dout)
        ,.prog_we_o(_i_sbox_x1y6se__prog_we_o)
        );
    sbox_sw_N_ex_e i_sbox_x1y6sw (
        .bi_u1v1n_L1(_i_sbox_x1y5sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x1y6sw__so_u1y0n_L1)
        ,.bi_x0v1w_L1(_i_sbox_x1y6se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x0y6__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x1y5nw__prog_we_o)
        ,.prog_din(_i_sbox_x1y5nw__prog_dout)
        ,.prog_dout(_i_sbox_x1y6sw__prog_dout)
        ,.prog_we_o(_i_sbox_x1y6sw__prog_we_o)
        );
    tile_clb i_tile_x1y7 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x1y7__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x1y7__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x1y7sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x0y7ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x1y7sw__prog_we_o)
        ,.prog_din(_i_sbox_x1y7sw__prog_dout)
        ,.prog_dout(_i_tile_x1y7__prog_dout)
        ,.prog_we_o(_i_tile_x1y7__prog_we_o)
        );
    sbox_ne_S i_sbox_x1y7ne (
        .bi_x0y0e_L1(_i_sbox_x1y7nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x1y7ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x1y8ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x2y8se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x1y7__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x1y8se__prog_we_o)
        ,.prog_din(_i_sbox_x1y8se__prog_dout)
        ,.prog_dout(_i_sbox_x1y7ne__prog_dout)
        ,.prog_we_o(_i_sbox_x1y7ne__prog_we_o)
        );
    sbox_nw_E_ex_e i_sbox_x1y7nw (
        .bi_u1y0n_L1(_i_sbox_x1y7sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x1y7nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x0y8ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x1y7__prog_we_o)
        ,.prog_din(_i_tile_x1y7__prog_dout)
        ,.prog_dout(_i_sbox_x1y7nw__prog_dout)
        ,.prog_we_o(_i_sbox_x1y7nw__prog_we_o)
        );
    sbox_se_W i_sbox_x1y7se (
        .bi_x0v1n_L1(_i_sbox_x2y6sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x1y7se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x1y7ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x2y7se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x1y7ne__prog_we_o)
        ,.prog_din(_i_sbox_x1y7ne__prog_dout)
        ,.prog_dout(_i_sbox_x1y7se__prog_dout)
        ,.prog_we_o(_i_sbox_x1y7se__prog_we_o)
        );
    sbox_sw_N_ex_e i_sbox_x1y7sw (
        .bi_u1v1n_L1(_i_sbox_x1y6sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x1y7sw__so_u1y0n_L1)
        ,.bi_x0v1w_L1(_i_sbox_x1y7se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x0y7__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x1y6nw__prog_we_o)
        ,.prog_din(_i_sbox_x1y6nw__prog_dout)
        ,.prog_dout(_i_sbox_x1y7sw__prog_dout)
        ,.prog_we_o(_i_sbox_x1y7sw__prog_we_o)
        );
    tile_clb i_tile_x1y8 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x1y8__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x1y8__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x1y8sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x0y8ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x1y8sw__prog_we_o)
        ,.prog_din(_i_sbox_x1y8sw__prog_dout)
        ,.prog_dout(_i_tile_x1y8__prog_dout)
        ,.prog_we_o(_i_tile_x1y8__prog_we_o)
        );
    sbox_ne_S_ex_s i_sbox_x1y8ne (
        .bi_x0y0e_L1(_i_sbox_x1y8nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x1y8ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x2y9se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x1y8__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x1y9se__prog_we_o)
        ,.prog_din(_i_sbox_x1y9se__prog_dout)
        ,.prog_dout(_i_sbox_x1y8ne__prog_dout)
        ,.prog_we_o(_i_sbox_x1y8ne__prog_we_o)
        );
    sbox_nw_E_ex_es i_sbox_x1y8nw (
        .bi_u1y0n_L1(_i_sbox_x1y8sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x1y8nw__so_x0y0e_L1)
        ,.cu_x0y0e_L1(_i_tile_x1y9__cu_x0v1e_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x1y8__prog_we_o)
        ,.prog_din(_i_tile_x1y8__prog_dout)
        ,.prog_dout(_i_sbox_x1y8nw__prog_dout)
        ,.prog_we_o(_i_sbox_x1y8nw__prog_we_o)
        );
    sbox_se_W i_sbox_x1y8se (
        .bi_x0v1n_L1(_i_sbox_x2y7sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x1y8se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x1y8ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x2y8se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x1y8ne__prog_we_o)
        ,.prog_din(_i_sbox_x1y8ne__prog_dout)
        ,.prog_dout(_i_sbox_x1y8se__prog_dout)
        ,.prog_we_o(_i_sbox_x1y8se__prog_we_o)
        );
    sbox_sw_N_ex_e i_sbox_x1y8sw (
        .bi_u1v1n_L1(_i_sbox_x1y7sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x1y8sw__so_u1y0n_L1)
        ,.bi_x0v1w_L1(_i_sbox_x1y8se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x0y8__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x1y7nw__prog_we_o)
        ,.prog_din(_i_sbox_x1y7nw__prog_dout)
        ,.prog_dout(_i_sbox_x1y8sw__prog_dout)
        ,.prog_we_o(_i_sbox_x1y8sw__prog_we_o)
        );
    t_io_n i_tile_x1y9 (
        .bi_x0v1e_L1(_i_sbox_x1y8nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x1y9se__so_x0v1w_L1)
        ,.cu_x0v1e_L1(_i_tile_x1y9__cu_x0v1e_L1)
        ,.cu_x0v1w_L1(_i_tile_x1y9__cu_x0v1w_L1)
        ,.ipin_x0y0_0(ipin_x1y9_0)
        ,.opin_x0y0_0(_i_tile_x1y9__opin_x0y0_0)
        ,.oe_x0y0_0(_i_tile_x1y9__oe_x0y0_0)
        ,.ipin_x0y0_1(ipin_x1y9_1)
        ,.opin_x0y0_1(_i_tile_x1y9__opin_x0y0_1)
        ,.oe_x0y0_1(_i_tile_x1y9__oe_x0y0_1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x1y8nw__prog_we_o)
        ,.prog_din(_i_sbox_x1y8nw__prog_dout)
        ,.prog_dout(_i_tile_x1y9__prog_dout)
        ,.prog_we_o(_i_tile_x1y9__prog_we_o)
        );
    sbox_se_W_ex_s i_sbox_x1y9se (
        .bi_x0v1n_L1(_i_sbox_x2y8sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x1y9se__so_x0v1w_L1)
        ,.bi_x1v1w_L1(_i_sbox_x2y9se__so_x0v1w_L1)
        ,.cu_x0v1w_L1(_i_tile_x1y9__cu_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x1y9__prog_we_o)
        ,.prog_din(_i_tile_x1y9__prog_dout)
        ,.prog_dout(_i_sbox_x1y9se__prog_dout)
        ,.prog_we_o(_i_sbox_x1y9se__prog_we_o)
        );
    sbox_sw_s_ex_es i_sbox_x1y9sw (
        .bi_x0v1w_L1(_i_sbox_x1y9se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_ne_n_ex_n i_sbox_x2y0ne (
        .bi_x0y0e_L1(_i_sbox_x2y0nw__so_x0y0e_L1)
        ,.bi_x1y0w_L1(_i_sbox_x3y1se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_nw_E_ex_n i_sbox_x2y0nw (
        .bi_u1y0e_L1(_i_sbox_x1y0nw__so_x0y0e_L1)
        ,.so_x0y0e_L1(_i_sbox_x2y0nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x1y1ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x1y1se__prog_we_o)
        ,.prog_din(_i_sbox_x1y1se__prog_dout)
        ,.prog_dout(_i_sbox_x2y0nw__prog_dout)
        ,.prog_we_o(_i_sbox_x2y0nw__prog_we_o)
        );
    tile_clb i_tile_x2y1 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x2y1__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x2y1__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x2y1sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x1y1ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x2y1sw__prog_we_o)
        ,.prog_din(_i_sbox_x2y1sw__prog_dout)
        ,.prog_dout(_i_tile_x2y1__prog_dout)
        ,.prog_we_o(_i_tile_x2y1__prog_we_o)
        );
    sbox_ne_S i_sbox_x2y1ne (
        .bi_x0y0e_L1(_i_sbox_x2y1nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x2y1ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x2y2ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x3y2se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x2y1__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x2y2se__prog_we_o)
        ,.prog_din(_i_sbox_x2y2se__prog_dout)
        ,.prog_dout(_i_sbox_x2y1ne__prog_dout)
        ,.prog_we_o(_i_sbox_x2y1ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x2y1nw (
        .bi_u1y0n_L1(_i_sbox_x2y1sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x2y1nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x1y1nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x1y2ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x2y1__prog_we_o)
        ,.prog_din(_i_tile_x2y1__prog_dout)
        ,.prog_dout(_i_sbox_x2y1nw__prog_dout)
        ,.prog_we_o(_i_sbox_x2y1nw__prog_we_o)
        );
    sbox_se_W_ex_n i_sbox_x2y1se (
        .bi_x0y0s_L1(_i_sbox_x2y1ne__so_x0y0s_L1)
        ,.so_x0v1w_L1(_i_sbox_x2y1se__so_x0v1w_L1)
        ,.bi_x1v1w_L1(_i_sbox_x3y1se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x2y1ne__prog_we_o)
        ,.prog_din(_i_sbox_x2y1ne__prog_dout)
        ,.prog_dout(_i_sbox_x2y1se__prog_dout)
        ,.prog_we_o(_i_sbox_x2y1se__prog_we_o)
        );
    sbox_sw_N_ex_n i_sbox_x2y1sw (
        .bi_u1v1e_L1(_i_sbox_x1y0nw__so_x0y0e_L1)
        ,.so_u1y0n_L1(_i_sbox_x2y1sw__so_u1y0n_L1)
        ,.bi_x0v1w_L1(_i_sbox_x2y1se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x1y1__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x2y0nw__prog_we_o)
        ,.prog_din(_i_sbox_x2y0nw__prog_dout)
        ,.prog_dout(_i_sbox_x2y1sw__prog_dout)
        ,.prog_we_o(_i_sbox_x2y1sw__prog_we_o)
        );
    tile_clb i_tile_x2y2 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x2y2__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x2y2__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x2y2sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x1y2ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x2y2sw__prog_we_o)
        ,.prog_din(_i_sbox_x2y2sw__prog_dout)
        ,.prog_dout(_i_tile_x2y2__prog_dout)
        ,.prog_we_o(_i_tile_x2y2__prog_we_o)
        );
    sbox_ne_S i_sbox_x2y2ne (
        .bi_x0y0e_L1(_i_sbox_x2y2nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x2y2ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x2y3ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x3y3se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x2y2__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x2y3se__prog_we_o)
        ,.prog_din(_i_sbox_x2y3se__prog_dout)
        ,.prog_dout(_i_sbox_x2y2ne__prog_dout)
        ,.prog_we_o(_i_sbox_x2y2ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x2y2nw (
        .bi_u1y0n_L1(_i_sbox_x2y2sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x2y2nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x1y2nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x1y3ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x2y2__prog_we_o)
        ,.prog_din(_i_tile_x2y2__prog_dout)
        ,.prog_dout(_i_sbox_x2y2nw__prog_dout)
        ,.prog_we_o(_i_sbox_x2y2nw__prog_we_o)
        );
    sbox_se_W i_sbox_x2y2se (
        .bi_x0v1n_L1(_i_sbox_x3y1sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x2y2se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x2y2ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x3y2se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x2y2ne__prog_we_o)
        ,.prog_din(_i_sbox_x2y2ne__prog_dout)
        ,.prog_dout(_i_sbox_x2y2se__prog_dout)
        ,.prog_we_o(_i_sbox_x2y2se__prog_we_o)
        );
    sbox_sw_N i_sbox_x2y2sw (
        .bi_u1v1n_L1(_i_sbox_x2y1sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x2y2sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x1y1nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x2y2se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x1y2__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x2y1nw__prog_we_o)
        ,.prog_din(_i_sbox_x2y1nw__prog_dout)
        ,.prog_dout(_i_sbox_x2y2sw__prog_dout)
        ,.prog_we_o(_i_sbox_x2y2sw__prog_we_o)
        );
    tile_clb i_tile_x2y3 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x2y3__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x2y3__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x2y3sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x1y3ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x2y3sw__prog_we_o)
        ,.prog_din(_i_sbox_x2y3sw__prog_dout)
        ,.prog_dout(_i_tile_x2y3__prog_dout)
        ,.prog_we_o(_i_tile_x2y3__prog_we_o)
        );
    sbox_ne_S i_sbox_x2y3ne (
        .bi_x0y0e_L1(_i_sbox_x2y3nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x2y3ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x2y4ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x3y4se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x2y3__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x2y4se__prog_we_o)
        ,.prog_din(_i_sbox_x2y4se__prog_dout)
        ,.prog_dout(_i_sbox_x2y3ne__prog_dout)
        ,.prog_we_o(_i_sbox_x2y3ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x2y3nw (
        .bi_u1y0n_L1(_i_sbox_x2y3sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x2y3nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x1y3nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x1y4ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x2y3__prog_we_o)
        ,.prog_din(_i_tile_x2y3__prog_dout)
        ,.prog_dout(_i_sbox_x2y3nw__prog_dout)
        ,.prog_we_o(_i_sbox_x2y3nw__prog_we_o)
        );
    sbox_se_W i_sbox_x2y3se (
        .bi_x0v1n_L1(_i_sbox_x3y2sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x2y3se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x2y3ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x3y3se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x2y3ne__prog_we_o)
        ,.prog_din(_i_sbox_x2y3ne__prog_dout)
        ,.prog_dout(_i_sbox_x2y3se__prog_dout)
        ,.prog_we_o(_i_sbox_x2y3se__prog_we_o)
        );
    sbox_sw_N i_sbox_x2y3sw (
        .bi_u1v1n_L1(_i_sbox_x2y2sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x2y3sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x1y2nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x2y3se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x1y3__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x2y2nw__prog_we_o)
        ,.prog_din(_i_sbox_x2y2nw__prog_dout)
        ,.prog_dout(_i_sbox_x2y3sw__prog_dout)
        ,.prog_we_o(_i_sbox_x2y3sw__prog_we_o)
        );
    tile_clb i_tile_x2y4 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x2y4__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x2y4__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x2y4sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x1y4ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x2y4sw__prog_we_o)
        ,.prog_din(_i_sbox_x2y4sw__prog_dout)
        ,.prog_dout(_i_tile_x2y4__prog_dout)
        ,.prog_we_o(_i_tile_x2y4__prog_we_o)
        );
    sbox_ne_S i_sbox_x2y4ne (
        .bi_x0y0e_L1(_i_sbox_x2y4nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x2y4ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x2y5ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x3y5se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x2y4__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x2y5se__prog_we_o)
        ,.prog_din(_i_sbox_x2y5se__prog_dout)
        ,.prog_dout(_i_sbox_x2y4ne__prog_dout)
        ,.prog_we_o(_i_sbox_x2y4ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x2y4nw (
        .bi_u1y0n_L1(_i_sbox_x2y4sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x2y4nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x1y4nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x1y5ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x2y4__prog_we_o)
        ,.prog_din(_i_tile_x2y4__prog_dout)
        ,.prog_dout(_i_sbox_x2y4nw__prog_dout)
        ,.prog_we_o(_i_sbox_x2y4nw__prog_we_o)
        );
    sbox_se_W i_sbox_x2y4se (
        .bi_x0v1n_L1(_i_sbox_x3y3sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x2y4se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x2y4ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x3y4se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x2y4ne__prog_we_o)
        ,.prog_din(_i_sbox_x2y4ne__prog_dout)
        ,.prog_dout(_i_sbox_x2y4se__prog_dout)
        ,.prog_we_o(_i_sbox_x2y4se__prog_we_o)
        );
    sbox_sw_N i_sbox_x2y4sw (
        .bi_u1v1n_L1(_i_sbox_x2y3sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x2y4sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x1y3nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x2y4se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x1y4__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x2y3nw__prog_we_o)
        ,.prog_din(_i_sbox_x2y3nw__prog_dout)
        ,.prog_dout(_i_sbox_x2y4sw__prog_dout)
        ,.prog_we_o(_i_sbox_x2y4sw__prog_we_o)
        );
    tile_clb i_tile_x2y5 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x2y5__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x2y5__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x2y5sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x1y5ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x2y5sw__prog_we_o)
        ,.prog_din(_i_sbox_x2y5sw__prog_dout)
        ,.prog_dout(_i_tile_x2y5__prog_dout)
        ,.prog_we_o(_i_tile_x2y5__prog_we_o)
        );
    sbox_ne_S i_sbox_x2y5ne (
        .bi_x0y0e_L1(_i_sbox_x2y5nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x2y5ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x2y6ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x3y6se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x2y5__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x2y6se__prog_we_o)
        ,.prog_din(_i_sbox_x2y6se__prog_dout)
        ,.prog_dout(_i_sbox_x2y5ne__prog_dout)
        ,.prog_we_o(_i_sbox_x2y5ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x2y5nw (
        .bi_u1y0n_L1(_i_sbox_x2y5sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x2y5nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x1y5nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x1y6ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x2y5__prog_we_o)
        ,.prog_din(_i_tile_x2y5__prog_dout)
        ,.prog_dout(_i_sbox_x2y5nw__prog_dout)
        ,.prog_we_o(_i_sbox_x2y5nw__prog_we_o)
        );
    sbox_se_W i_sbox_x2y5se (
        .bi_x0v1n_L1(_i_sbox_x3y4sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x2y5se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x2y5ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x3y5se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x2y5ne__prog_we_o)
        ,.prog_din(_i_sbox_x2y5ne__prog_dout)
        ,.prog_dout(_i_sbox_x2y5se__prog_dout)
        ,.prog_we_o(_i_sbox_x2y5se__prog_we_o)
        );
    sbox_sw_N i_sbox_x2y5sw (
        .bi_u1v1n_L1(_i_sbox_x2y4sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x2y5sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x1y4nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x2y5se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x1y5__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x2y4nw__prog_we_o)
        ,.prog_din(_i_sbox_x2y4nw__prog_dout)
        ,.prog_dout(_i_sbox_x2y5sw__prog_dout)
        ,.prog_we_o(_i_sbox_x2y5sw__prog_we_o)
        );
    tile_clb i_tile_x2y6 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x2y6__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x2y6__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x2y6sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x1y6ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x2y6sw__prog_we_o)
        ,.prog_din(_i_sbox_x2y6sw__prog_dout)
        ,.prog_dout(_i_tile_x2y6__prog_dout)
        ,.prog_we_o(_i_tile_x2y6__prog_we_o)
        );
    sbox_ne_S i_sbox_x2y6ne (
        .bi_x0y0e_L1(_i_sbox_x2y6nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x2y6ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x2y7ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x3y7se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x2y6__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x2y7se__prog_we_o)
        ,.prog_din(_i_sbox_x2y7se__prog_dout)
        ,.prog_dout(_i_sbox_x2y6ne__prog_dout)
        ,.prog_we_o(_i_sbox_x2y6ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x2y6nw (
        .bi_u1y0n_L1(_i_sbox_x2y6sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x2y6nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x1y6nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x1y7ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x2y6__prog_we_o)
        ,.prog_din(_i_tile_x2y6__prog_dout)
        ,.prog_dout(_i_sbox_x2y6nw__prog_dout)
        ,.prog_we_o(_i_sbox_x2y6nw__prog_we_o)
        );
    sbox_se_W i_sbox_x2y6se (
        .bi_x0v1n_L1(_i_sbox_x3y5sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x2y6se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x2y6ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x3y6se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x2y6ne__prog_we_o)
        ,.prog_din(_i_sbox_x2y6ne__prog_dout)
        ,.prog_dout(_i_sbox_x2y6se__prog_dout)
        ,.prog_we_o(_i_sbox_x2y6se__prog_we_o)
        );
    sbox_sw_N i_sbox_x2y6sw (
        .bi_u1v1n_L1(_i_sbox_x2y5sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x2y6sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x1y5nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x2y6se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x1y6__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x2y5nw__prog_we_o)
        ,.prog_din(_i_sbox_x2y5nw__prog_dout)
        ,.prog_dout(_i_sbox_x2y6sw__prog_dout)
        ,.prog_we_o(_i_sbox_x2y6sw__prog_we_o)
        );
    tile_clb i_tile_x2y7 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x2y7__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x2y7__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x2y7sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x1y7ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x2y7sw__prog_we_o)
        ,.prog_din(_i_sbox_x2y7sw__prog_dout)
        ,.prog_dout(_i_tile_x2y7__prog_dout)
        ,.prog_we_o(_i_tile_x2y7__prog_we_o)
        );
    sbox_ne_S i_sbox_x2y7ne (
        .bi_x0y0e_L1(_i_sbox_x2y7nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x2y7ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x2y8ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x3y8se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x2y7__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x2y8se__prog_we_o)
        ,.prog_din(_i_sbox_x2y8se__prog_dout)
        ,.prog_dout(_i_sbox_x2y7ne__prog_dout)
        ,.prog_we_o(_i_sbox_x2y7ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x2y7nw (
        .bi_u1y0n_L1(_i_sbox_x2y7sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x2y7nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x1y7nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x1y8ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x2y7__prog_we_o)
        ,.prog_din(_i_tile_x2y7__prog_dout)
        ,.prog_dout(_i_sbox_x2y7nw__prog_dout)
        ,.prog_we_o(_i_sbox_x2y7nw__prog_we_o)
        );
    sbox_se_W i_sbox_x2y7se (
        .bi_x0v1n_L1(_i_sbox_x3y6sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x2y7se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x2y7ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x3y7se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x2y7ne__prog_we_o)
        ,.prog_din(_i_sbox_x2y7ne__prog_dout)
        ,.prog_dout(_i_sbox_x2y7se__prog_dout)
        ,.prog_we_o(_i_sbox_x2y7se__prog_we_o)
        );
    sbox_sw_N i_sbox_x2y7sw (
        .bi_u1v1n_L1(_i_sbox_x2y6sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x2y7sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x1y6nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x2y7se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x1y7__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x2y6nw__prog_we_o)
        ,.prog_din(_i_sbox_x2y6nw__prog_dout)
        ,.prog_dout(_i_sbox_x2y7sw__prog_dout)
        ,.prog_we_o(_i_sbox_x2y7sw__prog_we_o)
        );
    tile_clb i_tile_x2y8 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x2y8__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x2y8__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x2y8sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x1y8ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x2y8sw__prog_we_o)
        ,.prog_din(_i_sbox_x2y8sw__prog_dout)
        ,.prog_dout(_i_tile_x2y8__prog_dout)
        ,.prog_we_o(_i_tile_x2y8__prog_we_o)
        );
    sbox_ne_S_ex_s i_sbox_x2y8ne (
        .bi_x0y0e_L1(_i_sbox_x2y8nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x2y8ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x3y9se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x2y8__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x2y9se__prog_we_o)
        ,.prog_din(_i_sbox_x2y9se__prog_dout)
        ,.prog_dout(_i_sbox_x2y8ne__prog_dout)
        ,.prog_we_o(_i_sbox_x2y8ne__prog_we_o)
        );
    sbox_nw_E_ex_s i_sbox_x2y8nw (
        .bi_u1y0n_L1(_i_sbox_x2y8sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x2y8nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x1y8nw__so_x0y0e_L1)
        ,.cu_x0y0e_L1(_i_tile_x2y9__cu_x0v1e_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x2y8__prog_we_o)
        ,.prog_din(_i_tile_x2y8__prog_dout)
        ,.prog_dout(_i_sbox_x2y8nw__prog_dout)
        ,.prog_we_o(_i_sbox_x2y8nw__prog_we_o)
        );
    sbox_se_W i_sbox_x2y8se (
        .bi_x0v1n_L1(_i_sbox_x3y7sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x2y8se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x2y8ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x3y8se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x2y8ne__prog_we_o)
        ,.prog_din(_i_sbox_x2y8ne__prog_dout)
        ,.prog_dout(_i_sbox_x2y8se__prog_dout)
        ,.prog_we_o(_i_sbox_x2y8se__prog_we_o)
        );
    sbox_sw_N i_sbox_x2y8sw (
        .bi_u1v1n_L1(_i_sbox_x2y7sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x2y8sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x1y7nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x2y8se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x1y8__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x2y7nw__prog_we_o)
        ,.prog_din(_i_sbox_x2y7nw__prog_dout)
        ,.prog_dout(_i_sbox_x2y8sw__prog_dout)
        ,.prog_we_o(_i_sbox_x2y8sw__prog_we_o)
        );
    t_io_n i_tile_x2y9 (
        .bi_x0v1e_L1(_i_sbox_x2y8nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x2y9se__so_x0v1w_L1)
        ,.cu_x0v1e_L1(_i_tile_x2y9__cu_x0v1e_L1)
        ,.cu_x0v1w_L1(_i_tile_x2y9__cu_x0v1w_L1)
        ,.ipin_x0y0_0(ipin_x2y9_0)
        ,.opin_x0y0_0(_i_tile_x2y9__opin_x0y0_0)
        ,.oe_x0y0_0(_i_tile_x2y9__oe_x0y0_0)
        ,.ipin_x0y0_1(ipin_x2y9_1)
        ,.opin_x0y0_1(_i_tile_x2y9__opin_x0y0_1)
        ,.oe_x0y0_1(_i_tile_x2y9__oe_x0y0_1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x2y8nw__prog_we_o)
        ,.prog_din(_i_sbox_x2y8nw__prog_dout)
        ,.prog_dout(_i_tile_x2y9__prog_dout)
        ,.prog_we_o(_i_tile_x2y9__prog_we_o)
        );
    sbox_se_W_ex_s i_sbox_x2y9se (
        .bi_x0v1n_L1(_i_sbox_x3y8sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x2y9se__so_x0v1w_L1)
        ,.bi_x1v1w_L1(_i_sbox_x3y9se__so_x0v1w_L1)
        ,.cu_x0v1w_L1(_i_tile_x2y9__cu_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x2y9__prog_we_o)
        ,.prog_din(_i_tile_x2y9__prog_dout)
        ,.prog_dout(_i_sbox_x2y9se__prog_dout)
        ,.prog_we_o(_i_sbox_x2y9se__prog_we_o)
        );
    sbox_sw_s_ex_s i_sbox_x2y9sw (
        .bi_u1v1e_L1(_i_sbox_x1y8nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x2y9se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_ne_n_ex_n i_sbox_x3y0ne (
        .bi_x0y0e_L1(_i_sbox_x3y0nw__so_x0y0e_L1)
        ,.bi_x1y0w_L1(_i_sbox_x4y1se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_nw_E_ex_n i_sbox_x3y0nw (
        .bi_u1y0e_L1(_i_sbox_x2y0nw__so_x0y0e_L1)
        ,.so_x0y0e_L1(_i_sbox_x3y0nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x2y1ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x2y1se__prog_we_o)
        ,.prog_din(_i_sbox_x2y1se__prog_dout)
        ,.prog_dout(_i_sbox_x3y0nw__prog_dout)
        ,.prog_we_o(_i_sbox_x3y0nw__prog_we_o)
        );
    tile_clb i_tile_x3y1 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x3y1__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x3y1__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x3y1sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x2y1ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x3y1sw__prog_we_o)
        ,.prog_din(_i_sbox_x3y1sw__prog_dout)
        ,.prog_dout(_i_tile_x3y1__prog_dout)
        ,.prog_we_o(_i_tile_x3y1__prog_we_o)
        );
    sbox_ne_S i_sbox_x3y1ne (
        .bi_x0y0e_L1(_i_sbox_x3y1nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x3y1ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x3y2ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x4y2se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x3y1__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x3y2se__prog_we_o)
        ,.prog_din(_i_sbox_x3y2se__prog_dout)
        ,.prog_dout(_i_sbox_x3y1ne__prog_dout)
        ,.prog_we_o(_i_sbox_x3y1ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x3y1nw (
        .bi_u1y0n_L1(_i_sbox_x3y1sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x3y1nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x2y1nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x2y2ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x3y1__prog_we_o)
        ,.prog_din(_i_tile_x3y1__prog_dout)
        ,.prog_dout(_i_sbox_x3y1nw__prog_dout)
        ,.prog_we_o(_i_sbox_x3y1nw__prog_we_o)
        );
    sbox_se_W_ex_n i_sbox_x3y1se (
        .bi_x0y0s_L1(_i_sbox_x3y1ne__so_x0y0s_L1)
        ,.so_x0v1w_L1(_i_sbox_x3y1se__so_x0v1w_L1)
        ,.bi_x1v1w_L1(_i_sbox_x4y1se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x3y1ne__prog_we_o)
        ,.prog_din(_i_sbox_x3y1ne__prog_dout)
        ,.prog_dout(_i_sbox_x3y1se__prog_dout)
        ,.prog_we_o(_i_sbox_x3y1se__prog_we_o)
        );
    sbox_sw_N_ex_n i_sbox_x3y1sw (
        .bi_u1v1e_L1(_i_sbox_x2y0nw__so_x0y0e_L1)
        ,.so_u1y0n_L1(_i_sbox_x3y1sw__so_u1y0n_L1)
        ,.bi_x0v1w_L1(_i_sbox_x3y1se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x2y1__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x3y0nw__prog_we_o)
        ,.prog_din(_i_sbox_x3y0nw__prog_dout)
        ,.prog_dout(_i_sbox_x3y1sw__prog_dout)
        ,.prog_we_o(_i_sbox_x3y1sw__prog_we_o)
        );
    tile_clb i_tile_x3y2 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x3y2__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x3y2__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x3y2sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x2y2ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x3y2sw__prog_we_o)
        ,.prog_din(_i_sbox_x3y2sw__prog_dout)
        ,.prog_dout(_i_tile_x3y2__prog_dout)
        ,.prog_we_o(_i_tile_x3y2__prog_we_o)
        );
    sbox_ne_S i_sbox_x3y2ne (
        .bi_x0y0e_L1(_i_sbox_x3y2nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x3y2ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x3y3ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x4y3se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x3y2__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x3y3se__prog_we_o)
        ,.prog_din(_i_sbox_x3y3se__prog_dout)
        ,.prog_dout(_i_sbox_x3y2ne__prog_dout)
        ,.prog_we_o(_i_sbox_x3y2ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x3y2nw (
        .bi_u1y0n_L1(_i_sbox_x3y2sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x3y2nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x2y2nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x2y3ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x3y2__prog_we_o)
        ,.prog_din(_i_tile_x3y2__prog_dout)
        ,.prog_dout(_i_sbox_x3y2nw__prog_dout)
        ,.prog_we_o(_i_sbox_x3y2nw__prog_we_o)
        );
    sbox_se_W i_sbox_x3y2se (
        .bi_x0v1n_L1(_i_sbox_x4y1sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x3y2se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x3y2ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x4y2se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x3y2ne__prog_we_o)
        ,.prog_din(_i_sbox_x3y2ne__prog_dout)
        ,.prog_dout(_i_sbox_x3y2se__prog_dout)
        ,.prog_we_o(_i_sbox_x3y2se__prog_we_o)
        );
    sbox_sw_N i_sbox_x3y2sw (
        .bi_u1v1n_L1(_i_sbox_x3y1sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x3y2sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x2y1nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x3y2se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x2y2__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x3y1nw__prog_we_o)
        ,.prog_din(_i_sbox_x3y1nw__prog_dout)
        ,.prog_dout(_i_sbox_x3y2sw__prog_dout)
        ,.prog_we_o(_i_sbox_x3y2sw__prog_we_o)
        );
    tile_clb i_tile_x3y3 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x3y3__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x3y3__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x3y3sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x2y3ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x3y3sw__prog_we_o)
        ,.prog_din(_i_sbox_x3y3sw__prog_dout)
        ,.prog_dout(_i_tile_x3y3__prog_dout)
        ,.prog_we_o(_i_tile_x3y3__prog_we_o)
        );
    sbox_ne_S i_sbox_x3y3ne (
        .bi_x0y0e_L1(_i_sbox_x3y3nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x3y3ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x3y4ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x4y4se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x3y3__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x3y4se__prog_we_o)
        ,.prog_din(_i_sbox_x3y4se__prog_dout)
        ,.prog_dout(_i_sbox_x3y3ne__prog_dout)
        ,.prog_we_o(_i_sbox_x3y3ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x3y3nw (
        .bi_u1y0n_L1(_i_sbox_x3y3sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x3y3nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x2y3nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x2y4ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x3y3__prog_we_o)
        ,.prog_din(_i_tile_x3y3__prog_dout)
        ,.prog_dout(_i_sbox_x3y3nw__prog_dout)
        ,.prog_we_o(_i_sbox_x3y3nw__prog_we_o)
        );
    sbox_se_W i_sbox_x3y3se (
        .bi_x0v1n_L1(_i_sbox_x4y2sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x3y3se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x3y3ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x4y3se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x3y3ne__prog_we_o)
        ,.prog_din(_i_sbox_x3y3ne__prog_dout)
        ,.prog_dout(_i_sbox_x3y3se__prog_dout)
        ,.prog_we_o(_i_sbox_x3y3se__prog_we_o)
        );
    sbox_sw_N i_sbox_x3y3sw (
        .bi_u1v1n_L1(_i_sbox_x3y2sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x3y3sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x2y2nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x3y3se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x2y3__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x3y2nw__prog_we_o)
        ,.prog_din(_i_sbox_x3y2nw__prog_dout)
        ,.prog_dout(_i_sbox_x3y3sw__prog_dout)
        ,.prog_we_o(_i_sbox_x3y3sw__prog_we_o)
        );
    tile_clb i_tile_x3y4 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x3y4__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x3y4__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x3y4sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x2y4ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x3y4sw__prog_we_o)
        ,.prog_din(_i_sbox_x3y4sw__prog_dout)
        ,.prog_dout(_i_tile_x3y4__prog_dout)
        ,.prog_we_o(_i_tile_x3y4__prog_we_o)
        );
    sbox_ne_S i_sbox_x3y4ne (
        .bi_x0y0e_L1(_i_sbox_x3y4nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x3y4ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x3y5ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x4y5se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x3y4__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x3y5se__prog_we_o)
        ,.prog_din(_i_sbox_x3y5se__prog_dout)
        ,.prog_dout(_i_sbox_x3y4ne__prog_dout)
        ,.prog_we_o(_i_sbox_x3y4ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x3y4nw (
        .bi_u1y0n_L1(_i_sbox_x3y4sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x3y4nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x2y4nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x2y5ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x3y4__prog_we_o)
        ,.prog_din(_i_tile_x3y4__prog_dout)
        ,.prog_dout(_i_sbox_x3y4nw__prog_dout)
        ,.prog_we_o(_i_sbox_x3y4nw__prog_we_o)
        );
    sbox_se_W i_sbox_x3y4se (
        .bi_x0v1n_L1(_i_sbox_x4y3sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x3y4se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x3y4ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x4y4se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x3y4ne__prog_we_o)
        ,.prog_din(_i_sbox_x3y4ne__prog_dout)
        ,.prog_dout(_i_sbox_x3y4se__prog_dout)
        ,.prog_we_o(_i_sbox_x3y4se__prog_we_o)
        );
    sbox_sw_N i_sbox_x3y4sw (
        .bi_u1v1n_L1(_i_sbox_x3y3sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x3y4sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x2y3nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x3y4se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x2y4__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x3y3nw__prog_we_o)
        ,.prog_din(_i_sbox_x3y3nw__prog_dout)
        ,.prog_dout(_i_sbox_x3y4sw__prog_dout)
        ,.prog_we_o(_i_sbox_x3y4sw__prog_we_o)
        );
    tile_clb i_tile_x3y5 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x3y5__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x3y5__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x3y5sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x2y5ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x3y5sw__prog_we_o)
        ,.prog_din(_i_sbox_x3y5sw__prog_dout)
        ,.prog_dout(_i_tile_x3y5__prog_dout)
        ,.prog_we_o(_i_tile_x3y5__prog_we_o)
        );
    sbox_ne_S i_sbox_x3y5ne (
        .bi_x0y0e_L1(_i_sbox_x3y5nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x3y5ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x3y6ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x4y6se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x3y5__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x3y6se__prog_we_o)
        ,.prog_din(_i_sbox_x3y6se__prog_dout)
        ,.prog_dout(_i_sbox_x3y5ne__prog_dout)
        ,.prog_we_o(_i_sbox_x3y5ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x3y5nw (
        .bi_u1y0n_L1(_i_sbox_x3y5sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x3y5nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x2y5nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x2y6ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x3y5__prog_we_o)
        ,.prog_din(_i_tile_x3y5__prog_dout)
        ,.prog_dout(_i_sbox_x3y5nw__prog_dout)
        ,.prog_we_o(_i_sbox_x3y5nw__prog_we_o)
        );
    sbox_se_W i_sbox_x3y5se (
        .bi_x0v1n_L1(_i_sbox_x4y4sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x3y5se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x3y5ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x4y5se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x3y5ne__prog_we_o)
        ,.prog_din(_i_sbox_x3y5ne__prog_dout)
        ,.prog_dout(_i_sbox_x3y5se__prog_dout)
        ,.prog_we_o(_i_sbox_x3y5se__prog_we_o)
        );
    sbox_sw_N i_sbox_x3y5sw (
        .bi_u1v1n_L1(_i_sbox_x3y4sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x3y5sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x2y4nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x3y5se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x2y5__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x3y4nw__prog_we_o)
        ,.prog_din(_i_sbox_x3y4nw__prog_dout)
        ,.prog_dout(_i_sbox_x3y5sw__prog_dout)
        ,.prog_we_o(_i_sbox_x3y5sw__prog_we_o)
        );
    tile_clb i_tile_x3y6 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x3y6__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x3y6__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x3y6sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x2y6ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x3y6sw__prog_we_o)
        ,.prog_din(_i_sbox_x3y6sw__prog_dout)
        ,.prog_dout(_i_tile_x3y6__prog_dout)
        ,.prog_we_o(_i_tile_x3y6__prog_we_o)
        );
    sbox_ne_S i_sbox_x3y6ne (
        .bi_x0y0e_L1(_i_sbox_x3y6nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x3y6ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x3y7ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x4y7se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x3y6__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x3y7se__prog_we_o)
        ,.prog_din(_i_sbox_x3y7se__prog_dout)
        ,.prog_dout(_i_sbox_x3y6ne__prog_dout)
        ,.prog_we_o(_i_sbox_x3y6ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x3y6nw (
        .bi_u1y0n_L1(_i_sbox_x3y6sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x3y6nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x2y6nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x2y7ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x3y6__prog_we_o)
        ,.prog_din(_i_tile_x3y6__prog_dout)
        ,.prog_dout(_i_sbox_x3y6nw__prog_dout)
        ,.prog_we_o(_i_sbox_x3y6nw__prog_we_o)
        );
    sbox_se_W i_sbox_x3y6se (
        .bi_x0v1n_L1(_i_sbox_x4y5sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x3y6se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x3y6ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x4y6se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x3y6ne__prog_we_o)
        ,.prog_din(_i_sbox_x3y6ne__prog_dout)
        ,.prog_dout(_i_sbox_x3y6se__prog_dout)
        ,.prog_we_o(_i_sbox_x3y6se__prog_we_o)
        );
    sbox_sw_N i_sbox_x3y6sw (
        .bi_u1v1n_L1(_i_sbox_x3y5sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x3y6sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x2y5nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x3y6se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x2y6__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x3y5nw__prog_we_o)
        ,.prog_din(_i_sbox_x3y5nw__prog_dout)
        ,.prog_dout(_i_sbox_x3y6sw__prog_dout)
        ,.prog_we_o(_i_sbox_x3y6sw__prog_we_o)
        );
    tile_clb i_tile_x3y7 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x3y7__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x3y7__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x3y7sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x2y7ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x3y7sw__prog_we_o)
        ,.prog_din(_i_sbox_x3y7sw__prog_dout)
        ,.prog_dout(_i_tile_x3y7__prog_dout)
        ,.prog_we_o(_i_tile_x3y7__prog_we_o)
        );
    sbox_ne_S i_sbox_x3y7ne (
        .bi_x0y0e_L1(_i_sbox_x3y7nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x3y7ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x3y8ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x4y8se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x3y7__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x3y8se__prog_we_o)
        ,.prog_din(_i_sbox_x3y8se__prog_dout)
        ,.prog_dout(_i_sbox_x3y7ne__prog_dout)
        ,.prog_we_o(_i_sbox_x3y7ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x3y7nw (
        .bi_u1y0n_L1(_i_sbox_x3y7sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x3y7nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x2y7nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x2y8ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x3y7__prog_we_o)
        ,.prog_din(_i_tile_x3y7__prog_dout)
        ,.prog_dout(_i_sbox_x3y7nw__prog_dout)
        ,.prog_we_o(_i_sbox_x3y7nw__prog_we_o)
        );
    sbox_se_W i_sbox_x3y7se (
        .bi_x0v1n_L1(_i_sbox_x4y6sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x3y7se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x3y7ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x4y7se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x3y7ne__prog_we_o)
        ,.prog_din(_i_sbox_x3y7ne__prog_dout)
        ,.prog_dout(_i_sbox_x3y7se__prog_dout)
        ,.prog_we_o(_i_sbox_x3y7se__prog_we_o)
        );
    sbox_sw_N i_sbox_x3y7sw (
        .bi_u1v1n_L1(_i_sbox_x3y6sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x3y7sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x2y6nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x3y7se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x2y7__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x3y6nw__prog_we_o)
        ,.prog_din(_i_sbox_x3y6nw__prog_dout)
        ,.prog_dout(_i_sbox_x3y7sw__prog_dout)
        ,.prog_we_o(_i_sbox_x3y7sw__prog_we_o)
        );
    tile_clb i_tile_x3y8 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x3y8__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x3y8__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x3y8sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x2y8ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x3y8sw__prog_we_o)
        ,.prog_din(_i_sbox_x3y8sw__prog_dout)
        ,.prog_dout(_i_tile_x3y8__prog_dout)
        ,.prog_we_o(_i_tile_x3y8__prog_we_o)
        );
    sbox_ne_S_ex_s i_sbox_x3y8ne (
        .bi_x0y0e_L1(_i_sbox_x3y8nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x3y8ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x4y9se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x3y8__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x3y9se__prog_we_o)
        ,.prog_din(_i_sbox_x3y9se__prog_dout)
        ,.prog_dout(_i_sbox_x3y8ne__prog_dout)
        ,.prog_we_o(_i_sbox_x3y8ne__prog_we_o)
        );
    sbox_nw_E_ex_s i_sbox_x3y8nw (
        .bi_u1y0n_L1(_i_sbox_x3y8sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x3y8nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x2y8nw__so_x0y0e_L1)
        ,.cu_x0y0e_L1(_i_tile_x3y9__cu_x0v1e_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x3y8__prog_we_o)
        ,.prog_din(_i_tile_x3y8__prog_dout)
        ,.prog_dout(_i_sbox_x3y8nw__prog_dout)
        ,.prog_we_o(_i_sbox_x3y8nw__prog_we_o)
        );
    sbox_se_W i_sbox_x3y8se (
        .bi_x0v1n_L1(_i_sbox_x4y7sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x3y8se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x3y8ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x4y8se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x3y8ne__prog_we_o)
        ,.prog_din(_i_sbox_x3y8ne__prog_dout)
        ,.prog_dout(_i_sbox_x3y8se__prog_dout)
        ,.prog_we_o(_i_sbox_x3y8se__prog_we_o)
        );
    sbox_sw_N i_sbox_x3y8sw (
        .bi_u1v1n_L1(_i_sbox_x3y7sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x3y8sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x2y7nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x3y8se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x2y8__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x3y7nw__prog_we_o)
        ,.prog_din(_i_sbox_x3y7nw__prog_dout)
        ,.prog_dout(_i_sbox_x3y8sw__prog_dout)
        ,.prog_we_o(_i_sbox_x3y8sw__prog_we_o)
        );
    t_io_n i_tile_x3y9 (
        .bi_x0v1e_L1(_i_sbox_x3y8nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x3y9se__so_x0v1w_L1)
        ,.cu_x0v1e_L1(_i_tile_x3y9__cu_x0v1e_L1)
        ,.cu_x0v1w_L1(_i_tile_x3y9__cu_x0v1w_L1)
        ,.ipin_x0y0_0(ipin_x3y9_0)
        ,.opin_x0y0_0(_i_tile_x3y9__opin_x0y0_0)
        ,.oe_x0y0_0(_i_tile_x3y9__oe_x0y0_0)
        ,.ipin_x0y0_1(ipin_x3y9_1)
        ,.opin_x0y0_1(_i_tile_x3y9__opin_x0y0_1)
        ,.oe_x0y0_1(_i_tile_x3y9__oe_x0y0_1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x3y8nw__prog_we_o)
        ,.prog_din(_i_sbox_x3y8nw__prog_dout)
        ,.prog_dout(_i_tile_x3y9__prog_dout)
        ,.prog_we_o(_i_tile_x3y9__prog_we_o)
        );
    sbox_se_W_ex_s i_sbox_x3y9se (
        .bi_x0v1n_L1(_i_sbox_x4y8sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x3y9se__so_x0v1w_L1)
        ,.bi_x1v1w_L1(_i_sbox_x4y9se__so_x0v1w_L1)
        ,.cu_x0v1w_L1(_i_tile_x3y9__cu_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x3y9__prog_we_o)
        ,.prog_din(_i_tile_x3y9__prog_dout)
        ,.prog_dout(_i_sbox_x3y9se__prog_dout)
        ,.prog_we_o(_i_sbox_x3y9se__prog_we_o)
        );
    sbox_sw_s_ex_s i_sbox_x3y9sw (
        .bi_u1v1e_L1(_i_sbox_x2y8nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x3y9se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_ne_n_ex_n i_sbox_x4y0ne (
        .bi_x0y0e_L1(_i_sbox_x4y0nw__so_x0y0e_L1)
        ,.bi_x1y0w_L1(_i_sbox_x5y1se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_nw_E_ex_n i_sbox_x4y0nw (
        .bi_u1y0e_L1(_i_sbox_x3y0nw__so_x0y0e_L1)
        ,.so_x0y0e_L1(_i_sbox_x4y0nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x3y1ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x3y1se__prog_we_o)
        ,.prog_din(_i_sbox_x3y1se__prog_dout)
        ,.prog_dout(_i_sbox_x4y0nw__prog_dout)
        ,.prog_we_o(_i_sbox_x4y0nw__prog_we_o)
        );
    tile_clb i_tile_x4y1 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x4y1__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x4y1__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x4y1sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x3y1ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x4y1sw__prog_we_o)
        ,.prog_din(_i_sbox_x4y1sw__prog_dout)
        ,.prog_dout(_i_tile_x4y1__prog_dout)
        ,.prog_we_o(_i_tile_x4y1__prog_we_o)
        );
    sbox_ne_S i_sbox_x4y1ne (
        .bi_x0y0e_L1(_i_sbox_x4y1nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x4y1ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x4y2ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x5y2se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x4y1__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x4y2se__prog_we_o)
        ,.prog_din(_i_sbox_x4y2se__prog_dout)
        ,.prog_dout(_i_sbox_x4y1ne__prog_dout)
        ,.prog_we_o(_i_sbox_x4y1ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x4y1nw (
        .bi_u1y0n_L1(_i_sbox_x4y1sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x4y1nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x3y1nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x3y2ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x4y1__prog_we_o)
        ,.prog_din(_i_tile_x4y1__prog_dout)
        ,.prog_dout(_i_sbox_x4y1nw__prog_dout)
        ,.prog_we_o(_i_sbox_x4y1nw__prog_we_o)
        );
    sbox_se_W_ex_n i_sbox_x4y1se (
        .bi_x0y0s_L1(_i_sbox_x4y1ne__so_x0y0s_L1)
        ,.so_x0v1w_L1(_i_sbox_x4y1se__so_x0v1w_L1)
        ,.bi_x1v1w_L1(_i_sbox_x5y1se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x4y1ne__prog_we_o)
        ,.prog_din(_i_sbox_x4y1ne__prog_dout)
        ,.prog_dout(_i_sbox_x4y1se__prog_dout)
        ,.prog_we_o(_i_sbox_x4y1se__prog_we_o)
        );
    sbox_sw_N_ex_n i_sbox_x4y1sw (
        .bi_u1v1e_L1(_i_sbox_x3y0nw__so_x0y0e_L1)
        ,.so_u1y0n_L1(_i_sbox_x4y1sw__so_u1y0n_L1)
        ,.bi_x0v1w_L1(_i_sbox_x4y1se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x3y1__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x4y0nw__prog_we_o)
        ,.prog_din(_i_sbox_x4y0nw__prog_dout)
        ,.prog_dout(_i_sbox_x4y1sw__prog_dout)
        ,.prog_we_o(_i_sbox_x4y1sw__prog_we_o)
        );
    tile_clb i_tile_x4y2 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x4y2__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x4y2__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x4y2sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x3y2ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x4y2sw__prog_we_o)
        ,.prog_din(_i_sbox_x4y2sw__prog_dout)
        ,.prog_dout(_i_tile_x4y2__prog_dout)
        ,.prog_we_o(_i_tile_x4y2__prog_we_o)
        );
    sbox_ne_S i_sbox_x4y2ne (
        .bi_x0y0e_L1(_i_sbox_x4y2nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x4y2ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x4y3ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x5y3se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x4y2__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x4y3se__prog_we_o)
        ,.prog_din(_i_sbox_x4y3se__prog_dout)
        ,.prog_dout(_i_sbox_x4y2ne__prog_dout)
        ,.prog_we_o(_i_sbox_x4y2ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x4y2nw (
        .bi_u1y0n_L1(_i_sbox_x4y2sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x4y2nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x3y2nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x3y3ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x4y2__prog_we_o)
        ,.prog_din(_i_tile_x4y2__prog_dout)
        ,.prog_dout(_i_sbox_x4y2nw__prog_dout)
        ,.prog_we_o(_i_sbox_x4y2nw__prog_we_o)
        );
    sbox_se_W i_sbox_x4y2se (
        .bi_x0v1n_L1(_i_sbox_x5y1sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x4y2se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x4y2ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x5y2se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x4y2ne__prog_we_o)
        ,.prog_din(_i_sbox_x4y2ne__prog_dout)
        ,.prog_dout(_i_sbox_x4y2se__prog_dout)
        ,.prog_we_o(_i_sbox_x4y2se__prog_we_o)
        );
    sbox_sw_N i_sbox_x4y2sw (
        .bi_u1v1n_L1(_i_sbox_x4y1sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x4y2sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x3y1nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x4y2se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x3y2__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x4y1nw__prog_we_o)
        ,.prog_din(_i_sbox_x4y1nw__prog_dout)
        ,.prog_dout(_i_sbox_x4y2sw__prog_dout)
        ,.prog_we_o(_i_sbox_x4y2sw__prog_we_o)
        );
    tile_clb i_tile_x4y3 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x4y3__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x4y3__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x4y3sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x3y3ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x4y3sw__prog_we_o)
        ,.prog_din(_i_sbox_x4y3sw__prog_dout)
        ,.prog_dout(_i_tile_x4y3__prog_dout)
        ,.prog_we_o(_i_tile_x4y3__prog_we_o)
        );
    sbox_ne_S i_sbox_x4y3ne (
        .bi_x0y0e_L1(_i_sbox_x4y3nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x4y3ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x4y4ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x5y4se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x4y3__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x4y4se__prog_we_o)
        ,.prog_din(_i_sbox_x4y4se__prog_dout)
        ,.prog_dout(_i_sbox_x4y3ne__prog_dout)
        ,.prog_we_o(_i_sbox_x4y3ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x4y3nw (
        .bi_u1y0n_L1(_i_sbox_x4y3sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x4y3nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x3y3nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x3y4ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x4y3__prog_we_o)
        ,.prog_din(_i_tile_x4y3__prog_dout)
        ,.prog_dout(_i_sbox_x4y3nw__prog_dout)
        ,.prog_we_o(_i_sbox_x4y3nw__prog_we_o)
        );
    sbox_se_W i_sbox_x4y3se (
        .bi_x0v1n_L1(_i_sbox_x5y2sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x4y3se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x4y3ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x5y3se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x4y3ne__prog_we_o)
        ,.prog_din(_i_sbox_x4y3ne__prog_dout)
        ,.prog_dout(_i_sbox_x4y3se__prog_dout)
        ,.prog_we_o(_i_sbox_x4y3se__prog_we_o)
        );
    sbox_sw_N i_sbox_x4y3sw (
        .bi_u1v1n_L1(_i_sbox_x4y2sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x4y3sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x3y2nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x4y3se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x3y3__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x4y2nw__prog_we_o)
        ,.prog_din(_i_sbox_x4y2nw__prog_dout)
        ,.prog_dout(_i_sbox_x4y3sw__prog_dout)
        ,.prog_we_o(_i_sbox_x4y3sw__prog_we_o)
        );
    tile_clb i_tile_x4y4 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x4y4__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x4y4__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x4y4sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x3y4ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x4y4sw__prog_we_o)
        ,.prog_din(_i_sbox_x4y4sw__prog_dout)
        ,.prog_dout(_i_tile_x4y4__prog_dout)
        ,.prog_we_o(_i_tile_x4y4__prog_we_o)
        );
    sbox_ne_S i_sbox_x4y4ne (
        .bi_x0y0e_L1(_i_sbox_x4y4nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x4y4ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x4y5ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x5y5se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x4y4__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x4y5se__prog_we_o)
        ,.prog_din(_i_sbox_x4y5se__prog_dout)
        ,.prog_dout(_i_sbox_x4y4ne__prog_dout)
        ,.prog_we_o(_i_sbox_x4y4ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x4y4nw (
        .bi_u1y0n_L1(_i_sbox_x4y4sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x4y4nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x3y4nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x3y5ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x4y4__prog_we_o)
        ,.prog_din(_i_tile_x4y4__prog_dout)
        ,.prog_dout(_i_sbox_x4y4nw__prog_dout)
        ,.prog_we_o(_i_sbox_x4y4nw__prog_we_o)
        );
    sbox_se_W i_sbox_x4y4se (
        .bi_x0v1n_L1(_i_sbox_x5y3sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x4y4se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x4y4ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x5y4se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x4y4ne__prog_we_o)
        ,.prog_din(_i_sbox_x4y4ne__prog_dout)
        ,.prog_dout(_i_sbox_x4y4se__prog_dout)
        ,.prog_we_o(_i_sbox_x4y4se__prog_we_o)
        );
    sbox_sw_N i_sbox_x4y4sw (
        .bi_u1v1n_L1(_i_sbox_x4y3sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x4y4sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x3y3nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x4y4se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x3y4__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x4y3nw__prog_we_o)
        ,.prog_din(_i_sbox_x4y3nw__prog_dout)
        ,.prog_dout(_i_sbox_x4y4sw__prog_dout)
        ,.prog_we_o(_i_sbox_x4y4sw__prog_we_o)
        );
    tile_clb i_tile_x4y5 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x4y5__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x4y5__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x4y5sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x3y5ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x4y5sw__prog_we_o)
        ,.prog_din(_i_sbox_x4y5sw__prog_dout)
        ,.prog_dout(_i_tile_x4y5__prog_dout)
        ,.prog_we_o(_i_tile_x4y5__prog_we_o)
        );
    sbox_ne_S i_sbox_x4y5ne (
        .bi_x0y0e_L1(_i_sbox_x4y5nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x4y5ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x4y6ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x5y6se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x4y5__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x4y6se__prog_we_o)
        ,.prog_din(_i_sbox_x4y6se__prog_dout)
        ,.prog_dout(_i_sbox_x4y5ne__prog_dout)
        ,.prog_we_o(_i_sbox_x4y5ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x4y5nw (
        .bi_u1y0n_L1(_i_sbox_x4y5sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x4y5nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x3y5nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x3y6ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x4y5__prog_we_o)
        ,.prog_din(_i_tile_x4y5__prog_dout)
        ,.prog_dout(_i_sbox_x4y5nw__prog_dout)
        ,.prog_we_o(_i_sbox_x4y5nw__prog_we_o)
        );
    sbox_se_W i_sbox_x4y5se (
        .bi_x0v1n_L1(_i_sbox_x5y4sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x4y5se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x4y5ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x5y5se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x4y5ne__prog_we_o)
        ,.prog_din(_i_sbox_x4y5ne__prog_dout)
        ,.prog_dout(_i_sbox_x4y5se__prog_dout)
        ,.prog_we_o(_i_sbox_x4y5se__prog_we_o)
        );
    sbox_sw_N i_sbox_x4y5sw (
        .bi_u1v1n_L1(_i_sbox_x4y4sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x4y5sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x3y4nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x4y5se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x3y5__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x4y4nw__prog_we_o)
        ,.prog_din(_i_sbox_x4y4nw__prog_dout)
        ,.prog_dout(_i_sbox_x4y5sw__prog_dout)
        ,.prog_we_o(_i_sbox_x4y5sw__prog_we_o)
        );
    tile_clb i_tile_x4y6 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x4y6__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x4y6__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x4y6sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x3y6ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x4y6sw__prog_we_o)
        ,.prog_din(_i_sbox_x4y6sw__prog_dout)
        ,.prog_dout(_i_tile_x4y6__prog_dout)
        ,.prog_we_o(_i_tile_x4y6__prog_we_o)
        );
    sbox_ne_S i_sbox_x4y6ne (
        .bi_x0y0e_L1(_i_sbox_x4y6nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x4y6ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x4y7ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x5y7se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x4y6__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x4y7se__prog_we_o)
        ,.prog_din(_i_sbox_x4y7se__prog_dout)
        ,.prog_dout(_i_sbox_x4y6ne__prog_dout)
        ,.prog_we_o(_i_sbox_x4y6ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x4y6nw (
        .bi_u1y0n_L1(_i_sbox_x4y6sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x4y6nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x3y6nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x3y7ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x4y6__prog_we_o)
        ,.prog_din(_i_tile_x4y6__prog_dout)
        ,.prog_dout(_i_sbox_x4y6nw__prog_dout)
        ,.prog_we_o(_i_sbox_x4y6nw__prog_we_o)
        );
    sbox_se_W i_sbox_x4y6se (
        .bi_x0v1n_L1(_i_sbox_x5y5sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x4y6se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x4y6ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x5y6se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x4y6ne__prog_we_o)
        ,.prog_din(_i_sbox_x4y6ne__prog_dout)
        ,.prog_dout(_i_sbox_x4y6se__prog_dout)
        ,.prog_we_o(_i_sbox_x4y6se__prog_we_o)
        );
    sbox_sw_N i_sbox_x4y6sw (
        .bi_u1v1n_L1(_i_sbox_x4y5sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x4y6sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x3y5nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x4y6se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x3y6__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x4y5nw__prog_we_o)
        ,.prog_din(_i_sbox_x4y5nw__prog_dout)
        ,.prog_dout(_i_sbox_x4y6sw__prog_dout)
        ,.prog_we_o(_i_sbox_x4y6sw__prog_we_o)
        );
    tile_clb i_tile_x4y7 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x4y7__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x4y7__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x4y7sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x3y7ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x4y7sw__prog_we_o)
        ,.prog_din(_i_sbox_x4y7sw__prog_dout)
        ,.prog_dout(_i_tile_x4y7__prog_dout)
        ,.prog_we_o(_i_tile_x4y7__prog_we_o)
        );
    sbox_ne_S i_sbox_x4y7ne (
        .bi_x0y0e_L1(_i_sbox_x4y7nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x4y7ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x4y8ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x5y8se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x4y7__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x4y8se__prog_we_o)
        ,.prog_din(_i_sbox_x4y8se__prog_dout)
        ,.prog_dout(_i_sbox_x4y7ne__prog_dout)
        ,.prog_we_o(_i_sbox_x4y7ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x4y7nw (
        .bi_u1y0n_L1(_i_sbox_x4y7sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x4y7nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x3y7nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x3y8ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x4y7__prog_we_o)
        ,.prog_din(_i_tile_x4y7__prog_dout)
        ,.prog_dout(_i_sbox_x4y7nw__prog_dout)
        ,.prog_we_o(_i_sbox_x4y7nw__prog_we_o)
        );
    sbox_se_W i_sbox_x4y7se (
        .bi_x0v1n_L1(_i_sbox_x5y6sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x4y7se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x4y7ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x5y7se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x4y7ne__prog_we_o)
        ,.prog_din(_i_sbox_x4y7ne__prog_dout)
        ,.prog_dout(_i_sbox_x4y7se__prog_dout)
        ,.prog_we_o(_i_sbox_x4y7se__prog_we_o)
        );
    sbox_sw_N i_sbox_x4y7sw (
        .bi_u1v1n_L1(_i_sbox_x4y6sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x4y7sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x3y6nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x4y7se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x3y7__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x4y6nw__prog_we_o)
        ,.prog_din(_i_sbox_x4y6nw__prog_dout)
        ,.prog_dout(_i_sbox_x4y7sw__prog_dout)
        ,.prog_we_o(_i_sbox_x4y7sw__prog_we_o)
        );
    tile_clb i_tile_x4y8 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x4y8__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x4y8__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x4y8sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x3y8ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x4y8sw__prog_we_o)
        ,.prog_din(_i_sbox_x4y8sw__prog_dout)
        ,.prog_dout(_i_tile_x4y8__prog_dout)
        ,.prog_we_o(_i_tile_x4y8__prog_we_o)
        );
    sbox_ne_S_ex_s i_sbox_x4y8ne (
        .bi_x0y0e_L1(_i_sbox_x4y8nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x4y8ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x5y9se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x4y8__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x4y9se__prog_we_o)
        ,.prog_din(_i_sbox_x4y9se__prog_dout)
        ,.prog_dout(_i_sbox_x4y8ne__prog_dout)
        ,.prog_we_o(_i_sbox_x4y8ne__prog_we_o)
        );
    sbox_nw_E_ex_s i_sbox_x4y8nw (
        .bi_u1y0n_L1(_i_sbox_x4y8sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x4y8nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x3y8nw__so_x0y0e_L1)
        ,.cu_x0y0e_L1(_i_tile_x4y9__cu_x0v1e_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x4y8__prog_we_o)
        ,.prog_din(_i_tile_x4y8__prog_dout)
        ,.prog_dout(_i_sbox_x4y8nw__prog_dout)
        ,.prog_we_o(_i_sbox_x4y8nw__prog_we_o)
        );
    sbox_se_W i_sbox_x4y8se (
        .bi_x0v1n_L1(_i_sbox_x5y7sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x4y8se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x4y8ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x5y8se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x4y8ne__prog_we_o)
        ,.prog_din(_i_sbox_x4y8ne__prog_dout)
        ,.prog_dout(_i_sbox_x4y8se__prog_dout)
        ,.prog_we_o(_i_sbox_x4y8se__prog_we_o)
        );
    sbox_sw_N i_sbox_x4y8sw (
        .bi_u1v1n_L1(_i_sbox_x4y7sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x4y8sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x3y7nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x4y8se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x3y8__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x4y7nw__prog_we_o)
        ,.prog_din(_i_sbox_x4y7nw__prog_dout)
        ,.prog_dout(_i_sbox_x4y8sw__prog_dout)
        ,.prog_we_o(_i_sbox_x4y8sw__prog_we_o)
        );
    t_io_n i_tile_x4y9 (
        .bi_x0v1e_L1(_i_sbox_x4y8nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x4y9se__so_x0v1w_L1)
        ,.cu_x0v1e_L1(_i_tile_x4y9__cu_x0v1e_L1)
        ,.cu_x0v1w_L1(_i_tile_x4y9__cu_x0v1w_L1)
        ,.ipin_x0y0_0(ipin_x4y9_0)
        ,.opin_x0y0_0(_i_tile_x4y9__opin_x0y0_0)
        ,.oe_x0y0_0(_i_tile_x4y9__oe_x0y0_0)
        ,.ipin_x0y0_1(ipin_x4y9_1)
        ,.opin_x0y0_1(_i_tile_x4y9__opin_x0y0_1)
        ,.oe_x0y0_1(_i_tile_x4y9__oe_x0y0_1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x4y8nw__prog_we_o)
        ,.prog_din(_i_sbox_x4y8nw__prog_dout)
        ,.prog_dout(_i_tile_x4y9__prog_dout)
        ,.prog_we_o(_i_tile_x4y9__prog_we_o)
        );
    sbox_se_W_ex_s i_sbox_x4y9se (
        .bi_x0v1n_L1(_i_sbox_x5y8sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x4y9se__so_x0v1w_L1)
        ,.bi_x1v1w_L1(_i_sbox_x5y9se__so_x0v1w_L1)
        ,.cu_x0v1w_L1(_i_tile_x4y9__cu_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x4y9__prog_we_o)
        ,.prog_din(_i_tile_x4y9__prog_dout)
        ,.prog_dout(_i_sbox_x4y9se__prog_dout)
        ,.prog_we_o(_i_sbox_x4y9se__prog_we_o)
        );
    sbox_sw_s_ex_s i_sbox_x4y9sw (
        .bi_u1v1e_L1(_i_sbox_x3y8nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x4y9se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_ne_n_ex_n i_sbox_x5y0ne (
        .bi_x0y0e_L1(_i_sbox_x5y0nw__so_x0y0e_L1)
        ,.bi_x1y0w_L1(_i_sbox_x6y1se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_nw_E_ex_n i_sbox_x5y0nw (
        .bi_u1y0e_L1(_i_sbox_x4y0nw__so_x0y0e_L1)
        ,.so_x0y0e_L1(_i_sbox_x5y0nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x4y1ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x4y1se__prog_we_o)
        ,.prog_din(_i_sbox_x4y1se__prog_dout)
        ,.prog_dout(_i_sbox_x5y0nw__prog_dout)
        ,.prog_we_o(_i_sbox_x5y0nw__prog_we_o)
        );
    tile_clb i_tile_x5y1 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x5y1__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x5y1__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x5y1sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x4y1ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x5y1sw__prog_we_o)
        ,.prog_din(_i_sbox_x5y1sw__prog_dout)
        ,.prog_dout(_i_tile_x5y1__prog_dout)
        ,.prog_we_o(_i_tile_x5y1__prog_we_o)
        );
    sbox_ne_S i_sbox_x5y1ne (
        .bi_x0y0e_L1(_i_sbox_x5y1nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x5y1ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x5y2ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x6y2se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x5y1__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x5y2se__prog_we_o)
        ,.prog_din(_i_sbox_x5y2se__prog_dout)
        ,.prog_dout(_i_sbox_x5y1ne__prog_dout)
        ,.prog_we_o(_i_sbox_x5y1ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x5y1nw (
        .bi_u1y0n_L1(_i_sbox_x5y1sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x5y1nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x4y1nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x4y2ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x5y1__prog_we_o)
        ,.prog_din(_i_tile_x5y1__prog_dout)
        ,.prog_dout(_i_sbox_x5y1nw__prog_dout)
        ,.prog_we_o(_i_sbox_x5y1nw__prog_we_o)
        );
    sbox_se_W_ex_n i_sbox_x5y1se (
        .bi_x0y0s_L1(_i_sbox_x5y1ne__so_x0y0s_L1)
        ,.so_x0v1w_L1(_i_sbox_x5y1se__so_x0v1w_L1)
        ,.bi_x1v1w_L1(_i_sbox_x6y1se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x5y1ne__prog_we_o)
        ,.prog_din(_i_sbox_x5y1ne__prog_dout)
        ,.prog_dout(_i_sbox_x5y1se__prog_dout)
        ,.prog_we_o(_i_sbox_x5y1se__prog_we_o)
        );
    sbox_sw_N_ex_n i_sbox_x5y1sw (
        .bi_u1v1e_L1(_i_sbox_x4y0nw__so_x0y0e_L1)
        ,.so_u1y0n_L1(_i_sbox_x5y1sw__so_u1y0n_L1)
        ,.bi_x0v1w_L1(_i_sbox_x5y1se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x4y1__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x5y0nw__prog_we_o)
        ,.prog_din(_i_sbox_x5y0nw__prog_dout)
        ,.prog_dout(_i_sbox_x5y1sw__prog_dout)
        ,.prog_we_o(_i_sbox_x5y1sw__prog_we_o)
        );
    tile_clb i_tile_x5y2 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x5y2__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x5y2__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x5y2sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x4y2ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x5y2sw__prog_we_o)
        ,.prog_din(_i_sbox_x5y2sw__prog_dout)
        ,.prog_dout(_i_tile_x5y2__prog_dout)
        ,.prog_we_o(_i_tile_x5y2__prog_we_o)
        );
    sbox_ne_S i_sbox_x5y2ne (
        .bi_x0y0e_L1(_i_sbox_x5y2nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x5y2ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x5y3ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x6y3se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x5y2__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x5y3se__prog_we_o)
        ,.prog_din(_i_sbox_x5y3se__prog_dout)
        ,.prog_dout(_i_sbox_x5y2ne__prog_dout)
        ,.prog_we_o(_i_sbox_x5y2ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x5y2nw (
        .bi_u1y0n_L1(_i_sbox_x5y2sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x5y2nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x4y2nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x4y3ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x5y2__prog_we_o)
        ,.prog_din(_i_tile_x5y2__prog_dout)
        ,.prog_dout(_i_sbox_x5y2nw__prog_dout)
        ,.prog_we_o(_i_sbox_x5y2nw__prog_we_o)
        );
    sbox_se_W i_sbox_x5y2se (
        .bi_x0v1n_L1(_i_sbox_x6y1sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x5y2se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x5y2ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x6y2se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x5y2ne__prog_we_o)
        ,.prog_din(_i_sbox_x5y2ne__prog_dout)
        ,.prog_dout(_i_sbox_x5y2se__prog_dout)
        ,.prog_we_o(_i_sbox_x5y2se__prog_we_o)
        );
    sbox_sw_N i_sbox_x5y2sw (
        .bi_u1v1n_L1(_i_sbox_x5y1sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x5y2sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x4y1nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x5y2se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x4y2__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x5y1nw__prog_we_o)
        ,.prog_din(_i_sbox_x5y1nw__prog_dout)
        ,.prog_dout(_i_sbox_x5y2sw__prog_dout)
        ,.prog_we_o(_i_sbox_x5y2sw__prog_we_o)
        );
    tile_clb i_tile_x5y3 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x5y3__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x5y3__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x5y3sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x4y3ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x5y3sw__prog_we_o)
        ,.prog_din(_i_sbox_x5y3sw__prog_dout)
        ,.prog_dout(_i_tile_x5y3__prog_dout)
        ,.prog_we_o(_i_tile_x5y3__prog_we_o)
        );
    sbox_ne_S i_sbox_x5y3ne (
        .bi_x0y0e_L1(_i_sbox_x5y3nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x5y3ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x5y4ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x6y4se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x5y3__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x5y4se__prog_we_o)
        ,.prog_din(_i_sbox_x5y4se__prog_dout)
        ,.prog_dout(_i_sbox_x5y3ne__prog_dout)
        ,.prog_we_o(_i_sbox_x5y3ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x5y3nw (
        .bi_u1y0n_L1(_i_sbox_x5y3sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x5y3nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x4y3nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x4y4ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x5y3__prog_we_o)
        ,.prog_din(_i_tile_x5y3__prog_dout)
        ,.prog_dout(_i_sbox_x5y3nw__prog_dout)
        ,.prog_we_o(_i_sbox_x5y3nw__prog_we_o)
        );
    sbox_se_W i_sbox_x5y3se (
        .bi_x0v1n_L1(_i_sbox_x6y2sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x5y3se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x5y3ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x6y3se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x5y3ne__prog_we_o)
        ,.prog_din(_i_sbox_x5y3ne__prog_dout)
        ,.prog_dout(_i_sbox_x5y3se__prog_dout)
        ,.prog_we_o(_i_sbox_x5y3se__prog_we_o)
        );
    sbox_sw_N i_sbox_x5y3sw (
        .bi_u1v1n_L1(_i_sbox_x5y2sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x5y3sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x4y2nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x5y3se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x4y3__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x5y2nw__prog_we_o)
        ,.prog_din(_i_sbox_x5y2nw__prog_dout)
        ,.prog_dout(_i_sbox_x5y3sw__prog_dout)
        ,.prog_we_o(_i_sbox_x5y3sw__prog_we_o)
        );
    tile_clb i_tile_x5y4 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x5y4__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x5y4__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x5y4sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x4y4ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x5y4sw__prog_we_o)
        ,.prog_din(_i_sbox_x5y4sw__prog_dout)
        ,.prog_dout(_i_tile_x5y4__prog_dout)
        ,.prog_we_o(_i_tile_x5y4__prog_we_o)
        );
    sbox_ne_S i_sbox_x5y4ne (
        .bi_x0y0e_L1(_i_sbox_x5y4nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x5y4ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x5y5ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x6y5se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x5y4__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x5y5se__prog_we_o)
        ,.prog_din(_i_sbox_x5y5se__prog_dout)
        ,.prog_dout(_i_sbox_x5y4ne__prog_dout)
        ,.prog_we_o(_i_sbox_x5y4ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x5y4nw (
        .bi_u1y0n_L1(_i_sbox_x5y4sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x5y4nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x4y4nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x4y5ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x5y4__prog_we_o)
        ,.prog_din(_i_tile_x5y4__prog_dout)
        ,.prog_dout(_i_sbox_x5y4nw__prog_dout)
        ,.prog_we_o(_i_sbox_x5y4nw__prog_we_o)
        );
    sbox_se_W i_sbox_x5y4se (
        .bi_x0v1n_L1(_i_sbox_x6y3sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x5y4se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x5y4ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x6y4se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x5y4ne__prog_we_o)
        ,.prog_din(_i_sbox_x5y4ne__prog_dout)
        ,.prog_dout(_i_sbox_x5y4se__prog_dout)
        ,.prog_we_o(_i_sbox_x5y4se__prog_we_o)
        );
    sbox_sw_N i_sbox_x5y4sw (
        .bi_u1v1n_L1(_i_sbox_x5y3sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x5y4sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x4y3nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x5y4se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x4y4__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x5y3nw__prog_we_o)
        ,.prog_din(_i_sbox_x5y3nw__prog_dout)
        ,.prog_dout(_i_sbox_x5y4sw__prog_dout)
        ,.prog_we_o(_i_sbox_x5y4sw__prog_we_o)
        );
    tile_clb i_tile_x5y5 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x5y5__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x5y5__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x5y5sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x4y5ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x5y5sw__prog_we_o)
        ,.prog_din(_i_sbox_x5y5sw__prog_dout)
        ,.prog_dout(_i_tile_x5y5__prog_dout)
        ,.prog_we_o(_i_tile_x5y5__prog_we_o)
        );
    sbox_ne_S i_sbox_x5y5ne (
        .bi_x0y0e_L1(_i_sbox_x5y5nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x5y5ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x5y6ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x6y6se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x5y5__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x5y6se__prog_we_o)
        ,.prog_din(_i_sbox_x5y6se__prog_dout)
        ,.prog_dout(_i_sbox_x5y5ne__prog_dout)
        ,.prog_we_o(_i_sbox_x5y5ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x5y5nw (
        .bi_u1y0n_L1(_i_sbox_x5y5sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x5y5nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x4y5nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x4y6ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x5y5__prog_we_o)
        ,.prog_din(_i_tile_x5y5__prog_dout)
        ,.prog_dout(_i_sbox_x5y5nw__prog_dout)
        ,.prog_we_o(_i_sbox_x5y5nw__prog_we_o)
        );
    sbox_se_W i_sbox_x5y5se (
        .bi_x0v1n_L1(_i_sbox_x6y4sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x5y5se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x5y5ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x6y5se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x5y5ne__prog_we_o)
        ,.prog_din(_i_sbox_x5y5ne__prog_dout)
        ,.prog_dout(_i_sbox_x5y5se__prog_dout)
        ,.prog_we_o(_i_sbox_x5y5se__prog_we_o)
        );
    sbox_sw_N i_sbox_x5y5sw (
        .bi_u1v1n_L1(_i_sbox_x5y4sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x5y5sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x4y4nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x5y5se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x4y5__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x5y4nw__prog_we_o)
        ,.prog_din(_i_sbox_x5y4nw__prog_dout)
        ,.prog_dout(_i_sbox_x5y5sw__prog_dout)
        ,.prog_we_o(_i_sbox_x5y5sw__prog_we_o)
        );
    tile_clb i_tile_x5y6 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x5y6__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x5y6__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x5y6sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x4y6ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x5y6sw__prog_we_o)
        ,.prog_din(_i_sbox_x5y6sw__prog_dout)
        ,.prog_dout(_i_tile_x5y6__prog_dout)
        ,.prog_we_o(_i_tile_x5y6__prog_we_o)
        );
    sbox_ne_S i_sbox_x5y6ne (
        .bi_x0y0e_L1(_i_sbox_x5y6nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x5y6ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x5y7ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x6y7se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x5y6__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x5y7se__prog_we_o)
        ,.prog_din(_i_sbox_x5y7se__prog_dout)
        ,.prog_dout(_i_sbox_x5y6ne__prog_dout)
        ,.prog_we_o(_i_sbox_x5y6ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x5y6nw (
        .bi_u1y0n_L1(_i_sbox_x5y6sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x5y6nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x4y6nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x4y7ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x5y6__prog_we_o)
        ,.prog_din(_i_tile_x5y6__prog_dout)
        ,.prog_dout(_i_sbox_x5y6nw__prog_dout)
        ,.prog_we_o(_i_sbox_x5y6nw__prog_we_o)
        );
    sbox_se_W i_sbox_x5y6se (
        .bi_x0v1n_L1(_i_sbox_x6y5sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x5y6se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x5y6ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x6y6se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x5y6ne__prog_we_o)
        ,.prog_din(_i_sbox_x5y6ne__prog_dout)
        ,.prog_dout(_i_sbox_x5y6se__prog_dout)
        ,.prog_we_o(_i_sbox_x5y6se__prog_we_o)
        );
    sbox_sw_N i_sbox_x5y6sw (
        .bi_u1v1n_L1(_i_sbox_x5y5sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x5y6sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x4y5nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x5y6se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x4y6__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x5y5nw__prog_we_o)
        ,.prog_din(_i_sbox_x5y5nw__prog_dout)
        ,.prog_dout(_i_sbox_x5y6sw__prog_dout)
        ,.prog_we_o(_i_sbox_x5y6sw__prog_we_o)
        );
    tile_clb i_tile_x5y7 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x5y7__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x5y7__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x5y7sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x4y7ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x5y7sw__prog_we_o)
        ,.prog_din(_i_sbox_x5y7sw__prog_dout)
        ,.prog_dout(_i_tile_x5y7__prog_dout)
        ,.prog_we_o(_i_tile_x5y7__prog_we_o)
        );
    sbox_ne_S i_sbox_x5y7ne (
        .bi_x0y0e_L1(_i_sbox_x5y7nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x5y7ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x5y8ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x6y8se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x5y7__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x5y8se__prog_we_o)
        ,.prog_din(_i_sbox_x5y8se__prog_dout)
        ,.prog_dout(_i_sbox_x5y7ne__prog_dout)
        ,.prog_we_o(_i_sbox_x5y7ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x5y7nw (
        .bi_u1y0n_L1(_i_sbox_x5y7sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x5y7nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x4y7nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x4y8ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x5y7__prog_we_o)
        ,.prog_din(_i_tile_x5y7__prog_dout)
        ,.prog_dout(_i_sbox_x5y7nw__prog_dout)
        ,.prog_we_o(_i_sbox_x5y7nw__prog_we_o)
        );
    sbox_se_W i_sbox_x5y7se (
        .bi_x0v1n_L1(_i_sbox_x6y6sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x5y7se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x5y7ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x6y7se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x5y7ne__prog_we_o)
        ,.prog_din(_i_sbox_x5y7ne__prog_dout)
        ,.prog_dout(_i_sbox_x5y7se__prog_dout)
        ,.prog_we_o(_i_sbox_x5y7se__prog_we_o)
        );
    sbox_sw_N i_sbox_x5y7sw (
        .bi_u1v1n_L1(_i_sbox_x5y6sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x5y7sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x4y6nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x5y7se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x4y7__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x5y6nw__prog_we_o)
        ,.prog_din(_i_sbox_x5y6nw__prog_dout)
        ,.prog_dout(_i_sbox_x5y7sw__prog_dout)
        ,.prog_we_o(_i_sbox_x5y7sw__prog_we_o)
        );
    tile_clb i_tile_x5y8 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x5y8__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x5y8__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x5y8sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x4y8ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x5y8sw__prog_we_o)
        ,.prog_din(_i_sbox_x5y8sw__prog_dout)
        ,.prog_dout(_i_tile_x5y8__prog_dout)
        ,.prog_we_o(_i_tile_x5y8__prog_we_o)
        );
    sbox_ne_S_ex_s i_sbox_x5y8ne (
        .bi_x0y0e_L1(_i_sbox_x5y8nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x5y8ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x6y9se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x5y8__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x5y9se__prog_we_o)
        ,.prog_din(_i_sbox_x5y9se__prog_dout)
        ,.prog_dout(_i_sbox_x5y8ne__prog_dout)
        ,.prog_we_o(_i_sbox_x5y8ne__prog_we_o)
        );
    sbox_nw_E_ex_s i_sbox_x5y8nw (
        .bi_u1y0n_L1(_i_sbox_x5y8sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x5y8nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x4y8nw__so_x0y0e_L1)
        ,.cu_x0y0e_L1(_i_tile_x5y9__cu_x0v1e_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x5y8__prog_we_o)
        ,.prog_din(_i_tile_x5y8__prog_dout)
        ,.prog_dout(_i_sbox_x5y8nw__prog_dout)
        ,.prog_we_o(_i_sbox_x5y8nw__prog_we_o)
        );
    sbox_se_W i_sbox_x5y8se (
        .bi_x0v1n_L1(_i_sbox_x6y7sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x5y8se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x5y8ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x6y8se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x5y8ne__prog_we_o)
        ,.prog_din(_i_sbox_x5y8ne__prog_dout)
        ,.prog_dout(_i_sbox_x5y8se__prog_dout)
        ,.prog_we_o(_i_sbox_x5y8se__prog_we_o)
        );
    sbox_sw_N i_sbox_x5y8sw (
        .bi_u1v1n_L1(_i_sbox_x5y7sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x5y8sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x4y7nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x5y8se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x4y8__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x5y7nw__prog_we_o)
        ,.prog_din(_i_sbox_x5y7nw__prog_dout)
        ,.prog_dout(_i_sbox_x5y8sw__prog_dout)
        ,.prog_we_o(_i_sbox_x5y8sw__prog_we_o)
        );
    t_io_n i_tile_x5y9 (
        .bi_x0v1e_L1(_i_sbox_x5y8nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x5y9se__so_x0v1w_L1)
        ,.cu_x0v1e_L1(_i_tile_x5y9__cu_x0v1e_L1)
        ,.cu_x0v1w_L1(_i_tile_x5y9__cu_x0v1w_L1)
        ,.ipin_x0y0_0(ipin_x5y9_0)
        ,.opin_x0y0_0(_i_tile_x5y9__opin_x0y0_0)
        ,.oe_x0y0_0(_i_tile_x5y9__oe_x0y0_0)
        ,.ipin_x0y0_1(ipin_x5y9_1)
        ,.opin_x0y0_1(_i_tile_x5y9__opin_x0y0_1)
        ,.oe_x0y0_1(_i_tile_x5y9__oe_x0y0_1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x5y8nw__prog_we_o)
        ,.prog_din(_i_sbox_x5y8nw__prog_dout)
        ,.prog_dout(_i_tile_x5y9__prog_dout)
        ,.prog_we_o(_i_tile_x5y9__prog_we_o)
        );
    sbox_se_W_ex_s i_sbox_x5y9se (
        .bi_x0v1n_L1(_i_sbox_x6y8sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x5y9se__so_x0v1w_L1)
        ,.bi_x1v1w_L1(_i_sbox_x6y9se__so_x0v1w_L1)
        ,.cu_x0v1w_L1(_i_tile_x5y9__cu_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x5y9__prog_we_o)
        ,.prog_din(_i_tile_x5y9__prog_dout)
        ,.prog_dout(_i_sbox_x5y9se__prog_dout)
        ,.prog_we_o(_i_sbox_x5y9se__prog_we_o)
        );
    sbox_sw_s_ex_s i_sbox_x5y9sw (
        .bi_u1v1e_L1(_i_sbox_x4y8nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x5y9se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_ne_n_ex_n i_sbox_x6y0ne (
        .bi_x0y0e_L1(_i_sbox_x6y0nw__so_x0y0e_L1)
        ,.bi_x1y0w_L1(_i_sbox_x7y1se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_nw_E_ex_n i_sbox_x6y0nw (
        .bi_u1y0e_L1(_i_sbox_x5y0nw__so_x0y0e_L1)
        ,.so_x0y0e_L1(_i_sbox_x6y0nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x5y1ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x5y1se__prog_we_o)
        ,.prog_din(_i_sbox_x5y1se__prog_dout)
        ,.prog_dout(_i_sbox_x6y0nw__prog_dout)
        ,.prog_we_o(_i_sbox_x6y0nw__prog_we_o)
        );
    tile_clb i_tile_x6y1 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x6y1__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x6y1__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x6y1sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x5y1ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x6y1sw__prog_we_o)
        ,.prog_din(_i_sbox_x6y1sw__prog_dout)
        ,.prog_dout(_i_tile_x6y1__prog_dout)
        ,.prog_we_o(_i_tile_x6y1__prog_we_o)
        );
    sbox_ne_S i_sbox_x6y1ne (
        .bi_x0y0e_L1(_i_sbox_x6y1nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x6y1ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x6y2ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x7y2se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x6y1__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x6y2se__prog_we_o)
        ,.prog_din(_i_sbox_x6y2se__prog_dout)
        ,.prog_dout(_i_sbox_x6y1ne__prog_dout)
        ,.prog_we_o(_i_sbox_x6y1ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x6y1nw (
        .bi_u1y0n_L1(_i_sbox_x6y1sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x6y1nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x5y1nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x5y2ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x6y1__prog_we_o)
        ,.prog_din(_i_tile_x6y1__prog_dout)
        ,.prog_dout(_i_sbox_x6y1nw__prog_dout)
        ,.prog_we_o(_i_sbox_x6y1nw__prog_we_o)
        );
    sbox_se_W_ex_n i_sbox_x6y1se (
        .bi_x0y0s_L1(_i_sbox_x6y1ne__so_x0y0s_L1)
        ,.so_x0v1w_L1(_i_sbox_x6y1se__so_x0v1w_L1)
        ,.bi_x1v1w_L1(_i_sbox_x7y1se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x6y1ne__prog_we_o)
        ,.prog_din(_i_sbox_x6y1ne__prog_dout)
        ,.prog_dout(_i_sbox_x6y1se__prog_dout)
        ,.prog_we_o(_i_sbox_x6y1se__prog_we_o)
        );
    sbox_sw_N_ex_n i_sbox_x6y1sw (
        .bi_u1v1e_L1(_i_sbox_x5y0nw__so_x0y0e_L1)
        ,.so_u1y0n_L1(_i_sbox_x6y1sw__so_u1y0n_L1)
        ,.bi_x0v1w_L1(_i_sbox_x6y1se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x5y1__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x6y0nw__prog_we_o)
        ,.prog_din(_i_sbox_x6y0nw__prog_dout)
        ,.prog_dout(_i_sbox_x6y1sw__prog_dout)
        ,.prog_we_o(_i_sbox_x6y1sw__prog_we_o)
        );
    tile_clb i_tile_x6y2 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x6y2__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x6y2__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x6y2sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x5y2ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x6y2sw__prog_we_o)
        ,.prog_din(_i_sbox_x6y2sw__prog_dout)
        ,.prog_dout(_i_tile_x6y2__prog_dout)
        ,.prog_we_o(_i_tile_x6y2__prog_we_o)
        );
    sbox_ne_S i_sbox_x6y2ne (
        .bi_x0y0e_L1(_i_sbox_x6y2nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x6y2ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x6y3ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x7y3se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x6y2__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x6y3se__prog_we_o)
        ,.prog_din(_i_sbox_x6y3se__prog_dout)
        ,.prog_dout(_i_sbox_x6y2ne__prog_dout)
        ,.prog_we_o(_i_sbox_x6y2ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x6y2nw (
        .bi_u1y0n_L1(_i_sbox_x6y2sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x6y2nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x5y2nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x5y3ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x6y2__prog_we_o)
        ,.prog_din(_i_tile_x6y2__prog_dout)
        ,.prog_dout(_i_sbox_x6y2nw__prog_dout)
        ,.prog_we_o(_i_sbox_x6y2nw__prog_we_o)
        );
    sbox_se_W i_sbox_x6y2se (
        .bi_x0v1n_L1(_i_sbox_x7y1sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x6y2se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x6y2ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x7y2se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x6y2ne__prog_we_o)
        ,.prog_din(_i_sbox_x6y2ne__prog_dout)
        ,.prog_dout(_i_sbox_x6y2se__prog_dout)
        ,.prog_we_o(_i_sbox_x6y2se__prog_we_o)
        );
    sbox_sw_N i_sbox_x6y2sw (
        .bi_u1v1n_L1(_i_sbox_x6y1sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x6y2sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x5y1nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x6y2se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x5y2__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x6y1nw__prog_we_o)
        ,.prog_din(_i_sbox_x6y1nw__prog_dout)
        ,.prog_dout(_i_sbox_x6y2sw__prog_dout)
        ,.prog_we_o(_i_sbox_x6y2sw__prog_we_o)
        );
    tile_clb i_tile_x6y3 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x6y3__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x6y3__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x6y3sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x5y3ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x6y3sw__prog_we_o)
        ,.prog_din(_i_sbox_x6y3sw__prog_dout)
        ,.prog_dout(_i_tile_x6y3__prog_dout)
        ,.prog_we_o(_i_tile_x6y3__prog_we_o)
        );
    sbox_ne_S i_sbox_x6y3ne (
        .bi_x0y0e_L1(_i_sbox_x6y3nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x6y3ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x6y4ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x7y4se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x6y3__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x6y4se__prog_we_o)
        ,.prog_din(_i_sbox_x6y4se__prog_dout)
        ,.prog_dout(_i_sbox_x6y3ne__prog_dout)
        ,.prog_we_o(_i_sbox_x6y3ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x6y3nw (
        .bi_u1y0n_L1(_i_sbox_x6y3sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x6y3nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x5y3nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x5y4ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x6y3__prog_we_o)
        ,.prog_din(_i_tile_x6y3__prog_dout)
        ,.prog_dout(_i_sbox_x6y3nw__prog_dout)
        ,.prog_we_o(_i_sbox_x6y3nw__prog_we_o)
        );
    sbox_se_W i_sbox_x6y3se (
        .bi_x0v1n_L1(_i_sbox_x7y2sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x6y3se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x6y3ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x7y3se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x6y3ne__prog_we_o)
        ,.prog_din(_i_sbox_x6y3ne__prog_dout)
        ,.prog_dout(_i_sbox_x6y3se__prog_dout)
        ,.prog_we_o(_i_sbox_x6y3se__prog_we_o)
        );
    sbox_sw_N i_sbox_x6y3sw (
        .bi_u1v1n_L1(_i_sbox_x6y2sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x6y3sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x5y2nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x6y3se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x5y3__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x6y2nw__prog_we_o)
        ,.prog_din(_i_sbox_x6y2nw__prog_dout)
        ,.prog_dout(_i_sbox_x6y3sw__prog_dout)
        ,.prog_we_o(_i_sbox_x6y3sw__prog_we_o)
        );
    tile_clb i_tile_x6y4 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x6y4__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x6y4__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x6y4sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x5y4ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x6y4sw__prog_we_o)
        ,.prog_din(_i_sbox_x6y4sw__prog_dout)
        ,.prog_dout(_i_tile_x6y4__prog_dout)
        ,.prog_we_o(_i_tile_x6y4__prog_we_o)
        );
    sbox_ne_S i_sbox_x6y4ne (
        .bi_x0y0e_L1(_i_sbox_x6y4nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x6y4ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x6y5ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x7y5se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x6y4__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x6y5se__prog_we_o)
        ,.prog_din(_i_sbox_x6y5se__prog_dout)
        ,.prog_dout(_i_sbox_x6y4ne__prog_dout)
        ,.prog_we_o(_i_sbox_x6y4ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x6y4nw (
        .bi_u1y0n_L1(_i_sbox_x6y4sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x6y4nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x5y4nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x5y5ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x6y4__prog_we_o)
        ,.prog_din(_i_tile_x6y4__prog_dout)
        ,.prog_dout(_i_sbox_x6y4nw__prog_dout)
        ,.prog_we_o(_i_sbox_x6y4nw__prog_we_o)
        );
    sbox_se_W i_sbox_x6y4se (
        .bi_x0v1n_L1(_i_sbox_x7y3sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x6y4se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x6y4ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x7y4se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x6y4ne__prog_we_o)
        ,.prog_din(_i_sbox_x6y4ne__prog_dout)
        ,.prog_dout(_i_sbox_x6y4se__prog_dout)
        ,.prog_we_o(_i_sbox_x6y4se__prog_we_o)
        );
    sbox_sw_N i_sbox_x6y4sw (
        .bi_u1v1n_L1(_i_sbox_x6y3sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x6y4sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x5y3nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x6y4se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x5y4__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x6y3nw__prog_we_o)
        ,.prog_din(_i_sbox_x6y3nw__prog_dout)
        ,.prog_dout(_i_sbox_x6y4sw__prog_dout)
        ,.prog_we_o(_i_sbox_x6y4sw__prog_we_o)
        );
    tile_clb i_tile_x6y5 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x6y5__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x6y5__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x6y5sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x5y5ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x6y5sw__prog_we_o)
        ,.prog_din(_i_sbox_x6y5sw__prog_dout)
        ,.prog_dout(_i_tile_x6y5__prog_dout)
        ,.prog_we_o(_i_tile_x6y5__prog_we_o)
        );
    sbox_ne_S i_sbox_x6y5ne (
        .bi_x0y0e_L1(_i_sbox_x6y5nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x6y5ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x6y6ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x7y6se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x6y5__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x6y6se__prog_we_o)
        ,.prog_din(_i_sbox_x6y6se__prog_dout)
        ,.prog_dout(_i_sbox_x6y5ne__prog_dout)
        ,.prog_we_o(_i_sbox_x6y5ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x6y5nw (
        .bi_u1y0n_L1(_i_sbox_x6y5sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x6y5nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x5y5nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x5y6ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x6y5__prog_we_o)
        ,.prog_din(_i_tile_x6y5__prog_dout)
        ,.prog_dout(_i_sbox_x6y5nw__prog_dout)
        ,.prog_we_o(_i_sbox_x6y5nw__prog_we_o)
        );
    sbox_se_W i_sbox_x6y5se (
        .bi_x0v1n_L1(_i_sbox_x7y4sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x6y5se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x6y5ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x7y5se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x6y5ne__prog_we_o)
        ,.prog_din(_i_sbox_x6y5ne__prog_dout)
        ,.prog_dout(_i_sbox_x6y5se__prog_dout)
        ,.prog_we_o(_i_sbox_x6y5se__prog_we_o)
        );
    sbox_sw_N i_sbox_x6y5sw (
        .bi_u1v1n_L1(_i_sbox_x6y4sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x6y5sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x5y4nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x6y5se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x5y5__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x6y4nw__prog_we_o)
        ,.prog_din(_i_sbox_x6y4nw__prog_dout)
        ,.prog_dout(_i_sbox_x6y5sw__prog_dout)
        ,.prog_we_o(_i_sbox_x6y5sw__prog_we_o)
        );
    tile_clb i_tile_x6y6 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x6y6__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x6y6__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x6y6sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x5y6ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x6y6sw__prog_we_o)
        ,.prog_din(_i_sbox_x6y6sw__prog_dout)
        ,.prog_dout(_i_tile_x6y6__prog_dout)
        ,.prog_we_o(_i_tile_x6y6__prog_we_o)
        );
    sbox_ne_S i_sbox_x6y6ne (
        .bi_x0y0e_L1(_i_sbox_x6y6nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x6y6ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x6y7ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x7y7se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x6y6__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x6y7se__prog_we_o)
        ,.prog_din(_i_sbox_x6y7se__prog_dout)
        ,.prog_dout(_i_sbox_x6y6ne__prog_dout)
        ,.prog_we_o(_i_sbox_x6y6ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x6y6nw (
        .bi_u1y0n_L1(_i_sbox_x6y6sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x6y6nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x5y6nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x5y7ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x6y6__prog_we_o)
        ,.prog_din(_i_tile_x6y6__prog_dout)
        ,.prog_dout(_i_sbox_x6y6nw__prog_dout)
        ,.prog_we_o(_i_sbox_x6y6nw__prog_we_o)
        );
    sbox_se_W i_sbox_x6y6se (
        .bi_x0v1n_L1(_i_sbox_x7y5sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x6y6se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x6y6ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x7y6se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x6y6ne__prog_we_o)
        ,.prog_din(_i_sbox_x6y6ne__prog_dout)
        ,.prog_dout(_i_sbox_x6y6se__prog_dout)
        ,.prog_we_o(_i_sbox_x6y6se__prog_we_o)
        );
    sbox_sw_N i_sbox_x6y6sw (
        .bi_u1v1n_L1(_i_sbox_x6y5sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x6y6sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x5y5nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x6y6se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x5y6__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x6y5nw__prog_we_o)
        ,.prog_din(_i_sbox_x6y5nw__prog_dout)
        ,.prog_dout(_i_sbox_x6y6sw__prog_dout)
        ,.prog_we_o(_i_sbox_x6y6sw__prog_we_o)
        );
    tile_clb i_tile_x6y7 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x6y7__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x6y7__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x6y7sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x5y7ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x6y7sw__prog_we_o)
        ,.prog_din(_i_sbox_x6y7sw__prog_dout)
        ,.prog_dout(_i_tile_x6y7__prog_dout)
        ,.prog_we_o(_i_tile_x6y7__prog_we_o)
        );
    sbox_ne_S i_sbox_x6y7ne (
        .bi_x0y0e_L1(_i_sbox_x6y7nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x6y7ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x6y8ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x7y8se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x6y7__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x6y8se__prog_we_o)
        ,.prog_din(_i_sbox_x6y8se__prog_dout)
        ,.prog_dout(_i_sbox_x6y7ne__prog_dout)
        ,.prog_we_o(_i_sbox_x6y7ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x6y7nw (
        .bi_u1y0n_L1(_i_sbox_x6y7sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x6y7nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x5y7nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x5y8ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x6y7__prog_we_o)
        ,.prog_din(_i_tile_x6y7__prog_dout)
        ,.prog_dout(_i_sbox_x6y7nw__prog_dout)
        ,.prog_we_o(_i_sbox_x6y7nw__prog_we_o)
        );
    sbox_se_W i_sbox_x6y7se (
        .bi_x0v1n_L1(_i_sbox_x7y6sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x6y7se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x6y7ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x7y7se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x6y7ne__prog_we_o)
        ,.prog_din(_i_sbox_x6y7ne__prog_dout)
        ,.prog_dout(_i_sbox_x6y7se__prog_dout)
        ,.prog_we_o(_i_sbox_x6y7se__prog_we_o)
        );
    sbox_sw_N i_sbox_x6y7sw (
        .bi_u1v1n_L1(_i_sbox_x6y6sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x6y7sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x5y6nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x6y7se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x5y7__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x6y6nw__prog_we_o)
        ,.prog_din(_i_sbox_x6y6nw__prog_dout)
        ,.prog_dout(_i_sbox_x6y7sw__prog_dout)
        ,.prog_we_o(_i_sbox_x6y7sw__prog_we_o)
        );
    tile_clb i_tile_x6y8 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x6y8__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x6y8__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x6y8sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x5y8ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x6y8sw__prog_we_o)
        ,.prog_din(_i_sbox_x6y8sw__prog_dout)
        ,.prog_dout(_i_tile_x6y8__prog_dout)
        ,.prog_we_o(_i_tile_x6y8__prog_we_o)
        );
    sbox_ne_S_ex_s i_sbox_x6y8ne (
        .bi_x0y0e_L1(_i_sbox_x6y8nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x6y8ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x7y9se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x6y8__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x6y9se__prog_we_o)
        ,.prog_din(_i_sbox_x6y9se__prog_dout)
        ,.prog_dout(_i_sbox_x6y8ne__prog_dout)
        ,.prog_we_o(_i_sbox_x6y8ne__prog_we_o)
        );
    sbox_nw_E_ex_s i_sbox_x6y8nw (
        .bi_u1y0n_L1(_i_sbox_x6y8sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x6y8nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x5y8nw__so_x0y0e_L1)
        ,.cu_x0y0e_L1(_i_tile_x6y9__cu_x0v1e_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x6y8__prog_we_o)
        ,.prog_din(_i_tile_x6y8__prog_dout)
        ,.prog_dout(_i_sbox_x6y8nw__prog_dout)
        ,.prog_we_o(_i_sbox_x6y8nw__prog_we_o)
        );
    sbox_se_W i_sbox_x6y8se (
        .bi_x0v1n_L1(_i_sbox_x7y7sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x6y8se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x6y8ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x7y8se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x6y8ne__prog_we_o)
        ,.prog_din(_i_sbox_x6y8ne__prog_dout)
        ,.prog_dout(_i_sbox_x6y8se__prog_dout)
        ,.prog_we_o(_i_sbox_x6y8se__prog_we_o)
        );
    sbox_sw_N i_sbox_x6y8sw (
        .bi_u1v1n_L1(_i_sbox_x6y7sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x6y8sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x5y7nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x6y8se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x5y8__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x6y7nw__prog_we_o)
        ,.prog_din(_i_sbox_x6y7nw__prog_dout)
        ,.prog_dout(_i_sbox_x6y8sw__prog_dout)
        ,.prog_we_o(_i_sbox_x6y8sw__prog_we_o)
        );
    t_io_n i_tile_x6y9 (
        .bi_x0v1e_L1(_i_sbox_x6y8nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x6y9se__so_x0v1w_L1)
        ,.cu_x0v1e_L1(_i_tile_x6y9__cu_x0v1e_L1)
        ,.cu_x0v1w_L1(_i_tile_x6y9__cu_x0v1w_L1)
        ,.ipin_x0y0_0(ipin_x6y9_0)
        ,.opin_x0y0_0(_i_tile_x6y9__opin_x0y0_0)
        ,.oe_x0y0_0(_i_tile_x6y9__oe_x0y0_0)
        ,.ipin_x0y0_1(ipin_x6y9_1)
        ,.opin_x0y0_1(_i_tile_x6y9__opin_x0y0_1)
        ,.oe_x0y0_1(_i_tile_x6y9__oe_x0y0_1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x6y8nw__prog_we_o)
        ,.prog_din(_i_sbox_x6y8nw__prog_dout)
        ,.prog_dout(_i_tile_x6y9__prog_dout)
        ,.prog_we_o(_i_tile_x6y9__prog_we_o)
        );
    sbox_se_W_ex_s i_sbox_x6y9se (
        .bi_x0v1n_L1(_i_sbox_x7y8sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x6y9se__so_x0v1w_L1)
        ,.bi_x1v1w_L1(_i_sbox_x7y9se__so_x0v1w_L1)
        ,.cu_x0v1w_L1(_i_tile_x6y9__cu_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x6y9__prog_we_o)
        ,.prog_din(_i_tile_x6y9__prog_dout)
        ,.prog_dout(_i_sbox_x6y9se__prog_dout)
        ,.prog_we_o(_i_sbox_x6y9se__prog_we_o)
        );
    sbox_sw_s_ex_s i_sbox_x6y9sw (
        .bi_u1v1e_L1(_i_sbox_x5y8nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x6y9se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_ne_n_ex_n i_sbox_x7y0ne (
        .bi_x0y0e_L1(_i_sbox_x7y0nw__so_x0y0e_L1)
        ,.bi_x1y0w_L1(_i_sbox_x8y1se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_nw_E_ex_n i_sbox_x7y0nw (
        .bi_u1y0e_L1(_i_sbox_x6y0nw__so_x0y0e_L1)
        ,.so_x0y0e_L1(_i_sbox_x7y0nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x6y1ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x6y1se__prog_we_o)
        ,.prog_din(_i_sbox_x6y1se__prog_dout)
        ,.prog_dout(_i_sbox_x7y0nw__prog_dout)
        ,.prog_we_o(_i_sbox_x7y0nw__prog_we_o)
        );
    tile_clb i_tile_x7y1 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x7y1__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x7y1__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x7y1sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x6y1ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x7y1sw__prog_we_o)
        ,.prog_din(_i_sbox_x7y1sw__prog_dout)
        ,.prog_dout(_i_tile_x7y1__prog_dout)
        ,.prog_we_o(_i_tile_x7y1__prog_we_o)
        );
    sbox_ne_S i_sbox_x7y1ne (
        .bi_x0y0e_L1(_i_sbox_x7y1nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x7y1ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x7y2ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x8y2se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x7y1__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x7y2se__prog_we_o)
        ,.prog_din(_i_sbox_x7y2se__prog_dout)
        ,.prog_dout(_i_sbox_x7y1ne__prog_dout)
        ,.prog_we_o(_i_sbox_x7y1ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x7y1nw (
        .bi_u1y0n_L1(_i_sbox_x7y1sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x7y1nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x6y1nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x6y2ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x7y1__prog_we_o)
        ,.prog_din(_i_tile_x7y1__prog_dout)
        ,.prog_dout(_i_sbox_x7y1nw__prog_dout)
        ,.prog_we_o(_i_sbox_x7y1nw__prog_we_o)
        );
    sbox_se_W_ex_n i_sbox_x7y1se (
        .bi_x0y0s_L1(_i_sbox_x7y1ne__so_x0y0s_L1)
        ,.so_x0v1w_L1(_i_sbox_x7y1se__so_x0v1w_L1)
        ,.bi_x1v1w_L1(_i_sbox_x8y1se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x7y1ne__prog_we_o)
        ,.prog_din(_i_sbox_x7y1ne__prog_dout)
        ,.prog_dout(_i_sbox_x7y1se__prog_dout)
        ,.prog_we_o(_i_sbox_x7y1se__prog_we_o)
        );
    sbox_sw_N_ex_n i_sbox_x7y1sw (
        .bi_u1v1e_L1(_i_sbox_x6y0nw__so_x0y0e_L1)
        ,.so_u1y0n_L1(_i_sbox_x7y1sw__so_u1y0n_L1)
        ,.bi_x0v1w_L1(_i_sbox_x7y1se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x6y1__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x7y0nw__prog_we_o)
        ,.prog_din(_i_sbox_x7y0nw__prog_dout)
        ,.prog_dout(_i_sbox_x7y1sw__prog_dout)
        ,.prog_we_o(_i_sbox_x7y1sw__prog_we_o)
        );
    tile_clb i_tile_x7y2 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x7y2__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x7y2__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x7y2sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x6y2ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x7y2sw__prog_we_o)
        ,.prog_din(_i_sbox_x7y2sw__prog_dout)
        ,.prog_dout(_i_tile_x7y2__prog_dout)
        ,.prog_we_o(_i_tile_x7y2__prog_we_o)
        );
    sbox_ne_S i_sbox_x7y2ne (
        .bi_x0y0e_L1(_i_sbox_x7y2nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x7y2ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x7y3ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x8y3se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x7y2__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x7y3se__prog_we_o)
        ,.prog_din(_i_sbox_x7y3se__prog_dout)
        ,.prog_dout(_i_sbox_x7y2ne__prog_dout)
        ,.prog_we_o(_i_sbox_x7y2ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x7y2nw (
        .bi_u1y0n_L1(_i_sbox_x7y2sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x7y2nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x6y2nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x6y3ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x7y2__prog_we_o)
        ,.prog_din(_i_tile_x7y2__prog_dout)
        ,.prog_dout(_i_sbox_x7y2nw__prog_dout)
        ,.prog_we_o(_i_sbox_x7y2nw__prog_we_o)
        );
    sbox_se_W i_sbox_x7y2se (
        .bi_x0v1n_L1(_i_sbox_x8y1sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x7y2se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x7y2ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x8y2se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x7y2ne__prog_we_o)
        ,.prog_din(_i_sbox_x7y2ne__prog_dout)
        ,.prog_dout(_i_sbox_x7y2se__prog_dout)
        ,.prog_we_o(_i_sbox_x7y2se__prog_we_o)
        );
    sbox_sw_N i_sbox_x7y2sw (
        .bi_u1v1n_L1(_i_sbox_x7y1sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x7y2sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x6y1nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x7y2se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x6y2__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x7y1nw__prog_we_o)
        ,.prog_din(_i_sbox_x7y1nw__prog_dout)
        ,.prog_dout(_i_sbox_x7y2sw__prog_dout)
        ,.prog_we_o(_i_sbox_x7y2sw__prog_we_o)
        );
    tile_clb i_tile_x7y3 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x7y3__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x7y3__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x7y3sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x6y3ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x7y3sw__prog_we_o)
        ,.prog_din(_i_sbox_x7y3sw__prog_dout)
        ,.prog_dout(_i_tile_x7y3__prog_dout)
        ,.prog_we_o(_i_tile_x7y3__prog_we_o)
        );
    sbox_ne_S i_sbox_x7y3ne (
        .bi_x0y0e_L1(_i_sbox_x7y3nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x7y3ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x7y4ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x8y4se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x7y3__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x7y4se__prog_we_o)
        ,.prog_din(_i_sbox_x7y4se__prog_dout)
        ,.prog_dout(_i_sbox_x7y3ne__prog_dout)
        ,.prog_we_o(_i_sbox_x7y3ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x7y3nw (
        .bi_u1y0n_L1(_i_sbox_x7y3sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x7y3nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x6y3nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x6y4ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x7y3__prog_we_o)
        ,.prog_din(_i_tile_x7y3__prog_dout)
        ,.prog_dout(_i_sbox_x7y3nw__prog_dout)
        ,.prog_we_o(_i_sbox_x7y3nw__prog_we_o)
        );
    sbox_se_W i_sbox_x7y3se (
        .bi_x0v1n_L1(_i_sbox_x8y2sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x7y3se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x7y3ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x8y3se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x7y3ne__prog_we_o)
        ,.prog_din(_i_sbox_x7y3ne__prog_dout)
        ,.prog_dout(_i_sbox_x7y3se__prog_dout)
        ,.prog_we_o(_i_sbox_x7y3se__prog_we_o)
        );
    sbox_sw_N i_sbox_x7y3sw (
        .bi_u1v1n_L1(_i_sbox_x7y2sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x7y3sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x6y2nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x7y3se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x6y3__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x7y2nw__prog_we_o)
        ,.prog_din(_i_sbox_x7y2nw__prog_dout)
        ,.prog_dout(_i_sbox_x7y3sw__prog_dout)
        ,.prog_we_o(_i_sbox_x7y3sw__prog_we_o)
        );
    tile_clb i_tile_x7y4 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x7y4__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x7y4__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x7y4sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x6y4ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x7y4sw__prog_we_o)
        ,.prog_din(_i_sbox_x7y4sw__prog_dout)
        ,.prog_dout(_i_tile_x7y4__prog_dout)
        ,.prog_we_o(_i_tile_x7y4__prog_we_o)
        );
    sbox_ne_S i_sbox_x7y4ne (
        .bi_x0y0e_L1(_i_sbox_x7y4nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x7y4ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x7y5ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x8y5se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x7y4__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x7y5se__prog_we_o)
        ,.prog_din(_i_sbox_x7y5se__prog_dout)
        ,.prog_dout(_i_sbox_x7y4ne__prog_dout)
        ,.prog_we_o(_i_sbox_x7y4ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x7y4nw (
        .bi_u1y0n_L1(_i_sbox_x7y4sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x7y4nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x6y4nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x6y5ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x7y4__prog_we_o)
        ,.prog_din(_i_tile_x7y4__prog_dout)
        ,.prog_dout(_i_sbox_x7y4nw__prog_dout)
        ,.prog_we_o(_i_sbox_x7y4nw__prog_we_o)
        );
    sbox_se_W i_sbox_x7y4se (
        .bi_x0v1n_L1(_i_sbox_x8y3sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x7y4se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x7y4ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x8y4se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x7y4ne__prog_we_o)
        ,.prog_din(_i_sbox_x7y4ne__prog_dout)
        ,.prog_dout(_i_sbox_x7y4se__prog_dout)
        ,.prog_we_o(_i_sbox_x7y4se__prog_we_o)
        );
    sbox_sw_N i_sbox_x7y4sw (
        .bi_u1v1n_L1(_i_sbox_x7y3sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x7y4sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x6y3nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x7y4se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x6y4__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x7y3nw__prog_we_o)
        ,.prog_din(_i_sbox_x7y3nw__prog_dout)
        ,.prog_dout(_i_sbox_x7y4sw__prog_dout)
        ,.prog_we_o(_i_sbox_x7y4sw__prog_we_o)
        );
    tile_clb i_tile_x7y5 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x7y5__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x7y5__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x7y5sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x6y5ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x7y5sw__prog_we_o)
        ,.prog_din(_i_sbox_x7y5sw__prog_dout)
        ,.prog_dout(_i_tile_x7y5__prog_dout)
        ,.prog_we_o(_i_tile_x7y5__prog_we_o)
        );
    sbox_ne_S i_sbox_x7y5ne (
        .bi_x0y0e_L1(_i_sbox_x7y5nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x7y5ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x7y6ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x8y6se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x7y5__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x7y6se__prog_we_o)
        ,.prog_din(_i_sbox_x7y6se__prog_dout)
        ,.prog_dout(_i_sbox_x7y5ne__prog_dout)
        ,.prog_we_o(_i_sbox_x7y5ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x7y5nw (
        .bi_u1y0n_L1(_i_sbox_x7y5sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x7y5nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x6y5nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x6y6ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x7y5__prog_we_o)
        ,.prog_din(_i_tile_x7y5__prog_dout)
        ,.prog_dout(_i_sbox_x7y5nw__prog_dout)
        ,.prog_we_o(_i_sbox_x7y5nw__prog_we_o)
        );
    sbox_se_W i_sbox_x7y5se (
        .bi_x0v1n_L1(_i_sbox_x8y4sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x7y5se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x7y5ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x8y5se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x7y5ne__prog_we_o)
        ,.prog_din(_i_sbox_x7y5ne__prog_dout)
        ,.prog_dout(_i_sbox_x7y5se__prog_dout)
        ,.prog_we_o(_i_sbox_x7y5se__prog_we_o)
        );
    sbox_sw_N i_sbox_x7y5sw (
        .bi_u1v1n_L1(_i_sbox_x7y4sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x7y5sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x6y4nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x7y5se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x6y5__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x7y4nw__prog_we_o)
        ,.prog_din(_i_sbox_x7y4nw__prog_dout)
        ,.prog_dout(_i_sbox_x7y5sw__prog_dout)
        ,.prog_we_o(_i_sbox_x7y5sw__prog_we_o)
        );
    tile_clb i_tile_x7y6 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x7y6__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x7y6__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x7y6sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x6y6ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x7y6sw__prog_we_o)
        ,.prog_din(_i_sbox_x7y6sw__prog_dout)
        ,.prog_dout(_i_tile_x7y6__prog_dout)
        ,.prog_we_o(_i_tile_x7y6__prog_we_o)
        );
    sbox_ne_S i_sbox_x7y6ne (
        .bi_x0y0e_L1(_i_sbox_x7y6nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x7y6ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x7y7ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x8y7se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x7y6__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x7y7se__prog_we_o)
        ,.prog_din(_i_sbox_x7y7se__prog_dout)
        ,.prog_dout(_i_sbox_x7y6ne__prog_dout)
        ,.prog_we_o(_i_sbox_x7y6ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x7y6nw (
        .bi_u1y0n_L1(_i_sbox_x7y6sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x7y6nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x6y6nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x6y7ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x7y6__prog_we_o)
        ,.prog_din(_i_tile_x7y6__prog_dout)
        ,.prog_dout(_i_sbox_x7y6nw__prog_dout)
        ,.prog_we_o(_i_sbox_x7y6nw__prog_we_o)
        );
    sbox_se_W i_sbox_x7y6se (
        .bi_x0v1n_L1(_i_sbox_x8y5sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x7y6se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x7y6ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x8y6se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x7y6ne__prog_we_o)
        ,.prog_din(_i_sbox_x7y6ne__prog_dout)
        ,.prog_dout(_i_sbox_x7y6se__prog_dout)
        ,.prog_we_o(_i_sbox_x7y6se__prog_we_o)
        );
    sbox_sw_N i_sbox_x7y6sw (
        .bi_u1v1n_L1(_i_sbox_x7y5sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x7y6sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x6y5nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x7y6se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x6y6__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x7y5nw__prog_we_o)
        ,.prog_din(_i_sbox_x7y5nw__prog_dout)
        ,.prog_dout(_i_sbox_x7y6sw__prog_dout)
        ,.prog_we_o(_i_sbox_x7y6sw__prog_we_o)
        );
    tile_clb i_tile_x7y7 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x7y7__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x7y7__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x7y7sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x6y7ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x7y7sw__prog_we_o)
        ,.prog_din(_i_sbox_x7y7sw__prog_dout)
        ,.prog_dout(_i_tile_x7y7__prog_dout)
        ,.prog_we_o(_i_tile_x7y7__prog_we_o)
        );
    sbox_ne_S i_sbox_x7y7ne (
        .bi_x0y0e_L1(_i_sbox_x7y7nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x7y7ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x7y8ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x8y8se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x7y7__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x7y8se__prog_we_o)
        ,.prog_din(_i_sbox_x7y8se__prog_dout)
        ,.prog_dout(_i_sbox_x7y7ne__prog_dout)
        ,.prog_we_o(_i_sbox_x7y7ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x7y7nw (
        .bi_u1y0n_L1(_i_sbox_x7y7sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x7y7nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x6y7nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x6y8ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x7y7__prog_we_o)
        ,.prog_din(_i_tile_x7y7__prog_dout)
        ,.prog_dout(_i_sbox_x7y7nw__prog_dout)
        ,.prog_we_o(_i_sbox_x7y7nw__prog_we_o)
        );
    sbox_se_W i_sbox_x7y7se (
        .bi_x0v1n_L1(_i_sbox_x8y6sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x7y7se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x7y7ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x8y7se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x7y7ne__prog_we_o)
        ,.prog_din(_i_sbox_x7y7ne__prog_dout)
        ,.prog_dout(_i_sbox_x7y7se__prog_dout)
        ,.prog_we_o(_i_sbox_x7y7se__prog_we_o)
        );
    sbox_sw_N i_sbox_x7y7sw (
        .bi_u1v1n_L1(_i_sbox_x7y6sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x7y7sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x6y6nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x7y7se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x6y7__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x7y6nw__prog_we_o)
        ,.prog_din(_i_sbox_x7y6nw__prog_dout)
        ,.prog_dout(_i_sbox_x7y7sw__prog_dout)
        ,.prog_we_o(_i_sbox_x7y7sw__prog_we_o)
        );
    tile_clb i_tile_x7y8 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x7y8__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x7y8__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x7y8sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x6y8ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x7y8sw__prog_we_o)
        ,.prog_din(_i_sbox_x7y8sw__prog_dout)
        ,.prog_dout(_i_tile_x7y8__prog_dout)
        ,.prog_we_o(_i_tile_x7y8__prog_we_o)
        );
    sbox_ne_S_ex_s i_sbox_x7y8ne (
        .bi_x0y0e_L1(_i_sbox_x7y8nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x7y8ne__so_x0y0s_L1)
        ,.bi_x1y0w_L1(_i_sbox_x8y9se__so_x0v1w_L1)
        ,.cu_x0y0s_L1(_i_tile_x7y8__cu_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x7y9se__prog_we_o)
        ,.prog_din(_i_sbox_x7y9se__prog_dout)
        ,.prog_dout(_i_sbox_x7y8ne__prog_dout)
        ,.prog_we_o(_i_sbox_x7y8ne__prog_we_o)
        );
    sbox_nw_E_ex_s i_sbox_x7y8nw (
        .bi_u1y0n_L1(_i_sbox_x7y8sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x7y8nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x6y8nw__so_x0y0e_L1)
        ,.cu_x0y0e_L1(_i_tile_x7y9__cu_x0v1e_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x7y8__prog_we_o)
        ,.prog_din(_i_tile_x7y8__prog_dout)
        ,.prog_dout(_i_sbox_x7y8nw__prog_dout)
        ,.prog_we_o(_i_sbox_x7y8nw__prog_we_o)
        );
    sbox_se_W i_sbox_x7y8se (
        .bi_x0v1n_L1(_i_sbox_x8y7sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x7y8se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x7y8ne__so_x0y0s_L1)
        ,.bi_x1v1w_L1(_i_sbox_x8y8se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x7y8ne__prog_we_o)
        ,.prog_din(_i_sbox_x7y8ne__prog_dout)
        ,.prog_dout(_i_sbox_x7y8se__prog_dout)
        ,.prog_we_o(_i_sbox_x7y8se__prog_we_o)
        );
    sbox_sw_N i_sbox_x7y8sw (
        .bi_u1v1n_L1(_i_sbox_x7y7sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x7y8sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x6y7nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x7y8se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x6y8__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x7y7nw__prog_we_o)
        ,.prog_din(_i_sbox_x7y7nw__prog_dout)
        ,.prog_dout(_i_sbox_x7y8sw__prog_dout)
        ,.prog_we_o(_i_sbox_x7y8sw__prog_we_o)
        );
    t_io_n i_tile_x7y9 (
        .bi_x0v1e_L1(_i_sbox_x7y8nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x7y9se__so_x0v1w_L1)
        ,.cu_x0v1e_L1(_i_tile_x7y9__cu_x0v1e_L1)
        ,.cu_x0v1w_L1(_i_tile_x7y9__cu_x0v1w_L1)
        ,.ipin_x0y0_0(ipin_x7y9_0)
        ,.opin_x0y0_0(_i_tile_x7y9__opin_x0y0_0)
        ,.oe_x0y0_0(_i_tile_x7y9__oe_x0y0_0)
        ,.ipin_x0y0_1(ipin_x7y9_1)
        ,.opin_x0y0_1(_i_tile_x7y9__opin_x0y0_1)
        ,.oe_x0y0_1(_i_tile_x7y9__oe_x0y0_1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x7y8nw__prog_we_o)
        ,.prog_din(_i_sbox_x7y8nw__prog_dout)
        ,.prog_dout(_i_tile_x7y9__prog_dout)
        ,.prog_we_o(_i_tile_x7y9__prog_we_o)
        );
    sbox_se_W_ex_s i_sbox_x7y9se (
        .bi_x0v1n_L1(_i_sbox_x8y8sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x7y9se__so_x0v1w_L1)
        ,.bi_x1v1w_L1(_i_sbox_x8y9se__so_x0v1w_L1)
        ,.cu_x0v1w_L1(_i_tile_x7y9__cu_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x7y9__prog_we_o)
        ,.prog_din(_i_tile_x7y9__prog_dout)
        ,.prog_dout(_i_sbox_x7y9se__prog_dout)
        ,.prog_we_o(_i_sbox_x7y9se__prog_we_o)
        );
    sbox_sw_s_ex_s i_sbox_x7y9sw (
        .bi_u1v1e_L1(_i_sbox_x6y8nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x7y9se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_ne_n_ex_nw i_sbox_x8y0ne (
        .bi_x0y0e_L1(_i_sbox_x8y0nw__so_x0y0e_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_nw_E_ex_n i_sbox_x8y0nw (
        .bi_u1y0e_L1(_i_sbox_x7y0nw__so_x0y0e_L1)
        ,.so_x0y0e_L1(_i_sbox_x8y0nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x7y1ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x7y1se__prog_we_o)
        ,.prog_din(_i_sbox_x7y1se__prog_dout)
        ,.prog_dout(_i_sbox_x8y0nw__prog_dout)
        ,.prog_we_o(_i_sbox_x8y0nw__prog_we_o)
        );
    tile_clb i_tile_x8y1 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x8y1__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x8y1__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x8y1sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x7y1ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x8y1sw__prog_we_o)
        ,.prog_din(_i_sbox_x8y1sw__prog_dout)
        ,.prog_dout(_i_tile_x8y1__prog_dout)
        ,.prog_we_o(_i_tile_x8y1__prog_we_o)
        );
    sbox_ne_S_ex_w i_sbox_x8y1ne (
        .bi_x0y0e_L1(_i_sbox_x8y1nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x8y1ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x8y2ne__so_x0y0s_L1)
        ,.cu_x0y0s_L1(_i_tile_x8y1__cu_x0y0s_L1)
        ,.cv_x0y0s_L1(_i_tile_x9y1__cu_u1y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x8y2se__prog_we_o)
        ,.prog_din(_i_sbox_x8y2se__prog_dout)
        ,.prog_dout(_i_sbox_x8y1ne__prog_dout)
        ,.prog_we_o(_i_sbox_x8y1ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x8y1nw (
        .bi_u1y0n_L1(_i_sbox_x8y1sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x8y1nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x7y1nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x7y2ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x8y1__prog_we_o)
        ,.prog_din(_i_tile_x8y1__prog_dout)
        ,.prog_dout(_i_sbox_x8y1nw__prog_dout)
        ,.prog_we_o(_i_sbox_x8y1nw__prog_we_o)
        );
    sbox_se_W_ex_nw i_sbox_x8y1se (
        .bi_x0y0s_L1(_i_sbox_x8y1ne__so_x0y0s_L1)
        ,.so_x0v1w_L1(_i_sbox_x8y1se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x8y1ne__prog_we_o)
        ,.prog_din(_i_sbox_x8y1ne__prog_dout)
        ,.prog_dout(_i_sbox_x8y1se__prog_dout)
        ,.prog_we_o(_i_sbox_x8y1se__prog_we_o)
        );
    sbox_sw_N_ex_n i_sbox_x8y1sw (
        .bi_u1v1e_L1(_i_sbox_x7y0nw__so_x0y0e_L1)
        ,.so_u1y0n_L1(_i_sbox_x8y1sw__so_u1y0n_L1)
        ,.bi_x0v1w_L1(_i_sbox_x8y1se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x7y1__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x8y0nw__prog_we_o)
        ,.prog_din(_i_sbox_x8y0nw__prog_dout)
        ,.prog_dout(_i_sbox_x8y1sw__prog_dout)
        ,.prog_we_o(_i_sbox_x8y1sw__prog_we_o)
        );
    tile_clb i_tile_x8y2 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x8y2__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x8y2__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x8y2sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x7y2ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x8y2sw__prog_we_o)
        ,.prog_din(_i_sbox_x8y2sw__prog_dout)
        ,.prog_dout(_i_tile_x8y2__prog_dout)
        ,.prog_we_o(_i_tile_x8y2__prog_we_o)
        );
    sbox_ne_S_ex_w i_sbox_x8y2ne (
        .bi_x0y0e_L1(_i_sbox_x8y2nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x8y2ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x8y3ne__so_x0y0s_L1)
        ,.cu_x0y0s_L1(_i_tile_x8y2__cu_x0y0s_L1)
        ,.cv_x0y0s_L1(_i_tile_x9y2__cu_u1y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x8y3se__prog_we_o)
        ,.prog_din(_i_sbox_x8y3se__prog_dout)
        ,.prog_dout(_i_sbox_x8y2ne__prog_dout)
        ,.prog_we_o(_i_sbox_x8y2ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x8y2nw (
        .bi_u1y0n_L1(_i_sbox_x8y2sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x8y2nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x7y2nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x7y3ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x8y2__prog_we_o)
        ,.prog_din(_i_tile_x8y2__prog_dout)
        ,.prog_dout(_i_sbox_x8y2nw__prog_dout)
        ,.prog_we_o(_i_sbox_x8y2nw__prog_we_o)
        );
    sbox_se_W_ex_w i_sbox_x8y2se (
        .bi_x0v1n_L1(_i_sbox_x9y1sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x8y2se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x8y2ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x8y2ne__prog_we_o)
        ,.prog_din(_i_sbox_x8y2ne__prog_dout)
        ,.prog_dout(_i_sbox_x8y2se__prog_dout)
        ,.prog_we_o(_i_sbox_x8y2se__prog_we_o)
        );
    sbox_sw_N i_sbox_x8y2sw (
        .bi_u1v1n_L1(_i_sbox_x8y1sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x8y2sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x7y1nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x8y2se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x7y2__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x8y1nw__prog_we_o)
        ,.prog_din(_i_sbox_x8y1nw__prog_dout)
        ,.prog_dout(_i_sbox_x8y2sw__prog_dout)
        ,.prog_we_o(_i_sbox_x8y2sw__prog_we_o)
        );
    tile_clb i_tile_x8y3 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x8y3__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x8y3__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x8y3sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x7y3ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x8y3sw__prog_we_o)
        ,.prog_din(_i_sbox_x8y3sw__prog_dout)
        ,.prog_dout(_i_tile_x8y3__prog_dout)
        ,.prog_we_o(_i_tile_x8y3__prog_we_o)
        );
    sbox_ne_S_ex_w i_sbox_x8y3ne (
        .bi_x0y0e_L1(_i_sbox_x8y3nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x8y3ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x8y4ne__so_x0y0s_L1)
        ,.cu_x0y0s_L1(_i_tile_x8y3__cu_x0y0s_L1)
        ,.cv_x0y0s_L1(_i_tile_x9y3__cu_u1y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x8y4se__prog_we_o)
        ,.prog_din(_i_sbox_x8y4se__prog_dout)
        ,.prog_dout(_i_sbox_x8y3ne__prog_dout)
        ,.prog_we_o(_i_sbox_x8y3ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x8y3nw (
        .bi_u1y0n_L1(_i_sbox_x8y3sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x8y3nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x7y3nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x7y4ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x8y3__prog_we_o)
        ,.prog_din(_i_tile_x8y3__prog_dout)
        ,.prog_dout(_i_sbox_x8y3nw__prog_dout)
        ,.prog_we_o(_i_sbox_x8y3nw__prog_we_o)
        );
    sbox_se_W_ex_w i_sbox_x8y3se (
        .bi_x0v1n_L1(_i_sbox_x9y2sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x8y3se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x8y3ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x8y3ne__prog_we_o)
        ,.prog_din(_i_sbox_x8y3ne__prog_dout)
        ,.prog_dout(_i_sbox_x8y3se__prog_dout)
        ,.prog_we_o(_i_sbox_x8y3se__prog_we_o)
        );
    sbox_sw_N i_sbox_x8y3sw (
        .bi_u1v1n_L1(_i_sbox_x8y2sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x8y3sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x7y2nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x8y3se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x7y3__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x8y2nw__prog_we_o)
        ,.prog_din(_i_sbox_x8y2nw__prog_dout)
        ,.prog_dout(_i_sbox_x8y3sw__prog_dout)
        ,.prog_we_o(_i_sbox_x8y3sw__prog_we_o)
        );
    tile_clb i_tile_x8y4 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x8y4__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x8y4__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x8y4sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x7y4ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x8y4sw__prog_we_o)
        ,.prog_din(_i_sbox_x8y4sw__prog_dout)
        ,.prog_dout(_i_tile_x8y4__prog_dout)
        ,.prog_we_o(_i_tile_x8y4__prog_we_o)
        );
    sbox_ne_S_ex_w i_sbox_x8y4ne (
        .bi_x0y0e_L1(_i_sbox_x8y4nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x8y4ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x8y5ne__so_x0y0s_L1)
        ,.cu_x0y0s_L1(_i_tile_x8y4__cu_x0y0s_L1)
        ,.cv_x0y0s_L1(_i_tile_x9y4__cu_u1y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x8y5se__prog_we_o)
        ,.prog_din(_i_sbox_x8y5se__prog_dout)
        ,.prog_dout(_i_sbox_x8y4ne__prog_dout)
        ,.prog_we_o(_i_sbox_x8y4ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x8y4nw (
        .bi_u1y0n_L1(_i_sbox_x8y4sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x8y4nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x7y4nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x7y5ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x8y4__prog_we_o)
        ,.prog_din(_i_tile_x8y4__prog_dout)
        ,.prog_dout(_i_sbox_x8y4nw__prog_dout)
        ,.prog_we_o(_i_sbox_x8y4nw__prog_we_o)
        );
    sbox_se_W_ex_w i_sbox_x8y4se (
        .bi_x0v1n_L1(_i_sbox_x9y3sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x8y4se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x8y4ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x8y4ne__prog_we_o)
        ,.prog_din(_i_sbox_x8y4ne__prog_dout)
        ,.prog_dout(_i_sbox_x8y4se__prog_dout)
        ,.prog_we_o(_i_sbox_x8y4se__prog_we_o)
        );
    sbox_sw_N i_sbox_x8y4sw (
        .bi_u1v1n_L1(_i_sbox_x8y3sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x8y4sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x7y3nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x8y4se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x7y4__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x8y3nw__prog_we_o)
        ,.prog_din(_i_sbox_x8y3nw__prog_dout)
        ,.prog_dout(_i_sbox_x8y4sw__prog_dout)
        ,.prog_we_o(_i_sbox_x8y4sw__prog_we_o)
        );
    tile_clb i_tile_x8y5 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x8y5__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x8y5__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x8y5sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x7y5ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x8y5sw__prog_we_o)
        ,.prog_din(_i_sbox_x8y5sw__prog_dout)
        ,.prog_dout(_i_tile_x8y5__prog_dout)
        ,.prog_we_o(_i_tile_x8y5__prog_we_o)
        );
    sbox_ne_S_ex_w i_sbox_x8y5ne (
        .bi_x0y0e_L1(_i_sbox_x8y5nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x8y5ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x8y6ne__so_x0y0s_L1)
        ,.cu_x0y0s_L1(_i_tile_x8y5__cu_x0y0s_L1)
        ,.cv_x0y0s_L1(_i_tile_x9y5__cu_u1y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x8y6se__prog_we_o)
        ,.prog_din(_i_sbox_x8y6se__prog_dout)
        ,.prog_dout(_i_sbox_x8y5ne__prog_dout)
        ,.prog_we_o(_i_sbox_x8y5ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x8y5nw (
        .bi_u1y0n_L1(_i_sbox_x8y5sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x8y5nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x7y5nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x7y6ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x8y5__prog_we_o)
        ,.prog_din(_i_tile_x8y5__prog_dout)
        ,.prog_dout(_i_sbox_x8y5nw__prog_dout)
        ,.prog_we_o(_i_sbox_x8y5nw__prog_we_o)
        );
    sbox_se_W_ex_w i_sbox_x8y5se (
        .bi_x0v1n_L1(_i_sbox_x9y4sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x8y5se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x8y5ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x8y5ne__prog_we_o)
        ,.prog_din(_i_sbox_x8y5ne__prog_dout)
        ,.prog_dout(_i_sbox_x8y5se__prog_dout)
        ,.prog_we_o(_i_sbox_x8y5se__prog_we_o)
        );
    sbox_sw_N i_sbox_x8y5sw (
        .bi_u1v1n_L1(_i_sbox_x8y4sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x8y5sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x7y4nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x8y5se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x7y5__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x8y4nw__prog_we_o)
        ,.prog_din(_i_sbox_x8y4nw__prog_dout)
        ,.prog_dout(_i_sbox_x8y5sw__prog_dout)
        ,.prog_we_o(_i_sbox_x8y5sw__prog_we_o)
        );
    tile_clb i_tile_x8y6 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x8y6__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x8y6__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x8y6sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x7y6ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x8y6sw__prog_we_o)
        ,.prog_din(_i_sbox_x8y6sw__prog_dout)
        ,.prog_dout(_i_tile_x8y6__prog_dout)
        ,.prog_we_o(_i_tile_x8y6__prog_we_o)
        );
    sbox_ne_S_ex_w i_sbox_x8y6ne (
        .bi_x0y0e_L1(_i_sbox_x8y6nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x8y6ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x8y7ne__so_x0y0s_L1)
        ,.cu_x0y0s_L1(_i_tile_x8y6__cu_x0y0s_L1)
        ,.cv_x0y0s_L1(_i_tile_x9y6__cu_u1y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x8y7se__prog_we_o)
        ,.prog_din(_i_sbox_x8y7se__prog_dout)
        ,.prog_dout(_i_sbox_x8y6ne__prog_dout)
        ,.prog_we_o(_i_sbox_x8y6ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x8y6nw (
        .bi_u1y0n_L1(_i_sbox_x8y6sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x8y6nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x7y6nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x7y7ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x8y6__prog_we_o)
        ,.prog_din(_i_tile_x8y6__prog_dout)
        ,.prog_dout(_i_sbox_x8y6nw__prog_dout)
        ,.prog_we_o(_i_sbox_x8y6nw__prog_we_o)
        );
    sbox_se_W_ex_w i_sbox_x8y6se (
        .bi_x0v1n_L1(_i_sbox_x9y5sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x8y6se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x8y6ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x8y6ne__prog_we_o)
        ,.prog_din(_i_sbox_x8y6ne__prog_dout)
        ,.prog_dout(_i_sbox_x8y6se__prog_dout)
        ,.prog_we_o(_i_sbox_x8y6se__prog_we_o)
        );
    sbox_sw_N i_sbox_x8y6sw (
        .bi_u1v1n_L1(_i_sbox_x8y5sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x8y6sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x7y5nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x8y6se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x7y6__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x8y5nw__prog_we_o)
        ,.prog_din(_i_sbox_x8y5nw__prog_dout)
        ,.prog_dout(_i_sbox_x8y6sw__prog_dout)
        ,.prog_we_o(_i_sbox_x8y6sw__prog_we_o)
        );
    tile_clb i_tile_x8y7 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x8y7__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x8y7__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x8y7sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x7y7ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x8y7sw__prog_we_o)
        ,.prog_din(_i_sbox_x8y7sw__prog_dout)
        ,.prog_dout(_i_tile_x8y7__prog_dout)
        ,.prog_we_o(_i_tile_x8y7__prog_we_o)
        );
    sbox_ne_S_ex_w i_sbox_x8y7ne (
        .bi_x0y0e_L1(_i_sbox_x8y7nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x8y7ne__so_x0y0s_L1)
        ,.bi_x0y1s_L1(_i_sbox_x8y8ne__so_x0y0s_L1)
        ,.cu_x0y0s_L1(_i_tile_x8y7__cu_x0y0s_L1)
        ,.cv_x0y0s_L1(_i_tile_x9y7__cu_u1y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x8y8se__prog_we_o)
        ,.prog_din(_i_sbox_x8y8se__prog_dout)
        ,.prog_dout(_i_sbox_x8y7ne__prog_dout)
        ,.prog_we_o(_i_sbox_x8y7ne__prog_we_o)
        );
    sbox_nw_E i_sbox_x8y7nw (
        .bi_u1y0n_L1(_i_sbox_x8y7sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x8y7nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x7y7nw__so_x0y0e_L1)
        ,.bi_u1y1s_L1(_i_sbox_x7y8ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x8y7__prog_we_o)
        ,.prog_din(_i_tile_x8y7__prog_dout)
        ,.prog_dout(_i_sbox_x8y7nw__prog_dout)
        ,.prog_we_o(_i_sbox_x8y7nw__prog_we_o)
        );
    sbox_se_W_ex_w i_sbox_x8y7se (
        .bi_x0v1n_L1(_i_sbox_x9y6sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x8y7se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x8y7ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x8y7ne__prog_we_o)
        ,.prog_din(_i_sbox_x8y7ne__prog_dout)
        ,.prog_dout(_i_sbox_x8y7se__prog_dout)
        ,.prog_we_o(_i_sbox_x8y7se__prog_we_o)
        );
    sbox_sw_N i_sbox_x8y7sw (
        .bi_u1v1n_L1(_i_sbox_x8y6sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x8y7sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x7y6nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x8y7se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x7y7__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x8y6nw__prog_we_o)
        ,.prog_din(_i_sbox_x8y6nw__prog_dout)
        ,.prog_dout(_i_sbox_x8y7sw__prog_dout)
        ,.prog_we_o(_i_sbox_x8y7sw__prog_we_o)
        );
    tile_clb i_tile_x8y8 (
`ifdef USE_POWER_PINS
        .vssd1(vssd1),
        .vccd1(vccd1),
`endif
        .cu_x0y0n_L1(_i_tile_x8y8__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_tile_x8y8__cu_x0y0s_L1)
        ,.bi_u1y0n_L1(_i_sbox_x8y8sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x7y8ne__so_x0y0s_L1)
        ,.clk(ipin_x0y1_0)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x8y8sw__prog_we_o)
        ,.prog_din(_i_sbox_x8y8sw__prog_dout)
        ,.prog_dout(_i_tile_x8y8__prog_dout)
        ,.prog_we_o(_i_tile_x8y8__prog_we_o)
        );
    sbox_ne_S_ex_sw i_sbox_x8y8ne (
        .bi_x0y0e_L1(_i_sbox_x8y8nw__so_x0y0e_L1)
        ,.so_x0y0s_L1(_i_sbox_x8y8ne__so_x0y0s_L1)
        ,.cu_x0y0s_L1(_i_tile_x8y8__cu_x0y0s_L1)
        ,.cv_x0y0s_L1(_i_tile_x9y8__cu_u1y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x8y9se__prog_we_o)
        ,.prog_din(_i_sbox_x8y9se__prog_dout)
        ,.prog_dout(_i_sbox_x8y8ne__prog_dout)
        ,.prog_we_o(_i_sbox_x8y8ne__prog_we_o)
        );
    sbox_nw_E_ex_s i_sbox_x8y8nw (
        .bi_u1y0n_L1(_i_sbox_x8y8sw__so_u1y0n_L1)
        ,.so_x0y0e_L1(_i_sbox_x8y8nw__so_x0y0e_L1)
        ,.bi_u1y0e_L1(_i_sbox_x7y8nw__so_x0y0e_L1)
        ,.cu_x0y0e_L1(_i_tile_x8y9__cu_x0v1e_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x8y8__prog_we_o)
        ,.prog_din(_i_tile_x8y8__prog_dout)
        ,.prog_dout(_i_sbox_x8y8nw__prog_dout)
        ,.prog_we_o(_i_sbox_x8y8nw__prog_we_o)
        );
    sbox_se_W_ex_w i_sbox_x8y8se (
        .bi_x0v1n_L1(_i_sbox_x9y7sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x8y8se__so_x0v1w_L1)
        ,.bi_x0y0s_L1(_i_sbox_x8y8ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x8y8ne__prog_we_o)
        ,.prog_din(_i_sbox_x8y8ne__prog_dout)
        ,.prog_dout(_i_sbox_x8y8se__prog_dout)
        ,.prog_we_o(_i_sbox_x8y8se__prog_we_o)
        );
    sbox_sw_N i_sbox_x8y8sw (
        .bi_u1v1n_L1(_i_sbox_x8y7sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x8y8sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x7y7nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x8y8se__so_x0v1w_L1)
        ,.cu_u1y0n_L1(_i_tile_x7y8__cu_x0y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x8y7nw__prog_we_o)
        ,.prog_din(_i_sbox_x8y7nw__prog_dout)
        ,.prog_dout(_i_sbox_x8y8sw__prog_dout)
        ,.prog_we_o(_i_sbox_x8y8sw__prog_we_o)
        );
    t_io_n i_tile_x8y9 (
        .bi_x0v1e_L1(_i_sbox_x8y8nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x8y9se__so_x0v1w_L1)
        ,.cu_x0v1e_L1(_i_tile_x8y9__cu_x0v1e_L1)
        ,.cu_x0v1w_L1(_i_tile_x8y9__cu_x0v1w_L1)
        ,.ipin_x0y0_0(ipin_x8y9_0)
        ,.opin_x0y0_0(_i_tile_x8y9__opin_x0y0_0)
        ,.oe_x0y0_0(_i_tile_x8y9__oe_x0y0_0)
        ,.ipin_x0y0_1(ipin_x8y9_1)
        ,.opin_x0y0_1(_i_tile_x8y9__opin_x0y0_1)
        ,.oe_x0y0_1(_i_tile_x8y9__oe_x0y0_1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x8y8nw__prog_we_o)
        ,.prog_din(_i_sbox_x8y8nw__prog_dout)
        ,.prog_dout(_i_tile_x8y9__prog_dout)
        ,.prog_we_o(_i_tile_x8y9__prog_we_o)
        );
    sbox_se_W_ex_sw i_sbox_x8y9se (
        .bi_x0v1n_L1(_i_sbox_x9y8sw__so_u1y0n_L1)
        ,.so_x0v1w_L1(_i_sbox_x8y9se__so_x0v1w_L1)
        ,.cu_x0v1w_L1(_i_tile_x8y9__cu_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x8y9__prog_we_o)
        ,.prog_din(_i_tile_x8y9__prog_dout)
        ,.prog_dout(_i_sbox_x8y9se__prog_dout)
        ,.prog_we_o(_i_sbox_x8y9se__prog_we_o)
        );
    sbox_sw_s_ex_s i_sbox_x8y9sw (
        .bi_u1v1e_L1(_i_sbox_x7y8nw__so_x0y0e_L1)
        ,.bi_x0v1w_L1(_i_sbox_x8y9se__so_x0v1w_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_nw_w_ex_nw i_sbox_x9y0nw (
        .bi_u1y1s_L1(_i_sbox_x8y1ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    t_io_e i_tile_x9y1 (
        .bi_u1y0n_L1(_i_sbox_x9y1sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x8y1ne__so_x0y0s_L1)
        ,.cu_u1y0n_L1(_i_tile_x9y1__cu_u1y0n_L1)
        ,.cu_u1y0s_L1(_i_tile_x9y1__cu_u1y0s_L1)
        ,.ipin_x0y0_0(ipin_x9y1_0)
        ,.opin_x0y0_0(_i_tile_x9y1__opin_x0y0_0)
        ,.oe_x0y0_0(_i_tile_x9y1__oe_x0y0_0)
        ,.ipin_x0y0_1(ipin_x9y1_1)
        ,.opin_x0y0_1(_i_tile_x9y1__opin_x0y0_1)
        ,.oe_x0y0_1(_i_tile_x9y1__oe_x0y0_1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x9y1sw__prog_we_o)
        ,.prog_din(_i_sbox_x9y1sw__prog_dout)
        ,.prog_dout(_i_tile_x9y1__prog_dout)
        ,.prog_we_o(_i_tile_x9y1__prog_we_o)
        );
    sbox_nw_w_ex_w i_sbox_x9y1nw (
        .bi_u1y0n_L1(_i_sbox_x9y1sw__so_u1y0n_L1)
        ,.bi_u1y1s_L1(_i_sbox_x8y2ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_sw_N_ex_nw i_sbox_x9y1sw (
        .bi_u1v1e_L1(_i_sbox_x8y0nw__so_x0y0e_L1)
        ,.so_u1y0n_L1(_i_sbox_x9y1sw__so_u1y0n_L1)
        ,.cu_u1y0n_L1(_i_tile_x8y1__cu_x0y0n_L1)
        ,.cv_u1y0n_L1(_i_tile_x9y1__cu_u1y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_sbox_x8y1se__prog_we_o)
        ,.prog_din(_i_sbox_x8y1se__prog_dout)
        ,.prog_dout(_i_sbox_x9y1sw__prog_dout)
        ,.prog_we_o(_i_sbox_x9y1sw__prog_we_o)
        );
    t_io_e i_tile_x9y2 (
        .bi_u1y0n_L1(_i_sbox_x9y2sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x8y2ne__so_x0y0s_L1)
        ,.cu_u1y0n_L1(_i_tile_x9y2__cu_u1y0n_L1)
        ,.cu_u1y0s_L1(_i_tile_x9y2__cu_u1y0s_L1)
        ,.ipin_x0y0_0(ipin_x9y2_0)
        ,.opin_x0y0_0(_i_tile_x9y2__opin_x0y0_0)
        ,.oe_x0y0_0(_i_tile_x9y2__oe_x0y0_0)
        ,.ipin_x0y0_1(ipin_x9y2_1)
        ,.opin_x0y0_1(_i_tile_x9y2__opin_x0y0_1)
        ,.oe_x0y0_1(_i_tile_x9y2__oe_x0y0_1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x9y2sw__prog_we_o)
        ,.prog_din(_i_sbox_x9y2sw__prog_dout)
        ,.prog_dout(_i_tile_x9y2__prog_dout)
        ,.prog_we_o(_i_tile_x9y2__prog_we_o)
        );
    sbox_nw_w_ex_w i_sbox_x9y2nw (
        .bi_u1y0n_L1(_i_sbox_x9y2sw__so_u1y0n_L1)
        ,.bi_u1y1s_L1(_i_sbox_x8y3ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_sw_N_ex_w i_sbox_x9y2sw (
        .bi_u1v1n_L1(_i_sbox_x9y1sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x9y2sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x8y1nw__so_x0y0e_L1)
        ,.cu_u1y0n_L1(_i_tile_x8y2__cu_x0y0n_L1)
        ,.cv_u1y0n_L1(_i_tile_x9y2__cu_u1y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x9y1__prog_we_o)
        ,.prog_din(_i_tile_x9y1__prog_dout)
        ,.prog_dout(_i_sbox_x9y2sw__prog_dout)
        ,.prog_we_o(_i_sbox_x9y2sw__prog_we_o)
        );
    t_io_e i_tile_x9y3 (
        .bi_u1y0n_L1(_i_sbox_x9y3sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x8y3ne__so_x0y0s_L1)
        ,.cu_u1y0n_L1(_i_tile_x9y3__cu_u1y0n_L1)
        ,.cu_u1y0s_L1(_i_tile_x9y3__cu_u1y0s_L1)
        ,.ipin_x0y0_0(ipin_x9y3_0)
        ,.opin_x0y0_0(_i_tile_x9y3__opin_x0y0_0)
        ,.oe_x0y0_0(_i_tile_x9y3__oe_x0y0_0)
        ,.ipin_x0y0_1(ipin_x9y3_1)
        ,.opin_x0y0_1(_i_tile_x9y3__opin_x0y0_1)
        ,.oe_x0y0_1(_i_tile_x9y3__oe_x0y0_1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x9y3sw__prog_we_o)
        ,.prog_din(_i_sbox_x9y3sw__prog_dout)
        ,.prog_dout(_i_tile_x9y3__prog_dout)
        ,.prog_we_o(_i_tile_x9y3__prog_we_o)
        );
    sbox_nw_w_ex_w i_sbox_x9y3nw (
        .bi_u1y0n_L1(_i_sbox_x9y3sw__so_u1y0n_L1)
        ,.bi_u1y1s_L1(_i_sbox_x8y4ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_sw_N_ex_w i_sbox_x9y3sw (
        .bi_u1v1n_L1(_i_sbox_x9y2sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x9y3sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x8y2nw__so_x0y0e_L1)
        ,.cu_u1y0n_L1(_i_tile_x8y3__cu_x0y0n_L1)
        ,.cv_u1y0n_L1(_i_tile_x9y3__cu_u1y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x9y2__prog_we_o)
        ,.prog_din(_i_tile_x9y2__prog_dout)
        ,.prog_dout(_i_sbox_x9y3sw__prog_dout)
        ,.prog_we_o(_i_sbox_x9y3sw__prog_we_o)
        );
    t_io_e i_tile_x9y4 (
        .bi_u1y0n_L1(_i_sbox_x9y4sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x8y4ne__so_x0y0s_L1)
        ,.cu_u1y0n_L1(_i_tile_x9y4__cu_u1y0n_L1)
        ,.cu_u1y0s_L1(_i_tile_x9y4__cu_u1y0s_L1)
        ,.ipin_x0y0_0(ipin_x9y4_0)
        ,.opin_x0y0_0(_i_tile_x9y4__opin_x0y0_0)
        ,.oe_x0y0_0(_i_tile_x9y4__oe_x0y0_0)
        ,.ipin_x0y0_1(ipin_x9y4_1)
        ,.opin_x0y0_1(_i_tile_x9y4__opin_x0y0_1)
        ,.oe_x0y0_1(_i_tile_x9y4__oe_x0y0_1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x9y4sw__prog_we_o)
        ,.prog_din(_i_sbox_x9y4sw__prog_dout)
        ,.prog_dout(_i_tile_x9y4__prog_dout)
        ,.prog_we_o(_i_tile_x9y4__prog_we_o)
        );
    sbox_nw_w_ex_w i_sbox_x9y4nw (
        .bi_u1y0n_L1(_i_sbox_x9y4sw__so_u1y0n_L1)
        ,.bi_u1y1s_L1(_i_sbox_x8y5ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_sw_N_ex_w i_sbox_x9y4sw (
        .bi_u1v1n_L1(_i_sbox_x9y3sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x9y4sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x8y3nw__so_x0y0e_L1)
        ,.cu_u1y0n_L1(_i_tile_x8y4__cu_x0y0n_L1)
        ,.cv_u1y0n_L1(_i_tile_x9y4__cu_u1y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x9y3__prog_we_o)
        ,.prog_din(_i_tile_x9y3__prog_dout)
        ,.prog_dout(_i_sbox_x9y4sw__prog_dout)
        ,.prog_we_o(_i_sbox_x9y4sw__prog_we_o)
        );
    t_io_e i_tile_x9y5 (
        .bi_u1y0n_L1(_i_sbox_x9y5sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x8y5ne__so_x0y0s_L1)
        ,.cu_u1y0n_L1(_i_tile_x9y5__cu_u1y0n_L1)
        ,.cu_u1y0s_L1(_i_tile_x9y5__cu_u1y0s_L1)
        ,.ipin_x0y0_0(ipin_x9y5_0)
        ,.opin_x0y0_0(_i_tile_x9y5__opin_x0y0_0)
        ,.oe_x0y0_0(_i_tile_x9y5__oe_x0y0_0)
        ,.ipin_x0y0_1(ipin_x9y5_1)
        ,.opin_x0y0_1(_i_tile_x9y5__opin_x0y0_1)
        ,.oe_x0y0_1(_i_tile_x9y5__oe_x0y0_1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x9y5sw__prog_we_o)
        ,.prog_din(_i_sbox_x9y5sw__prog_dout)
        ,.prog_dout(_i_tile_x9y5__prog_dout)
        ,.prog_we_o(_i_tile_x9y5__prog_we_o)
        );
    sbox_nw_w_ex_w i_sbox_x9y5nw (
        .bi_u1y0n_L1(_i_sbox_x9y5sw__so_u1y0n_L1)
        ,.bi_u1y1s_L1(_i_sbox_x8y6ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_sw_N_ex_w i_sbox_x9y5sw (
        .bi_u1v1n_L1(_i_sbox_x9y4sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x9y5sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x8y4nw__so_x0y0e_L1)
        ,.cu_u1y0n_L1(_i_tile_x8y5__cu_x0y0n_L1)
        ,.cv_u1y0n_L1(_i_tile_x9y5__cu_u1y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x9y4__prog_we_o)
        ,.prog_din(_i_tile_x9y4__prog_dout)
        ,.prog_dout(_i_sbox_x9y5sw__prog_dout)
        ,.prog_we_o(_i_sbox_x9y5sw__prog_we_o)
        );
    t_io_e i_tile_x9y6 (
        .bi_u1y0n_L1(_i_sbox_x9y6sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x8y6ne__so_x0y0s_L1)
        ,.cu_u1y0n_L1(_i_tile_x9y6__cu_u1y0n_L1)
        ,.cu_u1y0s_L1(_i_tile_x9y6__cu_u1y0s_L1)
        ,.ipin_x0y0_0(ipin_x9y6_0)
        ,.opin_x0y0_0(_i_tile_x9y6__opin_x0y0_0)
        ,.oe_x0y0_0(_i_tile_x9y6__oe_x0y0_0)
        ,.ipin_x0y0_1(ipin_x9y6_1)
        ,.opin_x0y0_1(_i_tile_x9y6__opin_x0y0_1)
        ,.oe_x0y0_1(_i_tile_x9y6__oe_x0y0_1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x9y6sw__prog_we_o)
        ,.prog_din(_i_sbox_x9y6sw__prog_dout)
        ,.prog_dout(_i_tile_x9y6__prog_dout)
        ,.prog_we_o(_i_tile_x9y6__prog_we_o)
        );
    sbox_nw_w_ex_w i_sbox_x9y6nw (
        .bi_u1y0n_L1(_i_sbox_x9y6sw__so_u1y0n_L1)
        ,.bi_u1y1s_L1(_i_sbox_x8y7ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_sw_N_ex_w i_sbox_x9y6sw (
        .bi_u1v1n_L1(_i_sbox_x9y5sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x9y6sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x8y5nw__so_x0y0e_L1)
        ,.cu_u1y0n_L1(_i_tile_x8y6__cu_x0y0n_L1)
        ,.cv_u1y0n_L1(_i_tile_x9y6__cu_u1y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x9y5__prog_we_o)
        ,.prog_din(_i_tile_x9y5__prog_dout)
        ,.prog_dout(_i_sbox_x9y6sw__prog_dout)
        ,.prog_we_o(_i_sbox_x9y6sw__prog_we_o)
        );
    t_io_e i_tile_x9y7 (
        .bi_u1y0n_L1(_i_sbox_x9y7sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x8y7ne__so_x0y0s_L1)
        ,.cu_u1y0n_L1(_i_tile_x9y7__cu_u1y0n_L1)
        ,.cu_u1y0s_L1(_i_tile_x9y7__cu_u1y0s_L1)
        ,.ipin_x0y0_0(ipin_x9y7_0)
        ,.opin_x0y0_0(_i_tile_x9y7__opin_x0y0_0)
        ,.oe_x0y0_0(_i_tile_x9y7__oe_x0y0_0)
        ,.ipin_x0y0_1(ipin_x9y7_1)
        ,.opin_x0y0_1(_i_tile_x9y7__opin_x0y0_1)
        ,.oe_x0y0_1(_i_tile_x9y7__oe_x0y0_1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x9y7sw__prog_we_o)
        ,.prog_din(_i_sbox_x9y7sw__prog_dout)
        ,.prog_dout(_i_tile_x9y7__prog_dout)
        ,.prog_we_o(_i_tile_x9y7__prog_we_o)
        );
    sbox_nw_w_ex_w i_sbox_x9y7nw (
        .bi_u1y0n_L1(_i_sbox_x9y7sw__so_u1y0n_L1)
        ,.bi_u1y1s_L1(_i_sbox_x8y8ne__so_x0y0s_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_sw_N_ex_w i_sbox_x9y7sw (
        .bi_u1v1n_L1(_i_sbox_x9y6sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x9y7sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x8y6nw__so_x0y0e_L1)
        ,.cu_u1y0n_L1(_i_tile_x8y7__cu_x0y0n_L1)
        ,.cv_u1y0n_L1(_i_tile_x9y7__cu_u1y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x9y6__prog_we_o)
        ,.prog_din(_i_tile_x9y6__prog_dout)
        ,.prog_dout(_i_sbox_x9y7sw__prog_dout)
        ,.prog_we_o(_i_sbox_x9y7sw__prog_we_o)
        );
    t_io_e i_tile_x9y8 (
        .bi_u1y0n_L1(_i_sbox_x9y8sw__so_u1y0n_L1)
        ,.bi_u1y0s_L1(_i_sbox_x8y8ne__so_x0y0s_L1)
        ,.cu_u1y0n_L1(_i_tile_x9y8__cu_u1y0n_L1)
        ,.cu_u1y0s_L1(_i_tile_x9y8__cu_u1y0s_L1)
        ,.ipin_x0y0_0(ipin_x9y8_0)
        ,.opin_x0y0_0(_i_tile_x9y8__opin_x0y0_0)
        ,.oe_x0y0_0(_i_tile_x9y8__oe_x0y0_0)
        ,.ipin_x0y0_1(ipin_x9y8_1)
        ,.opin_x0y0_1(_i_tile_x9y8__opin_x0y0_1)
        ,.oe_x0y0_1(_i_tile_x9y8__oe_x0y0_1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l2__Q)
        ,.prog_done(_i_buf_prog_done_l2__Q)
        ,.prog_we(_i_sbox_x9y8sw__prog_we_o)
        ,.prog_din(_i_sbox_x9y8sw__prog_dout)
        ,.prog_dout(_i_tile_x9y8__prog_dout)
        ,.prog_we_o(_i_tile_x9y8__prog_we_o)
        );
    sbox_nw_w_ex_sw i_sbox_x9y8nw (
        .bi_u1y0n_L1(_i_sbox_x9y8sw__so_u1y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    sbox_sw_N_ex_w i_sbox_x9y8sw (
        .bi_u1v1n_L1(_i_sbox_x9y7sw__so_u1y0n_L1)
        ,.so_u1y0n_L1(_i_sbox_x9y8sw__so_u1y0n_L1)
        ,.bi_u1v1e_L1(_i_sbox_x8y7nw__so_x0y0e_L1)
        ,.cu_u1y0n_L1(_i_tile_x8y8__cu_x0y0n_L1)
        ,.cv_u1y0n_L1(_i_tile_x9y8__cu_u1y0n_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_tile_x9y7__prog_we_o)
        ,.prog_din(_i_tile_x9y7__prog_dout)
        ,.prog_dout(_i_sbox_x9y8sw__prog_dout)
        ,.prog_we_o(_i_sbox_x9y8sw__prog_we_o)
        );
    sbox_sw_s_ex_sw i_sbox_x9y9sw (
        .bi_u1v1e_L1(_i_sbox_x8y8nw__so_x0y0e_L1)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(_i_buf_prog_rst_l1__Q)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(_i_buf_prog_done_l1__Q)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    prga_simple_buf i_buf_prog_rst_l1 (
        .C(prog_clk)
        ,.D(_i_buf_prog_rst_l2__Q)
        ,.Q(_i_buf_prog_rst_l1__Q)
        );
    prga_simple_bufr i_buf_prog_done_l1 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(_i_buf_prog_done_l2__Q)
        ,.Q(_i_buf_prog_done_l1__Q)
        );
    prga_simple_buf i_buf_prog_rst_l2 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l2__Q)
        );
    prga_simple_bufr i_buf_prog_done_l2 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l2__Q)
        );
        
    assign opin_x0y1_0 = _i_tile_x0y1__opin_x0y0_0;
    assign oe_x0y1_0 = _i_tile_x0y1__oe_x0y0_0;
    assign opin_x0y1_1 = _i_tile_x0y1__opin_x0y0_1;
    assign oe_x0y1_1 = _i_tile_x0y1__oe_x0y0_1;
    assign opin_x0y2_0 = _i_tile_x0y2__opin_x0y0_0;
    assign oe_x0y2_0 = _i_tile_x0y2__oe_x0y0_0;
    assign opin_x0y2_1 = _i_tile_x0y2__opin_x0y0_1;
    assign oe_x0y2_1 = _i_tile_x0y2__oe_x0y0_1;
    assign opin_x0y3_0 = _i_tile_x0y3__opin_x0y0_0;
    assign oe_x0y3_0 = _i_tile_x0y3__oe_x0y0_0;
    assign opin_x0y3_1 = _i_tile_x0y3__opin_x0y0_1;
    assign oe_x0y3_1 = _i_tile_x0y3__oe_x0y0_1;
    assign opin_x0y4_0 = _i_tile_x0y4__opin_x0y0_0;
    assign oe_x0y4_0 = _i_tile_x0y4__oe_x0y0_0;
    assign opin_x0y4_1 = _i_tile_x0y4__opin_x0y0_1;
    assign oe_x0y4_1 = _i_tile_x0y4__oe_x0y0_1;
    assign opin_x0y5_0 = _i_tile_x0y5__opin_x0y0_0;
    assign oe_x0y5_0 = _i_tile_x0y5__oe_x0y0_0;
    assign opin_x0y5_1 = _i_tile_x0y5__opin_x0y0_1;
    assign oe_x0y5_1 = _i_tile_x0y5__oe_x0y0_1;
    assign opin_x0y6_0 = _i_tile_x0y6__opin_x0y0_0;
    assign oe_x0y6_0 = _i_tile_x0y6__oe_x0y0_0;
    assign opin_x0y6_1 = _i_tile_x0y6__opin_x0y0_1;
    assign oe_x0y6_1 = _i_tile_x0y6__oe_x0y0_1;
    assign opin_x0y7_0 = _i_tile_x0y7__opin_x0y0_0;
    assign oe_x0y7_0 = _i_tile_x0y7__oe_x0y0_0;
    assign opin_x0y7_1 = _i_tile_x0y7__opin_x0y0_1;
    assign oe_x0y7_1 = _i_tile_x0y7__oe_x0y0_1;
    assign opin_x0y8_0 = _i_tile_x0y8__opin_x0y0_0;
    assign oe_x0y8_0 = _i_tile_x0y8__oe_x0y0_0;
    assign opin_x0y8_1 = _i_tile_x0y8__opin_x0y0_1;
    assign oe_x0y8_1 = _i_tile_x0y8__oe_x0y0_1;
    assign opin_x1y9_0 = _i_tile_x1y9__opin_x0y0_0;
    assign oe_x1y9_0 = _i_tile_x1y9__oe_x0y0_0;
    assign opin_x1y9_1 = _i_tile_x1y9__opin_x0y0_1;
    assign oe_x1y9_1 = _i_tile_x1y9__oe_x0y0_1;
    assign opin_x2y9_0 = _i_tile_x2y9__opin_x0y0_0;
    assign oe_x2y9_0 = _i_tile_x2y9__oe_x0y0_0;
    assign opin_x2y9_1 = _i_tile_x2y9__opin_x0y0_1;
    assign oe_x2y9_1 = _i_tile_x2y9__oe_x0y0_1;
    assign opin_x3y9_0 = _i_tile_x3y9__opin_x0y0_0;
    assign oe_x3y9_0 = _i_tile_x3y9__oe_x0y0_0;
    assign opin_x3y9_1 = _i_tile_x3y9__opin_x0y0_1;
    assign oe_x3y9_1 = _i_tile_x3y9__oe_x0y0_1;
    assign opin_x4y9_0 = _i_tile_x4y9__opin_x0y0_0;
    assign oe_x4y9_0 = _i_tile_x4y9__oe_x0y0_0;
    assign opin_x4y9_1 = _i_tile_x4y9__opin_x0y0_1;
    assign oe_x4y9_1 = _i_tile_x4y9__oe_x0y0_1;
    assign opin_x5y9_0 = _i_tile_x5y9__opin_x0y0_0;
    assign oe_x5y9_0 = _i_tile_x5y9__oe_x0y0_0;
    assign opin_x5y9_1 = _i_tile_x5y9__opin_x0y0_1;
    assign oe_x5y9_1 = _i_tile_x5y9__oe_x0y0_1;
    assign opin_x6y9_0 = _i_tile_x6y9__opin_x0y0_0;
    assign oe_x6y9_0 = _i_tile_x6y9__oe_x0y0_0;
    assign opin_x6y9_1 = _i_tile_x6y9__opin_x0y0_1;
    assign oe_x6y9_1 = _i_tile_x6y9__oe_x0y0_1;
    assign opin_x7y9_0 = _i_tile_x7y9__opin_x0y0_0;
    assign oe_x7y9_0 = _i_tile_x7y9__oe_x0y0_0;
    assign opin_x7y9_1 = _i_tile_x7y9__opin_x0y0_1;
    assign oe_x7y9_1 = _i_tile_x7y9__oe_x0y0_1;
    assign opin_x8y9_0 = _i_tile_x8y9__opin_x0y0_0;
    assign oe_x8y9_0 = _i_tile_x8y9__oe_x0y0_0;
    assign opin_x8y9_1 = _i_tile_x8y9__opin_x0y0_1;
    assign oe_x8y9_1 = _i_tile_x8y9__oe_x0y0_1;
    assign opin_x9y1_0 = _i_tile_x9y1__opin_x0y0_0;
    assign oe_x9y1_0 = _i_tile_x9y1__oe_x0y0_0;
    assign opin_x9y1_1 = _i_tile_x9y1__opin_x0y0_1;
    assign oe_x9y1_1 = _i_tile_x9y1__oe_x0y0_1;
    assign opin_x9y2_0 = _i_tile_x9y2__opin_x0y0_0;
    assign oe_x9y2_0 = _i_tile_x9y2__oe_x0y0_0;
    assign opin_x9y2_1 = _i_tile_x9y2__opin_x0y0_1;
    assign oe_x9y2_1 = _i_tile_x9y2__oe_x0y0_1;
    assign opin_x9y3_0 = _i_tile_x9y3__opin_x0y0_0;
    assign oe_x9y3_0 = _i_tile_x9y3__oe_x0y0_0;
    assign opin_x9y3_1 = _i_tile_x9y3__opin_x0y0_1;
    assign oe_x9y3_1 = _i_tile_x9y3__oe_x0y0_1;
    assign opin_x9y4_0 = _i_tile_x9y4__opin_x0y0_0;
    assign oe_x9y4_0 = _i_tile_x9y4__oe_x0y0_0;
    assign opin_x9y4_1 = _i_tile_x9y4__opin_x0y0_1;
    assign oe_x9y4_1 = _i_tile_x9y4__oe_x0y0_1;
    assign opin_x9y5_0 = _i_tile_x9y5__opin_x0y0_0;
    assign oe_x9y5_0 = _i_tile_x9y5__oe_x0y0_0;
    assign opin_x9y5_1 = _i_tile_x9y5__opin_x0y0_1;
    assign oe_x9y5_1 = _i_tile_x9y5__oe_x0y0_1;
    assign opin_x9y6_0 = _i_tile_x9y6__opin_x0y0_0;
    assign oe_x9y6_0 = _i_tile_x9y6__oe_x0y0_0;
    assign opin_x9y6_1 = _i_tile_x9y6__opin_x0y0_1;
    assign oe_x9y6_1 = _i_tile_x9y6__oe_x0y0_1;
    assign opin_x9y7_0 = _i_tile_x9y7__opin_x0y0_0;
    assign oe_x9y7_0 = _i_tile_x9y7__oe_x0y0_0;
    assign opin_x9y7_1 = _i_tile_x9y7__opin_x0y0_1;
    assign oe_x9y7_1 = _i_tile_x9y7__oe_x0y0_1;
    assign opin_x9y8_0 = _i_tile_x9y8__opin_x0y0_0;
    assign oe_x9y8_0 = _i_tile_x9y8__oe_x0y0_0;
    assign opin_x9y8_1 = _i_tile_x9y8__opin_x0y0_1;
    assign oe_x9y8_1 = _i_tile_x9y8__oe_x0y0_1;
    assign prog_dout = _i_tile_x9y8__prog_dout;
    assign prog_we_o = _i_tile_x9y8__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_ne_n_ex_ne (
    input wire [11:0] bi_x1y0w_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    );
    
        
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
        
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
        

endmodule
// Automatically generated by PRGA's RTL generator
module t_io_w (
    input wire [11:0] bi_x0y0n_L1
    , input wire [11:0] bi_x0y0s_L1
    , output wire [11:0] cu_x0y0n_L1
    , output wire [11:0] cu_x0y0s_L1
    , input wire [0:0] ipin_x0y0_0
    , output wire [0:0] opin_x0y0_0
    , output wire [0:0] oe_x0y0_0
    , input wire [0:0] ipin_x0y0_1
    , output wire [0:0] opin_x0y0_1
    , output wire [0:0] oe_x0y0_1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_blk_i0__inpad;
    wire [0:0] _i_blk_i0__opin;
    wire [0:0] _i_blk_i0__oe;
    wire [0:0] _i_blk_i0__prog_dout;
    wire [0:0] _i_blk_i0__prog_we_o;
    wire [0:0] _i_blk_i1__inpad;
    wire [0:0] _i_blk_i1__opin;
    wire [0:0] _i_blk_i1__oe;
    wire [0:0] _i_blk_i1__prog_dout;
    wire [0:0] _i_blk_i1__prog_we_o;
    wire [0:0] _i_cbox_e0__bp_x0y0i0_outpad;
    wire [11:0] _i_cbox_e0__cu_x0y0n_L1;
    wire [11:0] _i_cbox_e0__cu_x0y0s_L1;
    wire [0:0] _i_cbox_e0__bp_x0y0i1_outpad;
    wire [0:0] _i_cbox_e0__prog_dout;
    wire [0:0] _i_cbox_e0__prog_we_o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_buf_prog_rst_l1__Q;
    wire [0:0] _i_buf_prog_done_l1__Q;
        
    iob i_blk_i0 (
        .outpad(_i_cbox_e0__bp_x0y0i0_outpad)
        ,.inpad(_i_blk_i0__inpad)
        ,.ipin(ipin_x0y0_0)
        ,.opin(_i_blk_i0__opin)
        ,.oe(_i_blk_i0__oe)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_blk_i0__prog_dout)
        ,.prog_we_o(_i_blk_i0__prog_we_o)
        );
    iob i_blk_i1 (
        .outpad(_i_cbox_e0__bp_x0y0i1_outpad)
        ,.inpad(_i_blk_i1__inpad)
        ,.ipin(ipin_x0y0_1)
        ,.opin(_i_blk_i1__opin)
        ,.oe(_i_blk_i1__oe)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_blk_i0__prog_we_o)
        ,.prog_din(_i_blk_i0__prog_dout)
        ,.prog_dout(_i_blk_i1__prog_dout)
        ,.prog_we_o(_i_blk_i1__prog_we_o)
        );
    cbox_t_io_w_e0 i_cbox_e0 (
        .bp_x0y0i0_outpad(_i_cbox_e0__bp_x0y0i0_outpad)
        ,.bi_x0y0n_L1(bi_x0y0n_L1)
        ,.bi_x0y0s_L1(bi_x0y0s_L1)
        ,.bp_x0y0i0_inpad(_i_blk_i0__inpad)
        ,.cu_x0y0n_L1(_i_cbox_e0__cu_x0y0n_L1)
        ,.cu_x0y0s_L1(_i_cbox_e0__cu_x0y0s_L1)
        ,.bp_x0y0i1_outpad(_i_cbox_e0__bp_x0y0i1_outpad)
        ,.bp_x0y0i1_inpad(_i_blk_i1__inpad)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_blk_i1__prog_we_o)
        ,.prog_din(_i_blk_i1__prog_dout)
        ,.prog_dout(_i_cbox_e0__prog_dout)
        ,.prog_we_o(_i_cbox_e0__prog_we_o)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(_i_buf_prog_rst_l1__Q)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(_i_buf_prog_done_l1__Q)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    prga_simple_buf i_buf_prog_rst_l1 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l1__Q)
        );
    prga_simple_bufr i_buf_prog_done_l1 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l1__Q)
        );
        
    assign cu_x0y0n_L1 = _i_cbox_e0__cu_x0y0n_L1;
    assign cu_x0y0s_L1 = _i_cbox_e0__cu_x0y0s_L1;
    assign opin_x0y0_0 = _i_blk_i0__opin;
    assign oe_x0y0_0 = _i_blk_i0__oe;
    assign opin_x0y0_1 = _i_blk_i1__opin;
    assign oe_x0y0_1 = _i_blk_i1__oe;
    assign prog_dout = _i_cbox_e0__prog_dout;
    assign prog_we_o = _i_cbox_e0__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_ne_S_ex_e (
    input wire [11:0] bi_x0y1s_L1
    , output wire [11:0] so_x0y0s_L1
    , input wire [11:0] bi_x1y0w_L1
    , input wire [11:0] cu_x0y0s_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_so_x0y0s_L1_0__o;
    wire [0:0] _i_sw_so_x0y0s_L1_1__o;
    wire [0:0] _i_sw_so_x0y0s_L1_2__o;
    wire [0:0] _i_sw_so_x0y0s_L1_3__o;
    wire [0:0] _i_sw_so_x0y0s_L1_4__o;
    wire [0:0] _i_sw_so_x0y0s_L1_5__o;
    wire [0:0] _i_sw_so_x0y0s_L1_6__o;
    wire [0:0] _i_sw_so_x0y0s_L1_7__o;
    wire [0:0] _i_sw_so_x0y0s_L1_8__o;
    wire [0:0] _i_sw_so_x0y0s_L1_9__o;
    wire [0:0] _i_sw_so_x0y0s_L1_10__o;
    wire [0:0] _i_sw_so_x0y0s_L1_11__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_4__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_4__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_5__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_5__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_6__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_7__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_8__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_9__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_9__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_10__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_10__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_11__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_11__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw3 i_sw_so_x0y0s_L1_0 (
        .i({cu_x0y0s_L1[0],
            bi_x1y0w_L1[0],
            bi_x0y1s_L1[0]})
        ,.o(_i_sw_so_x0y0s_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_0__prog_data)
        );
    sw2 i_sw_so_x0y0s_L1_1 (
        .i({cu_x0y0s_L1[1],
            bi_x0y1s_L1[1]})
        ,.o(_i_sw_so_x0y0s_L1_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_1__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_2 (
        .i({cu_x0y0s_L1[2],
            bi_x1y0w_L1[2],
            bi_x0y1s_L1[2]})
        ,.o(_i_sw_so_x0y0s_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_2__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_3 (
        .i({cu_x0y0s_L1[3],
            bi_x1y0w_L1[3],
            bi_x0y1s_L1[3]})
        ,.o(_i_sw_so_x0y0s_L1_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_3__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_4 (
        .i({cu_x0y0s_L1[4],
            bi_x1y0w_L1[4],
            bi_x0y1s_L1[4]})
        ,.o(_i_sw_so_x0y0s_L1_4__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_4__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_5 (
        .i({cu_x0y0s_L1[5],
            bi_x1y0w_L1[5],
            bi_x0y1s_L1[5]})
        ,.o(_i_sw_so_x0y0s_L1_5__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_5__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_6 (
        .i({cu_x0y0s_L1[6],
            bi_x1y0w_L1[6],
            bi_x0y1s_L1[6]})
        ,.o(_i_sw_so_x0y0s_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_6__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_7 (
        .i({cu_x0y0s_L1[7],
            bi_x1y0w_L1[7],
            bi_x0y1s_L1[7]})
        ,.o(_i_sw_so_x0y0s_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_7__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_8 (
        .i({cu_x0y0s_L1[8],
            bi_x1y0w_L1[8],
            bi_x0y1s_L1[8]})
        ,.o(_i_sw_so_x0y0s_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_8__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_9 (
        .i({cu_x0y0s_L1[9],
            bi_x1y0w_L1[9],
            bi_x0y1s_L1[9]})
        ,.o(_i_sw_so_x0y0s_L1_9__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_9__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_10 (
        .i({cu_x0y0s_L1[10],
            bi_x1y0w_L1[10],
            bi_x0y1s_L1[10]})
        ,.o(_i_sw_so_x0y0s_L1_10__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_10__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_11 (
        .i({cu_x0y0s_L1[11],
            bi_x1y0w_L1[11],
            bi_x0y1s_L1[11]})
        ,.o(_i_sw_so_x0y0s_L1_11__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_11__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_3__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_4 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_4__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_4__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_5 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_4__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_5__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_5__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_5__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_6__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_7__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_8__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_9 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_9__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_9__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_10 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_9__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_10__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_10__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_11 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_10__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_11__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_11__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_11__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign so_x0y0s_L1 = {_i_sw_so_x0y0s_L1_11__o,
        _i_sw_so_x0y0s_L1_10__o,
        _i_sw_so_x0y0s_L1_9__o,
        _i_sw_so_x0y0s_L1_8__o,
        _i_sw_so_x0y0s_L1_7__o,
        _i_sw_so_x0y0s_L1_6__o,
        _i_sw_so_x0y0s_L1_5__o,
        _i_sw_so_x0y0s_L1_4__o,
        _i_sw_so_x0y0s_L1_3__o,
        _i_sw_so_x0y0s_L1_2__o,
        _i_sw_so_x0y0s_L1_1__o,
        _i_sw_so_x0y0s_L1_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_se_e_ex_ne (
    input wire [11:0] bi_x0y0s_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    );
    
        
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
        
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
        

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_se_e_ex_e (
    input wire [11:0] bi_x0v1n_L1
    , input wire [11:0] bi_x0y0s_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    );
    
        
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
        
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
        

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_ne_S_ex_es (
    input wire [11:0] bi_x1y0w_L1
    , output wire [11:0] so_x0y0s_L1
    , input wire [11:0] cu_x0y0s_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_so_x0y0s_L1_0__o;
    wire [0:0] _i_sw_so_x0y0s_L1_1__o;
    wire [0:0] _i_sw_so_x0y0s_L1_2__o;
    wire [0:0] _i_sw_so_x0y0s_L1_3__o;
    wire [0:0] _i_sw_so_x0y0s_L1_4__o;
    wire [0:0] _i_sw_so_x0y0s_L1_5__o;
    wire [0:0] _i_sw_so_x0y0s_L1_6__o;
    wire [0:0] _i_sw_so_x0y0s_L1_7__o;
    wire [0:0] _i_sw_so_x0y0s_L1_8__o;
    wire [0:0] _i_sw_so_x0y0s_L1_9__o;
    wire [0:0] _i_sw_so_x0y0s_L1_10__o;
    wire [0:0] _i_sw_so_x0y0s_L1_11__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_1__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_4__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_4__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_5__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_5__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_6__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_7__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_8__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_9__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_9__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_10__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_10__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_11__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_11__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw2 i_sw_so_x0y0s_L1_0 (
        .i({cu_x0y0s_L1[0],
            bi_x1y0w_L1[0]})
        ,.o(_i_sw_so_x0y0s_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_0__prog_data)
        );
    sw1 i_sw_so_x0y0s_L1_1 (
        .i(cu_x0y0s_L1[1])
        ,.o(_i_sw_so_x0y0s_L1_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_1__prog_data)
        );
    sw2 i_sw_so_x0y0s_L1_2 (
        .i({cu_x0y0s_L1[2],
            bi_x1y0w_L1[2]})
        ,.o(_i_sw_so_x0y0s_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_2__prog_data)
        );
    sw2 i_sw_so_x0y0s_L1_3 (
        .i({cu_x0y0s_L1[3],
            bi_x1y0w_L1[3]})
        ,.o(_i_sw_so_x0y0s_L1_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_3__prog_data)
        );
    sw2 i_sw_so_x0y0s_L1_4 (
        .i({cu_x0y0s_L1[4],
            bi_x1y0w_L1[4]})
        ,.o(_i_sw_so_x0y0s_L1_4__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_4__prog_data)
        );
    sw2 i_sw_so_x0y0s_L1_5 (
        .i({cu_x0y0s_L1[5],
            bi_x1y0w_L1[5]})
        ,.o(_i_sw_so_x0y0s_L1_5__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_5__prog_data)
        );
    sw2 i_sw_so_x0y0s_L1_6 (
        .i({cu_x0y0s_L1[6],
            bi_x1y0w_L1[6]})
        ,.o(_i_sw_so_x0y0s_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_6__prog_data)
        );
    sw2 i_sw_so_x0y0s_L1_7 (
        .i({cu_x0y0s_L1[7],
            bi_x1y0w_L1[7]})
        ,.o(_i_sw_so_x0y0s_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_7__prog_data)
        );
    sw2 i_sw_so_x0y0s_L1_8 (
        .i({cu_x0y0s_L1[8],
            bi_x1y0w_L1[8]})
        ,.o(_i_sw_so_x0y0s_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_8__prog_data)
        );
    sw2 i_sw_so_x0y0s_L1_9 (
        .i({cu_x0y0s_L1[9],
            bi_x1y0w_L1[9]})
        ,.o(_i_sw_so_x0y0s_L1_9__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_9__prog_data)
        );
    sw2 i_sw_so_x0y0s_L1_10 (
        .i({cu_x0y0s_L1[10],
            bi_x1y0w_L1[10]})
        ,.o(_i_sw_so_x0y0s_L1_10__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_10__prog_data)
        );
    sw2 i_sw_so_x0y0s_L1_11 (
        .i({cu_x0y0s_L1[11],
            bi_x1y0w_L1[11]})
        ,.o(_i_sw_so_x0y0s_L1_11__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_11__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_0__prog_data)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0y0s_L1_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_3__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_4 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_4__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_4__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_5 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_4__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_5__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_5__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_5__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_6__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_7__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_8__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_9 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_9__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_9__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_10 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_9__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_10__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_10__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_11 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_10__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_11__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_11__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_11__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign so_x0y0s_L1 = {_i_sw_so_x0y0s_L1_11__o,
        _i_sw_so_x0y0s_L1_10__o,
        _i_sw_so_x0y0s_L1_9__o,
        _i_sw_so_x0y0s_L1_8__o,
        _i_sw_so_x0y0s_L1_7__o,
        _i_sw_so_x0y0s_L1_6__o,
        _i_sw_so_x0y0s_L1_5__o,
        _i_sw_so_x0y0s_L1_4__o,
        _i_sw_so_x0y0s_L1_3__o,
        _i_sw_so_x0y0s_L1_2__o,
        _i_sw_so_x0y0s_L1_1__o,
        _i_sw_so_x0y0s_L1_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_se_e_ex_es (
    input wire [11:0] bi_x0v1n_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    );
    
        
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
        
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
        

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_ne_n_ex_n (
    input wire [11:0] bi_x0y0e_L1
    , input wire [11:0] bi_x1y0w_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    );
    
        
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
        
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
        

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_nw_E_ex_ne (
    input wire [11:0] bi_u1y1s_L1
    , output wire [11:0] so_x0y0e_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_so_x0y0e_L1_0__o;
    wire [0:0] _i_sw_so_x0y0e_L1_1__o;
    wire [0:0] _i_sw_so_x0y0e_L1_2__o;
    wire [0:0] _i_sw_so_x0y0e_L1_3__o;
    wire [0:0] _i_sw_so_x0y0e_L1_4__o;
    wire [0:0] _i_sw_so_x0y0e_L1_5__o;
    wire [0:0] _i_sw_so_x0y0e_L1_6__o;
    wire [0:0] _i_sw_so_x0y0e_L1_7__o;
    wire [0:0] _i_sw_so_x0y0e_L1_8__o;
    wire [0:0] _i_sw_so_x0y0e_L1_9__o;
    wire [0:0] _i_sw_so_x0y0e_L1_10__o;
    wire [0:0] _i_sw_so_x0y0e_L1_11__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_0__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_1__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_2__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_3__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_4__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_4__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_5__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_5__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_6__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_7__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_8__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_9__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_9__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_10__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_10__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_11__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_11__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw1 i_sw_so_x0y0e_L1_0 (
        .i(bi_u1y1s_L1[1])
        ,.o(_i_sw_so_x0y0e_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_0__prog_data)
        );
    sw1 i_sw_so_x0y0e_L1_1 (
        .i(bi_u1y1s_L1[2])
        ,.o(_i_sw_so_x0y0e_L1_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_1__prog_data)
        );
    sw1 i_sw_so_x0y0e_L1_2 (
        .i(bi_u1y1s_L1[3])
        ,.o(_i_sw_so_x0y0e_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_2__prog_data)
        );
    sw1 i_sw_so_x0y0e_L1_3 (
        .i(bi_u1y1s_L1[4])
        ,.o(_i_sw_so_x0y0e_L1_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_3__prog_data)
        );
    sw1 i_sw_so_x0y0e_L1_4 (
        .i(bi_u1y1s_L1[5])
        ,.o(_i_sw_so_x0y0e_L1_4__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_4__prog_data)
        );
    sw1 i_sw_so_x0y0e_L1_5 (
        .i(bi_u1y1s_L1[6])
        ,.o(_i_sw_so_x0y0e_L1_5__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_5__prog_data)
        );
    sw1 i_sw_so_x0y0e_L1_6 (
        .i(bi_u1y1s_L1[7])
        ,.o(_i_sw_so_x0y0e_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_6__prog_data)
        );
    sw1 i_sw_so_x0y0e_L1_7 (
        .i(bi_u1y1s_L1[8])
        ,.o(_i_sw_so_x0y0e_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_7__prog_data)
        );
    sw1 i_sw_so_x0y0e_L1_8 (
        .i(bi_u1y1s_L1[9])
        ,.o(_i_sw_so_x0y0e_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_8__prog_data)
        );
    sw1 i_sw_so_x0y0e_L1_9 (
        .i(bi_u1y1s_L1[10])
        ,.o(_i_sw_so_x0y0e_L1_9__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_9__prog_data)
        );
    sw1 i_sw_so_x0y0e_L1_10 (
        .i(bi_u1y1s_L1[11])
        ,.o(_i_sw_so_x0y0e_L1_10__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_10__prog_data)
        );
    sw1 i_sw_so_x0y0e_L1_11 (
        .i(bi_u1y1s_L1[0])
        ,.o(_i_sw_so_x0y0e_L1_11__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_11__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0y0e_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_0__prog_data)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0y0e_L1_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_1__prog_data)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0y0e_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_2__prog_data)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0y0e_L1_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_3__prog_data)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0y0e_L1_4 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_4__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_4__prog_data)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0y0e_L1_5 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_4__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_5__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_5__prog_data)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0y0e_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_5__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_6__prog_data)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0y0e_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_7__prog_data)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0y0e_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_8__prog_data)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0y0e_L1_9 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_9__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_9__prog_data)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0y0e_L1_10 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_9__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_10__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_10__prog_data)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0y0e_L1_11 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_10__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_11__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_11__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_11__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign so_x0y0e_L1 = {_i_sw_so_x0y0e_L1_11__o,
        _i_sw_so_x0y0e_L1_10__o,
        _i_sw_so_x0y0e_L1_9__o,
        _i_sw_so_x0y0e_L1_8__o,
        _i_sw_so_x0y0e_L1_7__o,
        _i_sw_so_x0y0e_L1_6__o,
        _i_sw_so_x0y0e_L1_5__o,
        _i_sw_so_x0y0e_L1_4__o,
        _i_sw_so_x0y0e_L1_3__o,
        _i_sw_so_x0y0e_L1_2__o,
        _i_sw_so_x0y0e_L1_1__o,
        _i_sw_so_x0y0e_L1_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_ne_S (
    input wire [11:0] bi_x0y0e_L1
    , output wire [11:0] so_x0y0s_L1
    , input wire [11:0] bi_x0y1s_L1
    , input wire [11:0] bi_x1y0w_L1
    , input wire [11:0] cu_x0y0s_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_so_x0y0s_L1_0__o;
    wire [0:0] _i_sw_so_x0y0s_L1_1__o;
    wire [0:0] _i_sw_so_x0y0s_L1_2__o;
    wire [0:0] _i_sw_so_x0y0s_L1_3__o;
    wire [0:0] _i_sw_so_x0y0s_L1_4__o;
    wire [0:0] _i_sw_so_x0y0s_L1_5__o;
    wire [0:0] _i_sw_so_x0y0s_L1_6__o;
    wire [0:0] _i_sw_so_x0y0s_L1_7__o;
    wire [0:0] _i_sw_so_x0y0s_L1_8__o;
    wire [0:0] _i_sw_so_x0y0s_L1_9__o;
    wire [0:0] _i_sw_so_x0y0s_L1_10__o;
    wire [0:0] _i_sw_so_x0y0s_L1_11__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_0__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_x0y0s_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_2__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_x0y0s_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_3__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_x0y0s_L1_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_4__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_x0y0s_L1_4__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_5__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_x0y0s_L1_5__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_6__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_x0y0s_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_7__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_x0y0s_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_8__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_x0y0s_L1_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_9__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_x0y0s_L1_9__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_10__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_x0y0s_L1_10__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_11__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_x0y0s_L1_11__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw4 i_sw_so_x0y0s_L1_0 (
        .i({cu_x0y0s_L1[0],
            bi_x1y0w_L1[0],
            bi_x0y1s_L1[0],
            bi_x0y0e_L1[11]})
        ,.o(_i_sw_so_x0y0s_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_0__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_1 (
        .i({cu_x0y0s_L1[1],
            bi_x0y1s_L1[1],
            bi_x0y0e_L1[0]})
        ,.o(_i_sw_so_x0y0s_L1_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_1__prog_data)
        );
    sw4 i_sw_so_x0y0s_L1_2 (
        .i({cu_x0y0s_L1[2],
            bi_x1y0w_L1[2],
            bi_x0y1s_L1[2],
            bi_x0y0e_L1[1]})
        ,.o(_i_sw_so_x0y0s_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_2__prog_data)
        );
    sw4 i_sw_so_x0y0s_L1_3 (
        .i({cu_x0y0s_L1[3],
            bi_x1y0w_L1[3],
            bi_x0y1s_L1[3],
            bi_x0y0e_L1[2]})
        ,.o(_i_sw_so_x0y0s_L1_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_3__prog_data)
        );
    sw4 i_sw_so_x0y0s_L1_4 (
        .i({cu_x0y0s_L1[4],
            bi_x1y0w_L1[4],
            bi_x0y1s_L1[4],
            bi_x0y0e_L1[3]})
        ,.o(_i_sw_so_x0y0s_L1_4__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_4__prog_data)
        );
    sw4 i_sw_so_x0y0s_L1_5 (
        .i({cu_x0y0s_L1[5],
            bi_x1y0w_L1[5],
            bi_x0y1s_L1[5],
            bi_x0y0e_L1[4]})
        ,.o(_i_sw_so_x0y0s_L1_5__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_5__prog_data)
        );
    sw4 i_sw_so_x0y0s_L1_6 (
        .i({cu_x0y0s_L1[6],
            bi_x1y0w_L1[6],
            bi_x0y1s_L1[6],
            bi_x0y0e_L1[5]})
        ,.o(_i_sw_so_x0y0s_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_6__prog_data)
        );
    sw4 i_sw_so_x0y0s_L1_7 (
        .i({cu_x0y0s_L1[7],
            bi_x1y0w_L1[7],
            bi_x0y1s_L1[7],
            bi_x0y0e_L1[6]})
        ,.o(_i_sw_so_x0y0s_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_7__prog_data)
        );
    sw4 i_sw_so_x0y0s_L1_8 (
        .i({cu_x0y0s_L1[8],
            bi_x1y0w_L1[8],
            bi_x0y1s_L1[8],
            bi_x0y0e_L1[7]})
        ,.o(_i_sw_so_x0y0s_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_8__prog_data)
        );
    sw4 i_sw_so_x0y0s_L1_9 (
        .i({cu_x0y0s_L1[9],
            bi_x1y0w_L1[9],
            bi_x0y1s_L1[9],
            bi_x0y0e_L1[8]})
        ,.o(_i_sw_so_x0y0s_L1_9__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_9__prog_data)
        );
    sw4 i_sw_so_x0y0s_L1_10 (
        .i({cu_x0y0s_L1[10],
            bi_x1y0w_L1[10],
            bi_x0y1s_L1[10],
            bi_x0y0e_L1[9]})
        ,.o(_i_sw_so_x0y0s_L1_10__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_10__prog_data)
        );
    sw4 i_sw_so_x0y0s_L1_11 (
        .i({cu_x0y0s_L1[11],
            bi_x1y0w_L1[11],
            bi_x0y1s_L1[11],
            bi_x0y0e_L1[10]})
        ,.o(_i_sw_so_x0y0s_L1_11__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_11__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_x0y0s_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_1__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_x0y0s_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_2__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_x0y0s_L1_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_3__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_x0y0s_L1_4 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_4__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_4__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_x0y0s_L1_5 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_4__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_5__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_5__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_x0y0s_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_5__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_6__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_x0y0s_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_7__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_x0y0s_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_8__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_x0y0s_L1_9 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_9__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_9__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_x0y0s_L1_10 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_9__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_10__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_10__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_x0y0s_L1_11 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_10__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_11__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_11__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_11__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign so_x0y0s_L1 = {_i_sw_so_x0y0s_L1_11__o,
        _i_sw_so_x0y0s_L1_10__o,
        _i_sw_so_x0y0s_L1_9__o,
        _i_sw_so_x0y0s_L1_8__o,
        _i_sw_so_x0y0s_L1_7__o,
        _i_sw_so_x0y0s_L1_6__o,
        _i_sw_so_x0y0s_L1_5__o,
        _i_sw_so_x0y0s_L1_4__o,
        _i_sw_so_x0y0s_L1_3__o,
        _i_sw_so_x0y0s_L1_2__o,
        _i_sw_so_x0y0s_L1_1__o,
        _i_sw_so_x0y0s_L1_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_nw_E_ex_e (
    input wire [11:0] bi_u1y0n_L1
    , output wire [11:0] so_x0y0e_L1
    , input wire [11:0] bi_u1y1s_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_so_x0y0e_L1_0__o;
    wire [0:0] _i_sw_so_x0y0e_L1_1__o;
    wire [0:0] _i_sw_so_x0y0e_L1_2__o;
    wire [0:0] _i_sw_so_x0y0e_L1_3__o;
    wire [0:0] _i_sw_so_x0y0e_L1_4__o;
    wire [0:0] _i_sw_so_x0y0e_L1_5__o;
    wire [0:0] _i_sw_so_x0y0e_L1_6__o;
    wire [0:0] _i_sw_so_x0y0e_L1_7__o;
    wire [0:0] _i_sw_so_x0y0e_L1_8__o;
    wire [0:0] _i_sw_so_x0y0e_L1_9__o;
    wire [0:0] _i_sw_so_x0y0e_L1_10__o;
    wire [0:0] _i_sw_so_x0y0e_L1_11__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_0__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_4__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_4__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_5__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_5__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_6__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_7__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_8__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_9__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_9__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_10__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_10__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_11__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_11__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw1 i_sw_so_x0y0e_L1_0 (
        .i(bi_u1y1s_L1[1])
        ,.o(_i_sw_so_x0y0e_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_0__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_1 (
        .i({bi_u1y1s_L1[2],
            bi_u1y0n_L1[3]})
        ,.o(_i_sw_so_x0y0e_L1_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_1__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_2 (
        .i({bi_u1y1s_L1[3],
            bi_u1y0n_L1[4]})
        ,.o(_i_sw_so_x0y0e_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_2__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_3 (
        .i({bi_u1y1s_L1[4],
            bi_u1y0n_L1[5]})
        ,.o(_i_sw_so_x0y0e_L1_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_3__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_4 (
        .i({bi_u1y1s_L1[5],
            bi_u1y0n_L1[6]})
        ,.o(_i_sw_so_x0y0e_L1_4__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_4__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_5 (
        .i({bi_u1y1s_L1[6],
            bi_u1y0n_L1[7]})
        ,.o(_i_sw_so_x0y0e_L1_5__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_5__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_6 (
        .i({bi_u1y1s_L1[7],
            bi_u1y0n_L1[8]})
        ,.o(_i_sw_so_x0y0e_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_6__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_7 (
        .i({bi_u1y1s_L1[8],
            bi_u1y0n_L1[9]})
        ,.o(_i_sw_so_x0y0e_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_7__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_8 (
        .i({bi_u1y1s_L1[9],
            bi_u1y0n_L1[10]})
        ,.o(_i_sw_so_x0y0e_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_8__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_9 (
        .i({bi_u1y1s_L1[10],
            bi_u1y0n_L1[11]})
        ,.o(_i_sw_so_x0y0e_L1_9__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_9__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_10 (
        .i({bi_u1y1s_L1[11],
            bi_u1y0n_L1[0]})
        ,.o(_i_sw_so_x0y0e_L1_10__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_10__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_11 (
        .i({bi_u1y1s_L1[0],
            bi_u1y0n_L1[1]})
        ,.o(_i_sw_so_x0y0e_L1_11__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_11__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0y0e_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_3__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_4 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_4__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_4__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_5 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_4__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_5__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_5__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_5__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_6__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_7__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_8__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_9 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_9__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_9__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_10 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_9__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_10__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_10__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_11 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_10__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_11__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_11__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_11__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign so_x0y0e_L1 = {_i_sw_so_x0y0e_L1_11__o,
        _i_sw_so_x0y0e_L1_10__o,
        _i_sw_so_x0y0e_L1_9__o,
        _i_sw_so_x0y0e_L1_8__o,
        _i_sw_so_x0y0e_L1_7__o,
        _i_sw_so_x0y0e_L1_6__o,
        _i_sw_so_x0y0e_L1_5__o,
        _i_sw_so_x0y0e_L1_4__o,
        _i_sw_so_x0y0e_L1_3__o,
        _i_sw_so_x0y0e_L1_2__o,
        _i_sw_so_x0y0e_L1_1__o,
        _i_sw_so_x0y0e_L1_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_se_W_ex_n (
    input wire [11:0] bi_x0y0s_L1
    , output wire [11:0] so_x0v1w_L1
    , input wire [11:0] bi_x1v1w_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_so_x0v1w_L1_0__o;
    wire [0:0] _i_sw_so_x0v1w_L1_1__o;
    wire [0:0] _i_sw_so_x0v1w_L1_2__o;
    wire [0:0] _i_sw_so_x0v1w_L1_3__o;
    wire [0:0] _i_sw_so_x0v1w_L1_4__o;
    wire [0:0] _i_sw_so_x0v1w_L1_5__o;
    wire [0:0] _i_sw_so_x0v1w_L1_6__o;
    wire [0:0] _i_sw_so_x0v1w_L1_7__o;
    wire [0:0] _i_sw_so_x0v1w_L1_8__o;
    wire [0:0] _i_sw_so_x0v1w_L1_9__o;
    wire [0:0] _i_sw_so_x0v1w_L1_10__o;
    wire [0:0] _i_sw_so_x0v1w_L1_11__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_4__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_4__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_5__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_5__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_6__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_7__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_8__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_9__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_9__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_10__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_10__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_11__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_11__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw2 i_sw_so_x0v1w_L1_0 (
        .i({bi_x1v1w_L1[0],
            bi_x0y0s_L1[11]})
        ,.o(_i_sw_so_x0v1w_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_0__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_1 (
        .i({bi_x1v1w_L1[1],
            bi_x0y0s_L1[0]})
        ,.o(_i_sw_so_x0v1w_L1_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_1__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_2 (
        .i({bi_x1v1w_L1[2],
            bi_x0y0s_L1[1]})
        ,.o(_i_sw_so_x0v1w_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_2__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_3 (
        .i({bi_x1v1w_L1[3],
            bi_x0y0s_L1[2]})
        ,.o(_i_sw_so_x0v1w_L1_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_3__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_4 (
        .i({bi_x1v1w_L1[4],
            bi_x0y0s_L1[3]})
        ,.o(_i_sw_so_x0v1w_L1_4__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_4__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_5 (
        .i({bi_x1v1w_L1[5],
            bi_x0y0s_L1[4]})
        ,.o(_i_sw_so_x0v1w_L1_5__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_5__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_6 (
        .i({bi_x1v1w_L1[6],
            bi_x0y0s_L1[5]})
        ,.o(_i_sw_so_x0v1w_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_6__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_7 (
        .i({bi_x1v1w_L1[7],
            bi_x0y0s_L1[6]})
        ,.o(_i_sw_so_x0v1w_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_7__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_8 (
        .i({bi_x1v1w_L1[8],
            bi_x0y0s_L1[7]})
        ,.o(_i_sw_so_x0v1w_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_8__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_9 (
        .i({bi_x1v1w_L1[9],
            bi_x0y0s_L1[8]})
        ,.o(_i_sw_so_x0v1w_L1_9__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_9__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_10 (
        .i({bi_x1v1w_L1[10],
            bi_x0y0s_L1[9]})
        ,.o(_i_sw_so_x0v1w_L1_10__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_10__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_11 (
        .i({bi_x1v1w_L1[11],
            bi_x0y0s_L1[10]})
        ,.o(_i_sw_so_x0v1w_L1_11__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_11__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_3__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_4 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_4__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_4__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_5 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_4__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_5__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_5__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_5__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_6__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_7__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_8__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_9 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_9__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_9__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_10 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_9__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_10__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_10__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_11 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_10__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_11__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_11__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_11__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign so_x0v1w_L1 = {_i_sw_so_x0v1w_L1_11__o,
        _i_sw_so_x0v1w_L1_10__o,
        _i_sw_so_x0v1w_L1_9__o,
        _i_sw_so_x0v1w_L1_8__o,
        _i_sw_so_x0v1w_L1_7__o,
        _i_sw_so_x0v1w_L1_6__o,
        _i_sw_so_x0v1w_L1_5__o,
        _i_sw_so_x0v1w_L1_4__o,
        _i_sw_so_x0v1w_L1_3__o,
        _i_sw_so_x0v1w_L1_2__o,
        _i_sw_so_x0v1w_L1_1__o,
        _i_sw_so_x0v1w_L1_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_sw_N_ex_ne (
    input wire [11:0] bi_x0v1w_L1
    , output wire [11:0] so_u1y0n_L1
    , input wire [11:0] cu_u1y0n_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_so_u1y0n_L1_0__o;
    wire [0:0] _i_sw_so_u1y0n_L1_1__o;
    wire [0:0] _i_sw_so_u1y0n_L1_2__o;
    wire [0:0] _i_sw_so_u1y0n_L1_3__o;
    wire [0:0] _i_sw_so_u1y0n_L1_4__o;
    wire [0:0] _i_sw_so_u1y0n_L1_5__o;
    wire [0:0] _i_sw_so_u1y0n_L1_6__o;
    wire [0:0] _i_sw_so_u1y0n_L1_7__o;
    wire [0:0] _i_sw_so_u1y0n_L1_8__o;
    wire [0:0] _i_sw_so_u1y0n_L1_9__o;
    wire [0:0] _i_sw_so_u1y0n_L1_10__o;
    wire [0:0] _i_sw_so_u1y0n_L1_11__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_4__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_4__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_5__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_5__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_6__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_7__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_8__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_9__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_9__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_10__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_10__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_11__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_11__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw2 i_sw_so_u1y0n_L1_0 (
        .i({cu_u1y0n_L1[0],
            bi_x0v1w_L1[11]})
        ,.o(_i_sw_so_u1y0n_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_0__prog_data)
        );
    sw2 i_sw_so_u1y0n_L1_1 (
        .i({cu_u1y0n_L1[1],
            bi_x0v1w_L1[0]})
        ,.o(_i_sw_so_u1y0n_L1_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_1__prog_data)
        );
    sw2 i_sw_so_u1y0n_L1_2 (
        .i({cu_u1y0n_L1[2],
            bi_x0v1w_L1[1]})
        ,.o(_i_sw_so_u1y0n_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_2__prog_data)
        );
    sw2 i_sw_so_u1y0n_L1_3 (
        .i({cu_u1y0n_L1[3],
            bi_x0v1w_L1[2]})
        ,.o(_i_sw_so_u1y0n_L1_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_3__prog_data)
        );
    sw2 i_sw_so_u1y0n_L1_4 (
        .i({cu_u1y0n_L1[4],
            bi_x0v1w_L1[3]})
        ,.o(_i_sw_so_u1y0n_L1_4__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_4__prog_data)
        );
    sw2 i_sw_so_u1y0n_L1_5 (
        .i({cu_u1y0n_L1[5],
            bi_x0v1w_L1[4]})
        ,.o(_i_sw_so_u1y0n_L1_5__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_5__prog_data)
        );
    sw2 i_sw_so_u1y0n_L1_6 (
        .i({cu_u1y0n_L1[6],
            bi_x0v1w_L1[5]})
        ,.o(_i_sw_so_u1y0n_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_6__prog_data)
        );
    sw2 i_sw_so_u1y0n_L1_7 (
        .i({cu_u1y0n_L1[7],
            bi_x0v1w_L1[6]})
        ,.o(_i_sw_so_u1y0n_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_7__prog_data)
        );
    sw2 i_sw_so_u1y0n_L1_8 (
        .i({cu_u1y0n_L1[8],
            bi_x0v1w_L1[7]})
        ,.o(_i_sw_so_u1y0n_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_8__prog_data)
        );
    sw2 i_sw_so_u1y0n_L1_9 (
        .i({cu_u1y0n_L1[9],
            bi_x0v1w_L1[8]})
        ,.o(_i_sw_so_u1y0n_L1_9__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_9__prog_data)
        );
    sw2 i_sw_so_u1y0n_L1_10 (
        .i({cu_u1y0n_L1[10],
            bi_x0v1w_L1[9]})
        ,.o(_i_sw_so_u1y0n_L1_10__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_10__prog_data)
        );
    sw2 i_sw_so_u1y0n_L1_11 (
        .i({cu_u1y0n_L1[11],
            bi_x0v1w_L1[10]})
        ,.o(_i_sw_so_u1y0n_L1_11__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_11__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_3__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_4 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_4__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_4__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_5 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_4__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_5__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_5__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_5__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_6__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_7__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_8__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_9 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_9__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_9__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_10 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_9__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_10__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_10__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_11 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_10__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_11__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_11__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_11__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign so_u1y0n_L1 = {_i_sw_so_u1y0n_L1_11__o,
        _i_sw_so_u1y0n_L1_10__o,
        _i_sw_so_u1y0n_L1_9__o,
        _i_sw_so_u1y0n_L1_8__o,
        _i_sw_so_u1y0n_L1_7__o,
        _i_sw_so_u1y0n_L1_6__o,
        _i_sw_so_u1y0n_L1_5__o,
        _i_sw_so_u1y0n_L1_4__o,
        _i_sw_so_u1y0n_L1_3__o,
        _i_sw_so_u1y0n_L1_2__o,
        _i_sw_so_u1y0n_L1_1__o,
        _i_sw_so_u1y0n_L1_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_se_W (
    input wire [11:0] bi_x0v1n_L1
    , output wire [11:0] so_x0v1w_L1
    , input wire [11:0] bi_x0y0s_L1
    , input wire [11:0] bi_x1v1w_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_so_x0v1w_L1_0__o;
    wire [0:0] _i_sw_so_x0v1w_L1_1__o;
    wire [0:0] _i_sw_so_x0v1w_L1_2__o;
    wire [0:0] _i_sw_so_x0v1w_L1_3__o;
    wire [0:0] _i_sw_so_x0v1w_L1_4__o;
    wire [0:0] _i_sw_so_x0v1w_L1_5__o;
    wire [0:0] _i_sw_so_x0v1w_L1_6__o;
    wire [0:0] _i_sw_so_x0v1w_L1_7__o;
    wire [0:0] _i_sw_so_x0v1w_L1_8__o;
    wire [0:0] _i_sw_so_x0v1w_L1_9__o;
    wire [0:0] _i_sw_so_x0v1w_L1_10__o;
    wire [0:0] _i_sw_so_x0v1w_L1_11__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_4__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_4__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_5__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_5__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_6__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_7__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_8__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_9__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_9__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_10__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_10__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_11__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_11__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw3 i_sw_so_x0v1w_L1_0 (
        .i({bi_x1v1w_L1[0],
            bi_x0y0s_L1[11],
            bi_x0v1n_L1[1]})
        ,.o(_i_sw_so_x0v1w_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_0__prog_data)
        );
    sw3 i_sw_so_x0v1w_L1_1 (
        .i({bi_x1v1w_L1[1],
            bi_x0y0s_L1[0],
            bi_x0v1n_L1[2]})
        ,.o(_i_sw_so_x0v1w_L1_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_1__prog_data)
        );
    sw3 i_sw_so_x0v1w_L1_2 (
        .i({bi_x1v1w_L1[2],
            bi_x0y0s_L1[1],
            bi_x0v1n_L1[3]})
        ,.o(_i_sw_so_x0v1w_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_2__prog_data)
        );
    sw3 i_sw_so_x0v1w_L1_3 (
        .i({bi_x1v1w_L1[3],
            bi_x0y0s_L1[2],
            bi_x0v1n_L1[4]})
        ,.o(_i_sw_so_x0v1w_L1_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_3__prog_data)
        );
    sw3 i_sw_so_x0v1w_L1_4 (
        .i({bi_x1v1w_L1[4],
            bi_x0y0s_L1[3],
            bi_x0v1n_L1[5]})
        ,.o(_i_sw_so_x0v1w_L1_4__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_4__prog_data)
        );
    sw3 i_sw_so_x0v1w_L1_5 (
        .i({bi_x1v1w_L1[5],
            bi_x0y0s_L1[4],
            bi_x0v1n_L1[6]})
        ,.o(_i_sw_so_x0v1w_L1_5__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_5__prog_data)
        );
    sw3 i_sw_so_x0v1w_L1_6 (
        .i({bi_x1v1w_L1[6],
            bi_x0y0s_L1[5],
            bi_x0v1n_L1[7]})
        ,.o(_i_sw_so_x0v1w_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_6__prog_data)
        );
    sw3 i_sw_so_x0v1w_L1_7 (
        .i({bi_x1v1w_L1[7],
            bi_x0y0s_L1[6],
            bi_x0v1n_L1[8]})
        ,.o(_i_sw_so_x0v1w_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_7__prog_data)
        );
    sw3 i_sw_so_x0v1w_L1_8 (
        .i({bi_x1v1w_L1[8],
            bi_x0y0s_L1[7],
            bi_x0v1n_L1[9]})
        ,.o(_i_sw_so_x0v1w_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_8__prog_data)
        );
    sw3 i_sw_so_x0v1w_L1_9 (
        .i({bi_x1v1w_L1[9],
            bi_x0y0s_L1[8],
            bi_x0v1n_L1[10]})
        ,.o(_i_sw_so_x0v1w_L1_9__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_9__prog_data)
        );
    sw3 i_sw_so_x0v1w_L1_10 (
        .i({bi_x1v1w_L1[10],
            bi_x0y0s_L1[9],
            bi_x0v1n_L1[11]})
        ,.o(_i_sw_so_x0v1w_L1_10__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_10__prog_data)
        );
    sw3 i_sw_so_x0v1w_L1_11 (
        .i({bi_x1v1w_L1[11],
            bi_x0y0s_L1[10],
            bi_x0v1n_L1[0]})
        ,.o(_i_sw_so_x0v1w_L1_11__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_11__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_3__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_4 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_4__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_4__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_5 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_4__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_5__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_5__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_5__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_6__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_7__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_8__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_9 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_9__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_9__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_10 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_9__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_10__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_10__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_11 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_10__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_11__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_11__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_11__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign so_x0v1w_L1 = {_i_sw_so_x0v1w_L1_11__o,
        _i_sw_so_x0v1w_L1_10__o,
        _i_sw_so_x0v1w_L1_9__o,
        _i_sw_so_x0v1w_L1_8__o,
        _i_sw_so_x0v1w_L1_7__o,
        _i_sw_so_x0v1w_L1_6__o,
        _i_sw_so_x0v1w_L1_5__o,
        _i_sw_so_x0v1w_L1_4__o,
        _i_sw_so_x0v1w_L1_3__o,
        _i_sw_so_x0v1w_L1_2__o,
        _i_sw_so_x0v1w_L1_1__o,
        _i_sw_so_x0v1w_L1_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_sw_N_ex_e (
    input wire [11:0] bi_u1v1n_L1
    , output wire [11:0] so_u1y0n_L1
    , input wire [11:0] bi_x0v1w_L1
    , input wire [11:0] cu_u1y0n_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_so_u1y0n_L1_0__o;
    wire [0:0] _i_sw_so_u1y0n_L1_1__o;
    wire [0:0] _i_sw_so_u1y0n_L1_2__o;
    wire [0:0] _i_sw_so_u1y0n_L1_3__o;
    wire [0:0] _i_sw_so_u1y0n_L1_4__o;
    wire [0:0] _i_sw_so_u1y0n_L1_5__o;
    wire [0:0] _i_sw_so_u1y0n_L1_6__o;
    wire [0:0] _i_sw_so_u1y0n_L1_7__o;
    wire [0:0] _i_sw_so_u1y0n_L1_8__o;
    wire [0:0] _i_sw_so_u1y0n_L1_9__o;
    wire [0:0] _i_sw_so_u1y0n_L1_10__o;
    wire [0:0] _i_sw_so_u1y0n_L1_11__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_4__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_4__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_5__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_5__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_6__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_7__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_8__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_9__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_9__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_10__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_10__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_11__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_11__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw3 i_sw_so_u1y0n_L1_0 (
        .i({cu_u1y0n_L1[0],
            bi_x0v1w_L1[11],
            bi_u1v1n_L1[0]})
        ,.o(_i_sw_so_u1y0n_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_0__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_1 (
        .i({cu_u1y0n_L1[1],
            bi_x0v1w_L1[0],
            bi_u1v1n_L1[1]})
        ,.o(_i_sw_so_u1y0n_L1_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_1__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_2 (
        .i({cu_u1y0n_L1[2],
            bi_x0v1w_L1[1],
            bi_u1v1n_L1[2]})
        ,.o(_i_sw_so_u1y0n_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_2__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_3 (
        .i({cu_u1y0n_L1[3],
            bi_x0v1w_L1[2],
            bi_u1v1n_L1[3]})
        ,.o(_i_sw_so_u1y0n_L1_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_3__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_4 (
        .i({cu_u1y0n_L1[4],
            bi_x0v1w_L1[3],
            bi_u1v1n_L1[4]})
        ,.o(_i_sw_so_u1y0n_L1_4__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_4__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_5 (
        .i({cu_u1y0n_L1[5],
            bi_x0v1w_L1[4],
            bi_u1v1n_L1[5]})
        ,.o(_i_sw_so_u1y0n_L1_5__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_5__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_6 (
        .i({cu_u1y0n_L1[6],
            bi_x0v1w_L1[5],
            bi_u1v1n_L1[6]})
        ,.o(_i_sw_so_u1y0n_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_6__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_7 (
        .i({cu_u1y0n_L1[7],
            bi_x0v1w_L1[6],
            bi_u1v1n_L1[7]})
        ,.o(_i_sw_so_u1y0n_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_7__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_8 (
        .i({cu_u1y0n_L1[8],
            bi_x0v1w_L1[7],
            bi_u1v1n_L1[8]})
        ,.o(_i_sw_so_u1y0n_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_8__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_9 (
        .i({cu_u1y0n_L1[9],
            bi_x0v1w_L1[8],
            bi_u1v1n_L1[9]})
        ,.o(_i_sw_so_u1y0n_L1_9__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_9__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_10 (
        .i({cu_u1y0n_L1[10],
            bi_x0v1w_L1[9],
            bi_u1v1n_L1[10]})
        ,.o(_i_sw_so_u1y0n_L1_10__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_10__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_11 (
        .i({cu_u1y0n_L1[11],
            bi_x0v1w_L1[10],
            bi_u1v1n_L1[11]})
        ,.o(_i_sw_so_u1y0n_L1_11__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_11__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_3__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_4 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_4__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_4__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_5 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_4__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_5__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_5__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_5__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_6__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_7__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_8__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_9 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_9__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_9__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_10 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_9__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_10__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_10__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_11 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_10__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_11__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_11__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_11__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign so_u1y0n_L1 = {_i_sw_so_u1y0n_L1_11__o,
        _i_sw_so_u1y0n_L1_10__o,
        _i_sw_so_u1y0n_L1_9__o,
        _i_sw_so_u1y0n_L1_8__o,
        _i_sw_so_u1y0n_L1_7__o,
        _i_sw_so_u1y0n_L1_6__o,
        _i_sw_so_u1y0n_L1_5__o,
        _i_sw_so_u1y0n_L1_4__o,
        _i_sw_so_u1y0n_L1_3__o,
        _i_sw_so_u1y0n_L1_2__o,
        _i_sw_so_u1y0n_L1_1__o,
        _i_sw_so_u1y0n_L1_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_ne_S_ex_s (
    input wire [11:0] bi_x0y0e_L1
    , output wire [11:0] so_x0y0s_L1
    , input wire [11:0] bi_x1y0w_L1
    , input wire [11:0] cu_x0y0s_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_so_x0y0s_L1_0__o;
    wire [0:0] _i_sw_so_x0y0s_L1_1__o;
    wire [0:0] _i_sw_so_x0y0s_L1_2__o;
    wire [0:0] _i_sw_so_x0y0s_L1_3__o;
    wire [0:0] _i_sw_so_x0y0s_L1_4__o;
    wire [0:0] _i_sw_so_x0y0s_L1_5__o;
    wire [0:0] _i_sw_so_x0y0s_L1_6__o;
    wire [0:0] _i_sw_so_x0y0s_L1_7__o;
    wire [0:0] _i_sw_so_x0y0s_L1_8__o;
    wire [0:0] _i_sw_so_x0y0s_L1_9__o;
    wire [0:0] _i_sw_so_x0y0s_L1_10__o;
    wire [0:0] _i_sw_so_x0y0s_L1_11__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_4__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_4__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_5__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_5__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_6__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_7__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_8__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_9__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_9__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_10__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_10__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_11__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_11__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw3 i_sw_so_x0y0s_L1_0 (
        .i({cu_x0y0s_L1[0],
            bi_x1y0w_L1[0],
            bi_x0y0e_L1[11]})
        ,.o(_i_sw_so_x0y0s_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_0__prog_data)
        );
    sw2 i_sw_so_x0y0s_L1_1 (
        .i({cu_x0y0s_L1[1],
            bi_x0y0e_L1[0]})
        ,.o(_i_sw_so_x0y0s_L1_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_1__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_2 (
        .i({cu_x0y0s_L1[2],
            bi_x1y0w_L1[2],
            bi_x0y0e_L1[1]})
        ,.o(_i_sw_so_x0y0s_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_2__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_3 (
        .i({cu_x0y0s_L1[3],
            bi_x1y0w_L1[3],
            bi_x0y0e_L1[2]})
        ,.o(_i_sw_so_x0y0s_L1_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_3__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_4 (
        .i({cu_x0y0s_L1[4],
            bi_x1y0w_L1[4],
            bi_x0y0e_L1[3]})
        ,.o(_i_sw_so_x0y0s_L1_4__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_4__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_5 (
        .i({cu_x0y0s_L1[5],
            bi_x1y0w_L1[5],
            bi_x0y0e_L1[4]})
        ,.o(_i_sw_so_x0y0s_L1_5__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_5__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_6 (
        .i({cu_x0y0s_L1[6],
            bi_x1y0w_L1[6],
            bi_x0y0e_L1[5]})
        ,.o(_i_sw_so_x0y0s_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_6__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_7 (
        .i({cu_x0y0s_L1[7],
            bi_x1y0w_L1[7],
            bi_x0y0e_L1[6]})
        ,.o(_i_sw_so_x0y0s_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_7__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_8 (
        .i({cu_x0y0s_L1[8],
            bi_x1y0w_L1[8],
            bi_x0y0e_L1[7]})
        ,.o(_i_sw_so_x0y0s_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_8__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_9 (
        .i({cu_x0y0s_L1[9],
            bi_x1y0w_L1[9],
            bi_x0y0e_L1[8]})
        ,.o(_i_sw_so_x0y0s_L1_9__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_9__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_10 (
        .i({cu_x0y0s_L1[10],
            bi_x1y0w_L1[10],
            bi_x0y0e_L1[9]})
        ,.o(_i_sw_so_x0y0s_L1_10__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_10__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_11 (
        .i({cu_x0y0s_L1[11],
            bi_x1y0w_L1[11],
            bi_x0y0e_L1[10]})
        ,.o(_i_sw_so_x0y0s_L1_11__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_11__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_3__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_4 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_4__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_4__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_5 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_4__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_5__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_5__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_5__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_6__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_7__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_8__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_9 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_9__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_9__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_10 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_9__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_10__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_10__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_11 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_10__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_11__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_11__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_11__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign so_x0y0s_L1 = {_i_sw_so_x0y0s_L1_11__o,
        _i_sw_so_x0y0s_L1_10__o,
        _i_sw_so_x0y0s_L1_9__o,
        _i_sw_so_x0y0s_L1_8__o,
        _i_sw_so_x0y0s_L1_7__o,
        _i_sw_so_x0y0s_L1_6__o,
        _i_sw_so_x0y0s_L1_5__o,
        _i_sw_so_x0y0s_L1_4__o,
        _i_sw_so_x0y0s_L1_3__o,
        _i_sw_so_x0y0s_L1_2__o,
        _i_sw_so_x0y0s_L1_1__o,
        _i_sw_so_x0y0s_L1_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_nw_E_ex_es (
    input wire [11:0] bi_u1y0n_L1
    , output wire [11:0] so_x0y0e_L1
    , input wire [11:0] cu_x0y0e_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_so_x0y0e_L1_0__o;
    wire [0:0] _i_sw_so_x0y0e_L1_1__o;
    wire [0:0] _i_sw_so_x0y0e_L1_2__o;
    wire [0:0] _i_sw_so_x0y0e_L1_3__o;
    wire [0:0] _i_sw_so_x0y0e_L1_4__o;
    wire [0:0] _i_sw_so_x0y0e_L1_5__o;
    wire [0:0] _i_sw_so_x0y0e_L1_6__o;
    wire [0:0] _i_sw_so_x0y0e_L1_7__o;
    wire [0:0] _i_sw_so_x0y0e_L1_8__o;
    wire [0:0] _i_sw_so_x0y0e_L1_9__o;
    wire [0:0] _i_sw_so_x0y0e_L1_10__o;
    wire [0:0] _i_sw_so_x0y0e_L1_11__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_0__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_4__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_4__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_5__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_5__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_6__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_7__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_8__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_9__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_9__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_10__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_10__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_11__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_11__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw1 i_sw_so_x0y0e_L1_0 (
        .i(cu_x0y0e_L1[0])
        ,.o(_i_sw_so_x0y0e_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_0__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_1 (
        .i({cu_x0y0e_L1[1],
            bi_u1y0n_L1[3]})
        ,.o(_i_sw_so_x0y0e_L1_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_1__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_2 (
        .i({cu_x0y0e_L1[2],
            bi_u1y0n_L1[4]})
        ,.o(_i_sw_so_x0y0e_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_2__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_3 (
        .i({cu_x0y0e_L1[3],
            bi_u1y0n_L1[5]})
        ,.o(_i_sw_so_x0y0e_L1_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_3__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_4 (
        .i({cu_x0y0e_L1[4],
            bi_u1y0n_L1[6]})
        ,.o(_i_sw_so_x0y0e_L1_4__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_4__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_5 (
        .i({cu_x0y0e_L1[5],
            bi_u1y0n_L1[7]})
        ,.o(_i_sw_so_x0y0e_L1_5__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_5__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_6 (
        .i({cu_x0y0e_L1[6],
            bi_u1y0n_L1[8]})
        ,.o(_i_sw_so_x0y0e_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_6__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_7 (
        .i({cu_x0y0e_L1[7],
            bi_u1y0n_L1[9]})
        ,.o(_i_sw_so_x0y0e_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_7__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_8 (
        .i({cu_x0y0e_L1[8],
            bi_u1y0n_L1[10]})
        ,.o(_i_sw_so_x0y0e_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_8__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_9 (
        .i({cu_x0y0e_L1[9],
            bi_u1y0n_L1[11]})
        ,.o(_i_sw_so_x0y0e_L1_9__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_9__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_10 (
        .i({cu_x0y0e_L1[10],
            bi_u1y0n_L1[0]})
        ,.o(_i_sw_so_x0y0e_L1_10__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_10__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_11 (
        .i({cu_x0y0e_L1[11],
            bi_u1y0n_L1[1]})
        ,.o(_i_sw_so_x0y0e_L1_11__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_11__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0y0e_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_3__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_4 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_4__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_4__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_5 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_4__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_5__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_5__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_5__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_6__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_7__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_8__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_9 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_9__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_9__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_10 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_9__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_10__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_10__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_11 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_10__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_11__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_11__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_11__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign so_x0y0e_L1 = {_i_sw_so_x0y0e_L1_11__o,
        _i_sw_so_x0y0e_L1_10__o,
        _i_sw_so_x0y0e_L1_9__o,
        _i_sw_so_x0y0e_L1_8__o,
        _i_sw_so_x0y0e_L1_7__o,
        _i_sw_so_x0y0e_L1_6__o,
        _i_sw_so_x0y0e_L1_5__o,
        _i_sw_so_x0y0e_L1_4__o,
        _i_sw_so_x0y0e_L1_3__o,
        _i_sw_so_x0y0e_L1_2__o,
        _i_sw_so_x0y0e_L1_1__o,
        _i_sw_so_x0y0e_L1_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module t_io_n (
    input wire [11:0] bi_x0v1e_L1
    , input wire [11:0] bi_x0v1w_L1
    , output wire [11:0] cu_x0v1e_L1
    , output wire [11:0] cu_x0v1w_L1
    , input wire [0:0] ipin_x0y0_0
    , output wire [0:0] opin_x0y0_0
    , output wire [0:0] oe_x0y0_0
    , input wire [0:0] ipin_x0y0_1
    , output wire [0:0] opin_x0y0_1
    , output wire [0:0] oe_x0y0_1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_blk_i0__inpad;
    wire [0:0] _i_blk_i0__opin;
    wire [0:0] _i_blk_i0__oe;
    wire [0:0] _i_blk_i0__prog_dout;
    wire [0:0] _i_blk_i0__prog_we_o;
    wire [0:0] _i_blk_i1__inpad;
    wire [0:0] _i_blk_i1__opin;
    wire [0:0] _i_blk_i1__oe;
    wire [0:0] _i_blk_i1__prog_dout;
    wire [0:0] _i_blk_i1__prog_we_o;
    wire [0:0] _i_cbox_s0__bp_x0y0i0_outpad;
    wire [11:0] _i_cbox_s0__cu_x0v1e_L1;
    wire [11:0] _i_cbox_s0__cu_x0v1w_L1;
    wire [0:0] _i_cbox_s0__bp_x0y0i1_outpad;
    wire [0:0] _i_cbox_s0__prog_dout;
    wire [0:0] _i_cbox_s0__prog_we_o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_buf_prog_rst_l1__Q;
    wire [0:0] _i_buf_prog_done_l1__Q;
        
    iob i_blk_i0 (
        .outpad(_i_cbox_s0__bp_x0y0i0_outpad)
        ,.inpad(_i_blk_i0__inpad)
        ,.ipin(ipin_x0y0_0)
        ,.opin(_i_blk_i0__opin)
        ,.oe(_i_blk_i0__oe)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_blk_i0__prog_dout)
        ,.prog_we_o(_i_blk_i0__prog_we_o)
        );
    iob i_blk_i1 (
        .outpad(_i_cbox_s0__bp_x0y0i1_outpad)
        ,.inpad(_i_blk_i1__inpad)
        ,.ipin(ipin_x0y0_1)
        ,.opin(_i_blk_i1__opin)
        ,.oe(_i_blk_i1__oe)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_blk_i0__prog_we_o)
        ,.prog_din(_i_blk_i0__prog_dout)
        ,.prog_dout(_i_blk_i1__prog_dout)
        ,.prog_we_o(_i_blk_i1__prog_we_o)
        );
    cbox_t_io_n_s0 i_cbox_s0 (
        .bp_x0y0i0_outpad(_i_cbox_s0__bp_x0y0i0_outpad)
        ,.bi_x0v1e_L1(bi_x0v1e_L1)
        ,.bi_x0v1w_L1(bi_x0v1w_L1)
        ,.bp_x0y0i0_inpad(_i_blk_i0__inpad)
        ,.cu_x0v1e_L1(_i_cbox_s0__cu_x0v1e_L1)
        ,.cu_x0v1w_L1(_i_cbox_s0__cu_x0v1w_L1)
        ,.bp_x0y0i1_outpad(_i_cbox_s0__bp_x0y0i1_outpad)
        ,.bp_x0y0i1_inpad(_i_blk_i1__inpad)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_blk_i1__prog_we_o)
        ,.prog_din(_i_blk_i1__prog_dout)
        ,.prog_dout(_i_cbox_s0__prog_dout)
        ,.prog_we_o(_i_cbox_s0__prog_we_o)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(_i_buf_prog_rst_l1__Q)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(_i_buf_prog_done_l1__Q)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    prga_simple_buf i_buf_prog_rst_l1 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l1__Q)
        );
    prga_simple_bufr i_buf_prog_done_l1 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l1__Q)
        );
        
    assign cu_x0v1e_L1 = _i_cbox_s0__cu_x0v1e_L1;
    assign cu_x0v1w_L1 = _i_cbox_s0__cu_x0v1w_L1;
    assign opin_x0y0_0 = _i_blk_i0__opin;
    assign oe_x0y0_0 = _i_blk_i0__oe;
    assign opin_x0y0_1 = _i_blk_i1__opin;
    assign oe_x0y0_1 = _i_blk_i1__oe;
    assign prog_dout = _i_cbox_s0__prog_dout;
    assign prog_we_o = _i_cbox_s0__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_se_W_ex_s (
    input wire [11:0] bi_x0v1n_L1
    , output wire [11:0] so_x0v1w_L1
    , input wire [11:0] bi_x1v1w_L1
    , input wire [11:0] cu_x0v1w_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_so_x0v1w_L1_0__o;
    wire [0:0] _i_sw_so_x0v1w_L1_1__o;
    wire [0:0] _i_sw_so_x0v1w_L1_2__o;
    wire [0:0] _i_sw_so_x0v1w_L1_3__o;
    wire [0:0] _i_sw_so_x0v1w_L1_4__o;
    wire [0:0] _i_sw_so_x0v1w_L1_5__o;
    wire [0:0] _i_sw_so_x0v1w_L1_6__o;
    wire [0:0] _i_sw_so_x0v1w_L1_7__o;
    wire [0:0] _i_sw_so_x0v1w_L1_8__o;
    wire [0:0] _i_sw_so_x0v1w_L1_9__o;
    wire [0:0] _i_sw_so_x0v1w_L1_10__o;
    wire [0:0] _i_sw_so_x0v1w_L1_11__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_4__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_4__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_5__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_5__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_6__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_7__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_8__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_9__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_9__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_10__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_10__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_11__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_11__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw3 i_sw_so_x0v1w_L1_0 (
        .i({cu_x0v1w_L1[0],
            bi_x1v1w_L1[0],
            bi_x0v1n_L1[1]})
        ,.o(_i_sw_so_x0v1w_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_0__prog_data)
        );
    sw3 i_sw_so_x0v1w_L1_1 (
        .i({cu_x0v1w_L1[1],
            bi_x1v1w_L1[1],
            bi_x0v1n_L1[2]})
        ,.o(_i_sw_so_x0v1w_L1_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_1__prog_data)
        );
    sw3 i_sw_so_x0v1w_L1_2 (
        .i({cu_x0v1w_L1[2],
            bi_x1v1w_L1[2],
            bi_x0v1n_L1[3]})
        ,.o(_i_sw_so_x0v1w_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_2__prog_data)
        );
    sw3 i_sw_so_x0v1w_L1_3 (
        .i({cu_x0v1w_L1[3],
            bi_x1v1w_L1[3],
            bi_x0v1n_L1[4]})
        ,.o(_i_sw_so_x0v1w_L1_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_3__prog_data)
        );
    sw3 i_sw_so_x0v1w_L1_4 (
        .i({cu_x0v1w_L1[4],
            bi_x1v1w_L1[4],
            bi_x0v1n_L1[5]})
        ,.o(_i_sw_so_x0v1w_L1_4__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_4__prog_data)
        );
    sw3 i_sw_so_x0v1w_L1_5 (
        .i({cu_x0v1w_L1[5],
            bi_x1v1w_L1[5],
            bi_x0v1n_L1[6]})
        ,.o(_i_sw_so_x0v1w_L1_5__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_5__prog_data)
        );
    sw3 i_sw_so_x0v1w_L1_6 (
        .i({cu_x0v1w_L1[6],
            bi_x1v1w_L1[6],
            bi_x0v1n_L1[7]})
        ,.o(_i_sw_so_x0v1w_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_6__prog_data)
        );
    sw3 i_sw_so_x0v1w_L1_7 (
        .i({cu_x0v1w_L1[7],
            bi_x1v1w_L1[7],
            bi_x0v1n_L1[8]})
        ,.o(_i_sw_so_x0v1w_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_7__prog_data)
        );
    sw3 i_sw_so_x0v1w_L1_8 (
        .i({cu_x0v1w_L1[8],
            bi_x1v1w_L1[8],
            bi_x0v1n_L1[9]})
        ,.o(_i_sw_so_x0v1w_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_8__prog_data)
        );
    sw3 i_sw_so_x0v1w_L1_9 (
        .i({cu_x0v1w_L1[9],
            bi_x1v1w_L1[9],
            bi_x0v1n_L1[10]})
        ,.o(_i_sw_so_x0v1w_L1_9__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_9__prog_data)
        );
    sw3 i_sw_so_x0v1w_L1_10 (
        .i({cu_x0v1w_L1[10],
            bi_x1v1w_L1[10],
            bi_x0v1n_L1[11]})
        ,.o(_i_sw_so_x0v1w_L1_10__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_10__prog_data)
        );
    sw3 i_sw_so_x0v1w_L1_11 (
        .i({cu_x0v1w_L1[11],
            bi_x1v1w_L1[11],
            bi_x0v1n_L1[0]})
        ,.o(_i_sw_so_x0v1w_L1_11__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_11__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_3__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_4 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_4__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_4__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_5 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_4__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_5__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_5__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_5__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_6__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_7__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_8__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_9 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_9__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_9__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_10 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_9__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_10__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_10__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_11 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_10__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_11__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_11__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_11__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign so_x0v1w_L1 = {_i_sw_so_x0v1w_L1_11__o,
        _i_sw_so_x0v1w_L1_10__o,
        _i_sw_so_x0v1w_L1_9__o,
        _i_sw_so_x0v1w_L1_8__o,
        _i_sw_so_x0v1w_L1_7__o,
        _i_sw_so_x0v1w_L1_6__o,
        _i_sw_so_x0v1w_L1_5__o,
        _i_sw_so_x0v1w_L1_4__o,
        _i_sw_so_x0v1w_L1_3__o,
        _i_sw_so_x0v1w_L1_2__o,
        _i_sw_so_x0v1w_L1_1__o,
        _i_sw_so_x0v1w_L1_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_sw_s_ex_es (
    input wire [11:0] bi_x0v1w_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    );
    
        
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
        
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
        

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_nw_E_ex_n (
    input wire [11:0] bi_u1y0e_L1
    , output wire [11:0] so_x0y0e_L1
    , input wire [11:0] bi_u1y1s_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_so_x0y0e_L1_0__o;
    wire [0:0] _i_sw_so_x0y0e_L1_1__o;
    wire [0:0] _i_sw_so_x0y0e_L1_2__o;
    wire [0:0] _i_sw_so_x0y0e_L1_3__o;
    wire [0:0] _i_sw_so_x0y0e_L1_4__o;
    wire [0:0] _i_sw_so_x0y0e_L1_5__o;
    wire [0:0] _i_sw_so_x0y0e_L1_6__o;
    wire [0:0] _i_sw_so_x0y0e_L1_7__o;
    wire [0:0] _i_sw_so_x0y0e_L1_8__o;
    wire [0:0] _i_sw_so_x0y0e_L1_9__o;
    wire [0:0] _i_sw_so_x0y0e_L1_10__o;
    wire [0:0] _i_sw_so_x0y0e_L1_11__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_4__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_4__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_5__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_5__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_6__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_7__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_8__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_9__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_9__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_10__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_10__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_11__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_11__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw2 i_sw_so_x0y0e_L1_0 (
        .i({bi_u1y1s_L1[1],
            bi_u1y0e_L1[0]})
        ,.o(_i_sw_so_x0y0e_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_0__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_1 (
        .i({bi_u1y1s_L1[2],
            bi_u1y0e_L1[1]})
        ,.o(_i_sw_so_x0y0e_L1_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_1__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_2 (
        .i({bi_u1y1s_L1[3],
            bi_u1y0e_L1[2]})
        ,.o(_i_sw_so_x0y0e_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_2__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_3 (
        .i({bi_u1y1s_L1[4],
            bi_u1y0e_L1[3]})
        ,.o(_i_sw_so_x0y0e_L1_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_3__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_4 (
        .i({bi_u1y1s_L1[5],
            bi_u1y0e_L1[4]})
        ,.o(_i_sw_so_x0y0e_L1_4__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_4__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_5 (
        .i({bi_u1y1s_L1[6],
            bi_u1y0e_L1[5]})
        ,.o(_i_sw_so_x0y0e_L1_5__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_5__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_6 (
        .i({bi_u1y1s_L1[7],
            bi_u1y0e_L1[6]})
        ,.o(_i_sw_so_x0y0e_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_6__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_7 (
        .i({bi_u1y1s_L1[8],
            bi_u1y0e_L1[7]})
        ,.o(_i_sw_so_x0y0e_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_7__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_8 (
        .i({bi_u1y1s_L1[9],
            bi_u1y0e_L1[8]})
        ,.o(_i_sw_so_x0y0e_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_8__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_9 (
        .i({bi_u1y1s_L1[10],
            bi_u1y0e_L1[9]})
        ,.o(_i_sw_so_x0y0e_L1_9__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_9__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_10 (
        .i({bi_u1y1s_L1[11],
            bi_u1y0e_L1[10]})
        ,.o(_i_sw_so_x0y0e_L1_10__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_10__prog_data)
        );
    sw2 i_sw_so_x0y0e_L1_11 (
        .i({bi_u1y1s_L1[0],
            bi_u1y0e_L1[11]})
        ,.o(_i_sw_so_x0y0e_L1_11__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_11__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_3__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_4 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_4__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_4__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_5 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_4__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_5__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_5__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_5__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_6__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_7__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_8__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_9 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_9__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_9__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_10 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_9__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_10__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_10__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_11 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_10__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_11__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_11__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_11__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign so_x0y0e_L1 = {_i_sw_so_x0y0e_L1_11__o,
        _i_sw_so_x0y0e_L1_10__o,
        _i_sw_so_x0y0e_L1_9__o,
        _i_sw_so_x0y0e_L1_8__o,
        _i_sw_so_x0y0e_L1_7__o,
        _i_sw_so_x0y0e_L1_6__o,
        _i_sw_so_x0y0e_L1_5__o,
        _i_sw_so_x0y0e_L1_4__o,
        _i_sw_so_x0y0e_L1_3__o,
        _i_sw_so_x0y0e_L1_2__o,
        _i_sw_so_x0y0e_L1_1__o,
        _i_sw_so_x0y0e_L1_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_nw_E (
    input wire [11:0] bi_u1y0n_L1
    , output wire [11:0] so_x0y0e_L1
    , input wire [11:0] bi_u1y0e_L1
    , input wire [11:0] bi_u1y1s_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_so_x0y0e_L1_0__o;
    wire [0:0] _i_sw_so_x0y0e_L1_1__o;
    wire [0:0] _i_sw_so_x0y0e_L1_2__o;
    wire [0:0] _i_sw_so_x0y0e_L1_3__o;
    wire [0:0] _i_sw_so_x0y0e_L1_4__o;
    wire [0:0] _i_sw_so_x0y0e_L1_5__o;
    wire [0:0] _i_sw_so_x0y0e_L1_6__o;
    wire [0:0] _i_sw_so_x0y0e_L1_7__o;
    wire [0:0] _i_sw_so_x0y0e_L1_8__o;
    wire [0:0] _i_sw_so_x0y0e_L1_9__o;
    wire [0:0] _i_sw_so_x0y0e_L1_10__o;
    wire [0:0] _i_sw_so_x0y0e_L1_11__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_4__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_4__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_5__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_5__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_6__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_7__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_8__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_9__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_9__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_10__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_10__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_11__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_11__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw2 i_sw_so_x0y0e_L1_0 (
        .i({bi_u1y1s_L1[1],
            bi_u1y0e_L1[0]})
        ,.o(_i_sw_so_x0y0e_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_0__prog_data)
        );
    sw3 i_sw_so_x0y0e_L1_1 (
        .i({bi_u1y1s_L1[2],
            bi_u1y0e_L1[1],
            bi_u1y0n_L1[3]})
        ,.o(_i_sw_so_x0y0e_L1_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_1__prog_data)
        );
    sw3 i_sw_so_x0y0e_L1_2 (
        .i({bi_u1y1s_L1[3],
            bi_u1y0e_L1[2],
            bi_u1y0n_L1[4]})
        ,.o(_i_sw_so_x0y0e_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_2__prog_data)
        );
    sw3 i_sw_so_x0y0e_L1_3 (
        .i({bi_u1y1s_L1[4],
            bi_u1y0e_L1[3],
            bi_u1y0n_L1[5]})
        ,.o(_i_sw_so_x0y0e_L1_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_3__prog_data)
        );
    sw3 i_sw_so_x0y0e_L1_4 (
        .i({bi_u1y1s_L1[5],
            bi_u1y0e_L1[4],
            bi_u1y0n_L1[6]})
        ,.o(_i_sw_so_x0y0e_L1_4__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_4__prog_data)
        );
    sw3 i_sw_so_x0y0e_L1_5 (
        .i({bi_u1y1s_L1[6],
            bi_u1y0e_L1[5],
            bi_u1y0n_L1[7]})
        ,.o(_i_sw_so_x0y0e_L1_5__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_5__prog_data)
        );
    sw3 i_sw_so_x0y0e_L1_6 (
        .i({bi_u1y1s_L1[7],
            bi_u1y0e_L1[6],
            bi_u1y0n_L1[8]})
        ,.o(_i_sw_so_x0y0e_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_6__prog_data)
        );
    sw3 i_sw_so_x0y0e_L1_7 (
        .i({bi_u1y1s_L1[8],
            bi_u1y0e_L1[7],
            bi_u1y0n_L1[9]})
        ,.o(_i_sw_so_x0y0e_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_7__prog_data)
        );
    sw3 i_sw_so_x0y0e_L1_8 (
        .i({bi_u1y1s_L1[9],
            bi_u1y0e_L1[8],
            bi_u1y0n_L1[10]})
        ,.o(_i_sw_so_x0y0e_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_8__prog_data)
        );
    sw3 i_sw_so_x0y0e_L1_9 (
        .i({bi_u1y1s_L1[10],
            bi_u1y0e_L1[9],
            bi_u1y0n_L1[11]})
        ,.o(_i_sw_so_x0y0e_L1_9__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_9__prog_data)
        );
    sw3 i_sw_so_x0y0e_L1_10 (
        .i({bi_u1y1s_L1[11],
            bi_u1y0e_L1[10],
            bi_u1y0n_L1[0]})
        ,.o(_i_sw_so_x0y0e_L1_10__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_10__prog_data)
        );
    sw3 i_sw_so_x0y0e_L1_11 (
        .i({bi_u1y1s_L1[0],
            bi_u1y0e_L1[11],
            bi_u1y0n_L1[1]})
        ,.o(_i_sw_so_x0y0e_L1_11__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_11__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_3__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_4 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_4__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_4__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_5 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_4__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_5__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_5__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_5__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_6__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_7__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_8__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_9 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_9__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_9__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_10 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_9__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_10__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_10__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_11 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_10__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_11__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_11__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_11__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign so_x0y0e_L1 = {_i_sw_so_x0y0e_L1_11__o,
        _i_sw_so_x0y0e_L1_10__o,
        _i_sw_so_x0y0e_L1_9__o,
        _i_sw_so_x0y0e_L1_8__o,
        _i_sw_so_x0y0e_L1_7__o,
        _i_sw_so_x0y0e_L1_6__o,
        _i_sw_so_x0y0e_L1_5__o,
        _i_sw_so_x0y0e_L1_4__o,
        _i_sw_so_x0y0e_L1_3__o,
        _i_sw_so_x0y0e_L1_2__o,
        _i_sw_so_x0y0e_L1_1__o,
        _i_sw_so_x0y0e_L1_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_sw_N_ex_n (
    input wire [11:0] bi_u1v1e_L1
    , output wire [11:0] so_u1y0n_L1
    , input wire [11:0] bi_x0v1w_L1
    , input wire [11:0] cu_u1y0n_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_so_u1y0n_L1_0__o;
    wire [0:0] _i_sw_so_u1y0n_L1_1__o;
    wire [0:0] _i_sw_so_u1y0n_L1_2__o;
    wire [0:0] _i_sw_so_u1y0n_L1_3__o;
    wire [0:0] _i_sw_so_u1y0n_L1_4__o;
    wire [0:0] _i_sw_so_u1y0n_L1_5__o;
    wire [0:0] _i_sw_so_u1y0n_L1_6__o;
    wire [0:0] _i_sw_so_u1y0n_L1_7__o;
    wire [0:0] _i_sw_so_u1y0n_L1_8__o;
    wire [0:0] _i_sw_so_u1y0n_L1_9__o;
    wire [0:0] _i_sw_so_u1y0n_L1_10__o;
    wire [0:0] _i_sw_so_u1y0n_L1_11__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_4__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_4__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_5__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_5__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_6__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_7__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_8__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_9__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_9__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_10__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_10__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_11__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_11__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw3 i_sw_so_u1y0n_L1_0 (
        .i({cu_u1y0n_L1[0],
            bi_x0v1w_L1[11],
            bi_u1v1e_L1[9]})
        ,.o(_i_sw_so_u1y0n_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_0__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_1 (
        .i({cu_u1y0n_L1[1],
            bi_x0v1w_L1[0],
            bi_u1v1e_L1[10]})
        ,.o(_i_sw_so_u1y0n_L1_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_1__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_2 (
        .i({cu_u1y0n_L1[2],
            bi_x0v1w_L1[1],
            bi_u1v1e_L1[11]})
        ,.o(_i_sw_so_u1y0n_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_2__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_3 (
        .i({cu_u1y0n_L1[3],
            bi_x0v1w_L1[2],
            bi_u1v1e_L1[0]})
        ,.o(_i_sw_so_u1y0n_L1_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_3__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_4 (
        .i({cu_u1y0n_L1[4],
            bi_x0v1w_L1[3],
            bi_u1v1e_L1[1]})
        ,.o(_i_sw_so_u1y0n_L1_4__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_4__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_5 (
        .i({cu_u1y0n_L1[5],
            bi_x0v1w_L1[4],
            bi_u1v1e_L1[2]})
        ,.o(_i_sw_so_u1y0n_L1_5__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_5__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_6 (
        .i({cu_u1y0n_L1[6],
            bi_x0v1w_L1[5],
            bi_u1v1e_L1[3]})
        ,.o(_i_sw_so_u1y0n_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_6__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_7 (
        .i({cu_u1y0n_L1[7],
            bi_x0v1w_L1[6],
            bi_u1v1e_L1[4]})
        ,.o(_i_sw_so_u1y0n_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_7__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_8 (
        .i({cu_u1y0n_L1[8],
            bi_x0v1w_L1[7],
            bi_u1v1e_L1[5]})
        ,.o(_i_sw_so_u1y0n_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_8__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_9 (
        .i({cu_u1y0n_L1[9],
            bi_x0v1w_L1[8],
            bi_u1v1e_L1[6]})
        ,.o(_i_sw_so_u1y0n_L1_9__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_9__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_10 (
        .i({cu_u1y0n_L1[10],
            bi_x0v1w_L1[9],
            bi_u1v1e_L1[7]})
        ,.o(_i_sw_so_u1y0n_L1_10__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_10__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_11 (
        .i({cu_u1y0n_L1[11],
            bi_x0v1w_L1[10],
            bi_u1v1e_L1[8]})
        ,.o(_i_sw_so_u1y0n_L1_11__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_11__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_3__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_4 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_4__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_4__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_5 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_4__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_5__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_5__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_5__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_6__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_7__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_8__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_9 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_9__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_9__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_10 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_9__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_10__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_10__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_11 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_10__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_11__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_11__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_11__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign so_u1y0n_L1 = {_i_sw_so_u1y0n_L1_11__o,
        _i_sw_so_u1y0n_L1_10__o,
        _i_sw_so_u1y0n_L1_9__o,
        _i_sw_so_u1y0n_L1_8__o,
        _i_sw_so_u1y0n_L1_7__o,
        _i_sw_so_u1y0n_L1_6__o,
        _i_sw_so_u1y0n_L1_5__o,
        _i_sw_so_u1y0n_L1_4__o,
        _i_sw_so_u1y0n_L1_3__o,
        _i_sw_so_u1y0n_L1_2__o,
        _i_sw_so_u1y0n_L1_1__o,
        _i_sw_so_u1y0n_L1_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_sw_N (
    input wire [11:0] bi_u1v1n_L1
    , output wire [11:0] so_u1y0n_L1
    , input wire [11:0] bi_u1v1e_L1
    , input wire [11:0] bi_x0v1w_L1
    , input wire [11:0] cu_u1y0n_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_so_u1y0n_L1_0__o;
    wire [0:0] _i_sw_so_u1y0n_L1_1__o;
    wire [0:0] _i_sw_so_u1y0n_L1_2__o;
    wire [0:0] _i_sw_so_u1y0n_L1_3__o;
    wire [0:0] _i_sw_so_u1y0n_L1_4__o;
    wire [0:0] _i_sw_so_u1y0n_L1_5__o;
    wire [0:0] _i_sw_so_u1y0n_L1_6__o;
    wire [0:0] _i_sw_so_u1y0n_L1_7__o;
    wire [0:0] _i_sw_so_u1y0n_L1_8__o;
    wire [0:0] _i_sw_so_u1y0n_L1_9__o;
    wire [0:0] _i_sw_so_u1y0n_L1_10__o;
    wire [0:0] _i_sw_so_u1y0n_L1_11__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_0__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_u1y0n_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_1__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_u1y0n_L1_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_2__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_u1y0n_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_3__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_u1y0n_L1_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_4__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_u1y0n_L1_4__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_5__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_u1y0n_L1_5__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_6__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_u1y0n_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_7__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_u1y0n_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_8__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_u1y0n_L1_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_9__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_u1y0n_L1_9__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_10__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_u1y0n_L1_10__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_11__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_u1y0n_L1_11__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw4 i_sw_so_u1y0n_L1_0 (
        .i({cu_u1y0n_L1[0],
            bi_x0v1w_L1[11],
            bi_u1v1e_L1[9],
            bi_u1v1n_L1[0]})
        ,.o(_i_sw_so_u1y0n_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_0__prog_data)
        );
    sw4 i_sw_so_u1y0n_L1_1 (
        .i({cu_u1y0n_L1[1],
            bi_x0v1w_L1[0],
            bi_u1v1e_L1[10],
            bi_u1v1n_L1[1]})
        ,.o(_i_sw_so_u1y0n_L1_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_1__prog_data)
        );
    sw4 i_sw_so_u1y0n_L1_2 (
        .i({cu_u1y0n_L1[2],
            bi_x0v1w_L1[1],
            bi_u1v1e_L1[11],
            bi_u1v1n_L1[2]})
        ,.o(_i_sw_so_u1y0n_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_2__prog_data)
        );
    sw4 i_sw_so_u1y0n_L1_3 (
        .i({cu_u1y0n_L1[3],
            bi_x0v1w_L1[2],
            bi_u1v1e_L1[0],
            bi_u1v1n_L1[3]})
        ,.o(_i_sw_so_u1y0n_L1_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_3__prog_data)
        );
    sw4 i_sw_so_u1y0n_L1_4 (
        .i({cu_u1y0n_L1[4],
            bi_x0v1w_L1[3],
            bi_u1v1e_L1[1],
            bi_u1v1n_L1[4]})
        ,.o(_i_sw_so_u1y0n_L1_4__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_4__prog_data)
        );
    sw4 i_sw_so_u1y0n_L1_5 (
        .i({cu_u1y0n_L1[5],
            bi_x0v1w_L1[4],
            bi_u1v1e_L1[2],
            bi_u1v1n_L1[5]})
        ,.o(_i_sw_so_u1y0n_L1_5__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_5__prog_data)
        );
    sw4 i_sw_so_u1y0n_L1_6 (
        .i({cu_u1y0n_L1[6],
            bi_x0v1w_L1[5],
            bi_u1v1e_L1[3],
            bi_u1v1n_L1[6]})
        ,.o(_i_sw_so_u1y0n_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_6__prog_data)
        );
    sw4 i_sw_so_u1y0n_L1_7 (
        .i({cu_u1y0n_L1[7],
            bi_x0v1w_L1[6],
            bi_u1v1e_L1[4],
            bi_u1v1n_L1[7]})
        ,.o(_i_sw_so_u1y0n_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_7__prog_data)
        );
    sw4 i_sw_so_u1y0n_L1_8 (
        .i({cu_u1y0n_L1[8],
            bi_x0v1w_L1[7],
            bi_u1v1e_L1[5],
            bi_u1v1n_L1[8]})
        ,.o(_i_sw_so_u1y0n_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_8__prog_data)
        );
    sw4 i_sw_so_u1y0n_L1_9 (
        .i({cu_u1y0n_L1[9],
            bi_x0v1w_L1[8],
            bi_u1v1e_L1[6],
            bi_u1v1n_L1[9]})
        ,.o(_i_sw_so_u1y0n_L1_9__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_9__prog_data)
        );
    sw4 i_sw_so_u1y0n_L1_10 (
        .i({cu_u1y0n_L1[10],
            bi_x0v1w_L1[9],
            bi_u1v1e_L1[7],
            bi_u1v1n_L1[10]})
        ,.o(_i_sw_so_u1y0n_L1_10__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_10__prog_data)
        );
    sw4 i_sw_so_u1y0n_L1_11 (
        .i({cu_u1y0n_L1[11],
            bi_x0v1w_L1[10],
            bi_u1v1e_L1[8],
            bi_u1v1n_L1[11]})
        ,.o(_i_sw_so_u1y0n_L1_11__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_11__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_u1y0n_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_0__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_u1y0n_L1_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_1__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_u1y0n_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_2__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_u1y0n_L1_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_3__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_u1y0n_L1_4 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_4__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_4__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_u1y0n_L1_5 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_4__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_5__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_5__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_u1y0n_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_5__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_6__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_u1y0n_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_7__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_u1y0n_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_8__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_u1y0n_L1_9 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_9__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_9__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_u1y0n_L1_10 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_9__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_10__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_10__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_u1y0n_L1_11 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_10__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_11__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_11__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_11__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign so_u1y0n_L1 = {_i_sw_so_u1y0n_L1_11__o,
        _i_sw_so_u1y0n_L1_10__o,
        _i_sw_so_u1y0n_L1_9__o,
        _i_sw_so_u1y0n_L1_8__o,
        _i_sw_so_u1y0n_L1_7__o,
        _i_sw_so_u1y0n_L1_6__o,
        _i_sw_so_u1y0n_L1_5__o,
        _i_sw_so_u1y0n_L1_4__o,
        _i_sw_so_u1y0n_L1_3__o,
        _i_sw_so_u1y0n_L1_2__o,
        _i_sw_so_u1y0n_L1_1__o,
        _i_sw_so_u1y0n_L1_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_nw_E_ex_s (
    input wire [11:0] bi_u1y0n_L1
    , output wire [11:0] so_x0y0e_L1
    , input wire [11:0] bi_u1y0e_L1
    , input wire [11:0] cu_x0y0e_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_so_x0y0e_L1_0__o;
    wire [0:0] _i_sw_so_x0y0e_L1_1__o;
    wire [0:0] _i_sw_so_x0y0e_L1_2__o;
    wire [0:0] _i_sw_so_x0y0e_L1_3__o;
    wire [0:0] _i_sw_so_x0y0e_L1_4__o;
    wire [0:0] _i_sw_so_x0y0e_L1_5__o;
    wire [0:0] _i_sw_so_x0y0e_L1_6__o;
    wire [0:0] _i_sw_so_x0y0e_L1_7__o;
    wire [0:0] _i_sw_so_x0y0e_L1_8__o;
    wire [0:0] _i_sw_so_x0y0e_L1_9__o;
    wire [0:0] _i_sw_so_x0y0e_L1_10__o;
    wire [0:0] _i_sw_so_x0y0e_L1_11__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_4__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_4__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_5__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_5__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_6__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_7__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_8__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_9__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_9__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_10__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_10__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0e_L1_11__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0e_L1_11__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw2 i_sw_so_x0y0e_L1_0 (
        .i({cu_x0y0e_L1[0],
            bi_u1y0e_L1[0]})
        ,.o(_i_sw_so_x0y0e_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_0__prog_data)
        );
    sw3 i_sw_so_x0y0e_L1_1 (
        .i({cu_x0y0e_L1[1],
            bi_u1y0e_L1[1],
            bi_u1y0n_L1[3]})
        ,.o(_i_sw_so_x0y0e_L1_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_1__prog_data)
        );
    sw3 i_sw_so_x0y0e_L1_2 (
        .i({cu_x0y0e_L1[2],
            bi_u1y0e_L1[2],
            bi_u1y0n_L1[4]})
        ,.o(_i_sw_so_x0y0e_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_2__prog_data)
        );
    sw3 i_sw_so_x0y0e_L1_3 (
        .i({cu_x0y0e_L1[3],
            bi_u1y0e_L1[3],
            bi_u1y0n_L1[5]})
        ,.o(_i_sw_so_x0y0e_L1_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_3__prog_data)
        );
    sw3 i_sw_so_x0y0e_L1_4 (
        .i({cu_x0y0e_L1[4],
            bi_u1y0e_L1[4],
            bi_u1y0n_L1[6]})
        ,.o(_i_sw_so_x0y0e_L1_4__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_4__prog_data)
        );
    sw3 i_sw_so_x0y0e_L1_5 (
        .i({cu_x0y0e_L1[5],
            bi_u1y0e_L1[5],
            bi_u1y0n_L1[7]})
        ,.o(_i_sw_so_x0y0e_L1_5__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_5__prog_data)
        );
    sw3 i_sw_so_x0y0e_L1_6 (
        .i({cu_x0y0e_L1[6],
            bi_u1y0e_L1[6],
            bi_u1y0n_L1[8]})
        ,.o(_i_sw_so_x0y0e_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_6__prog_data)
        );
    sw3 i_sw_so_x0y0e_L1_7 (
        .i({cu_x0y0e_L1[7],
            bi_u1y0e_L1[7],
            bi_u1y0n_L1[9]})
        ,.o(_i_sw_so_x0y0e_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_7__prog_data)
        );
    sw3 i_sw_so_x0y0e_L1_8 (
        .i({cu_x0y0e_L1[8],
            bi_u1y0e_L1[8],
            bi_u1y0n_L1[10]})
        ,.o(_i_sw_so_x0y0e_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_8__prog_data)
        );
    sw3 i_sw_so_x0y0e_L1_9 (
        .i({cu_x0y0e_L1[9],
            bi_u1y0e_L1[9],
            bi_u1y0n_L1[11]})
        ,.o(_i_sw_so_x0y0e_L1_9__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_9__prog_data)
        );
    sw3 i_sw_so_x0y0e_L1_10 (
        .i({cu_x0y0e_L1[10],
            bi_u1y0e_L1[10],
            bi_u1y0n_L1[0]})
        ,.o(_i_sw_so_x0y0e_L1_10__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_10__prog_data)
        );
    sw3 i_sw_so_x0y0e_L1_11 (
        .i({cu_x0y0e_L1[11],
            bi_u1y0e_L1[11],
            bi_u1y0n_L1[1]})
        ,.o(_i_sw_so_x0y0e_L1_11__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_11__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_3__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_4 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_4__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_4__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_5 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_4__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_5__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_5__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_5__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_6__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_7__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_8__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_9 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_9__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_9__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_10 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_9__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_10__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_10__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0e_L1_11 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_10__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0e_L1_11__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0e_L1_11__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0e_L1_11__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign so_x0y0e_L1 = {_i_sw_so_x0y0e_L1_11__o,
        _i_sw_so_x0y0e_L1_10__o,
        _i_sw_so_x0y0e_L1_9__o,
        _i_sw_so_x0y0e_L1_8__o,
        _i_sw_so_x0y0e_L1_7__o,
        _i_sw_so_x0y0e_L1_6__o,
        _i_sw_so_x0y0e_L1_5__o,
        _i_sw_so_x0y0e_L1_4__o,
        _i_sw_so_x0y0e_L1_3__o,
        _i_sw_so_x0y0e_L1_2__o,
        _i_sw_so_x0y0e_L1_1__o,
        _i_sw_so_x0y0e_L1_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_sw_s_ex_s (
    input wire [11:0] bi_u1v1e_L1
    , input wire [11:0] bi_x0v1w_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    );
    
        
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
        
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
        

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_ne_n_ex_nw (
    input wire [11:0] bi_x0y0e_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    );
    
        
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
        
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
        

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_ne_S_ex_w (
    input wire [11:0] bi_x0y0e_L1
    , output wire [11:0] so_x0y0s_L1
    , input wire [11:0] bi_x0y1s_L1
    , input wire [11:0] cu_x0y0s_L1
    , input wire [11:0] cv_x0y0s_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_so_x0y0s_L1_0__o;
    wire [0:0] _i_sw_so_x0y0s_L1_1__o;
    wire [0:0] _i_sw_so_x0y0s_L1_2__o;
    wire [0:0] _i_sw_so_x0y0s_L1_3__o;
    wire [0:0] _i_sw_so_x0y0s_L1_4__o;
    wire [0:0] _i_sw_so_x0y0s_L1_5__o;
    wire [0:0] _i_sw_so_x0y0s_L1_6__o;
    wire [0:0] _i_sw_so_x0y0s_L1_7__o;
    wire [0:0] _i_sw_so_x0y0s_L1_8__o;
    wire [0:0] _i_sw_so_x0y0s_L1_9__o;
    wire [0:0] _i_sw_so_x0y0s_L1_10__o;
    wire [0:0] _i_sw_so_x0y0s_L1_11__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_0__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_x0y0s_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_1__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_x0y0s_L1_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_2__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_x0y0s_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_3__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_x0y0s_L1_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_4__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_x0y0s_L1_4__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_5__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_x0y0s_L1_5__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_6__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_x0y0s_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_7__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_x0y0s_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_8__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_x0y0s_L1_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_9__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_x0y0s_L1_9__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_10__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_x0y0s_L1_10__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_11__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_x0y0s_L1_11__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw4 i_sw_so_x0y0s_L1_0 (
        .i({cv_x0y0s_L1[0],
            cu_x0y0s_L1[0],
            bi_x0y1s_L1[0],
            bi_x0y0e_L1[11]})
        ,.o(_i_sw_so_x0y0s_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_0__prog_data)
        );
    sw4 i_sw_so_x0y0s_L1_1 (
        .i({cv_x0y0s_L1[1],
            cu_x0y0s_L1[1],
            bi_x0y1s_L1[1],
            bi_x0y0e_L1[0]})
        ,.o(_i_sw_so_x0y0s_L1_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_1__prog_data)
        );
    sw4 i_sw_so_x0y0s_L1_2 (
        .i({cv_x0y0s_L1[2],
            cu_x0y0s_L1[2],
            bi_x0y1s_L1[2],
            bi_x0y0e_L1[1]})
        ,.o(_i_sw_so_x0y0s_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_2__prog_data)
        );
    sw4 i_sw_so_x0y0s_L1_3 (
        .i({cv_x0y0s_L1[3],
            cu_x0y0s_L1[3],
            bi_x0y1s_L1[3],
            bi_x0y0e_L1[2]})
        ,.o(_i_sw_so_x0y0s_L1_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_3__prog_data)
        );
    sw4 i_sw_so_x0y0s_L1_4 (
        .i({cv_x0y0s_L1[4],
            cu_x0y0s_L1[4],
            bi_x0y1s_L1[4],
            bi_x0y0e_L1[3]})
        ,.o(_i_sw_so_x0y0s_L1_4__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_4__prog_data)
        );
    sw4 i_sw_so_x0y0s_L1_5 (
        .i({cv_x0y0s_L1[5],
            cu_x0y0s_L1[5],
            bi_x0y1s_L1[5],
            bi_x0y0e_L1[4]})
        ,.o(_i_sw_so_x0y0s_L1_5__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_5__prog_data)
        );
    sw4 i_sw_so_x0y0s_L1_6 (
        .i({cv_x0y0s_L1[6],
            cu_x0y0s_L1[6],
            bi_x0y1s_L1[6],
            bi_x0y0e_L1[5]})
        ,.o(_i_sw_so_x0y0s_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_6__prog_data)
        );
    sw4 i_sw_so_x0y0s_L1_7 (
        .i({cv_x0y0s_L1[7],
            cu_x0y0s_L1[7],
            bi_x0y1s_L1[7],
            bi_x0y0e_L1[6]})
        ,.o(_i_sw_so_x0y0s_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_7__prog_data)
        );
    sw4 i_sw_so_x0y0s_L1_8 (
        .i({cv_x0y0s_L1[8],
            cu_x0y0s_L1[8],
            bi_x0y1s_L1[8],
            bi_x0y0e_L1[7]})
        ,.o(_i_sw_so_x0y0s_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_8__prog_data)
        );
    sw4 i_sw_so_x0y0s_L1_9 (
        .i({cv_x0y0s_L1[9],
            cu_x0y0s_L1[9],
            bi_x0y1s_L1[9],
            bi_x0y0e_L1[8]})
        ,.o(_i_sw_so_x0y0s_L1_9__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_9__prog_data)
        );
    sw4 i_sw_so_x0y0s_L1_10 (
        .i({cv_x0y0s_L1[10],
            cu_x0y0s_L1[10],
            bi_x0y1s_L1[10],
            bi_x0y0e_L1[9]})
        ,.o(_i_sw_so_x0y0s_L1_10__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_10__prog_data)
        );
    sw4 i_sw_so_x0y0s_L1_11 (
        .i({cv_x0y0s_L1[11],
            cu_x0y0s_L1[11],
            bi_x0y1s_L1[11],
            bi_x0y0e_L1[10]})
        ,.o(_i_sw_so_x0y0s_L1_11__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_11__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_x0y0s_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_0__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_x0y0s_L1_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_1__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_x0y0s_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_2__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_x0y0s_L1_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_3__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_x0y0s_L1_4 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_4__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_4__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_x0y0s_L1_5 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_4__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_5__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_5__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_x0y0s_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_5__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_6__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_x0y0s_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_7__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_x0y0s_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_8__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_x0y0s_L1_9 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_9__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_9__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_x0y0s_L1_10 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_9__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_10__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_10__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_x0y0s_L1_11 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_10__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_11__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_11__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_11__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign so_x0y0s_L1 = {_i_sw_so_x0y0s_L1_11__o,
        _i_sw_so_x0y0s_L1_10__o,
        _i_sw_so_x0y0s_L1_9__o,
        _i_sw_so_x0y0s_L1_8__o,
        _i_sw_so_x0y0s_L1_7__o,
        _i_sw_so_x0y0s_L1_6__o,
        _i_sw_so_x0y0s_L1_5__o,
        _i_sw_so_x0y0s_L1_4__o,
        _i_sw_so_x0y0s_L1_3__o,
        _i_sw_so_x0y0s_L1_2__o,
        _i_sw_so_x0y0s_L1_1__o,
        _i_sw_so_x0y0s_L1_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_se_W_ex_nw (
    input wire [11:0] bi_x0y0s_L1
    , output wire [11:0] so_x0v1w_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_so_x0v1w_L1_0__o;
    wire [0:0] _i_sw_so_x0v1w_L1_1__o;
    wire [0:0] _i_sw_so_x0v1w_L1_2__o;
    wire [0:0] _i_sw_so_x0v1w_L1_3__o;
    wire [0:0] _i_sw_so_x0v1w_L1_4__o;
    wire [0:0] _i_sw_so_x0v1w_L1_5__o;
    wire [0:0] _i_sw_so_x0v1w_L1_6__o;
    wire [0:0] _i_sw_so_x0v1w_L1_7__o;
    wire [0:0] _i_sw_so_x0v1w_L1_8__o;
    wire [0:0] _i_sw_so_x0v1w_L1_9__o;
    wire [0:0] _i_sw_so_x0v1w_L1_10__o;
    wire [0:0] _i_sw_so_x0v1w_L1_11__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_0__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_1__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_2__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_3__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_4__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_4__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_5__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_5__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_6__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_7__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_8__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_9__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_9__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_10__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_10__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_11__prog_dout;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_11__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw1 i_sw_so_x0v1w_L1_0 (
        .i(bi_x0y0s_L1[11])
        ,.o(_i_sw_so_x0v1w_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_0__prog_data)
        );
    sw1 i_sw_so_x0v1w_L1_1 (
        .i(bi_x0y0s_L1[0])
        ,.o(_i_sw_so_x0v1w_L1_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_1__prog_data)
        );
    sw1 i_sw_so_x0v1w_L1_2 (
        .i(bi_x0y0s_L1[1])
        ,.o(_i_sw_so_x0v1w_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_2__prog_data)
        );
    sw1 i_sw_so_x0v1w_L1_3 (
        .i(bi_x0y0s_L1[2])
        ,.o(_i_sw_so_x0v1w_L1_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_3__prog_data)
        );
    sw1 i_sw_so_x0v1w_L1_4 (
        .i(bi_x0y0s_L1[3])
        ,.o(_i_sw_so_x0v1w_L1_4__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_4__prog_data)
        );
    sw1 i_sw_so_x0v1w_L1_5 (
        .i(bi_x0y0s_L1[4])
        ,.o(_i_sw_so_x0v1w_L1_5__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_5__prog_data)
        );
    sw1 i_sw_so_x0v1w_L1_6 (
        .i(bi_x0y0s_L1[5])
        ,.o(_i_sw_so_x0v1w_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_6__prog_data)
        );
    sw1 i_sw_so_x0v1w_L1_7 (
        .i(bi_x0y0s_L1[6])
        ,.o(_i_sw_so_x0v1w_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_7__prog_data)
        );
    sw1 i_sw_so_x0v1w_L1_8 (
        .i(bi_x0y0s_L1[7])
        ,.o(_i_sw_so_x0v1w_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_8__prog_data)
        );
    sw1 i_sw_so_x0v1w_L1_9 (
        .i(bi_x0y0s_L1[8])
        ,.o(_i_sw_so_x0v1w_L1_9__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_9__prog_data)
        );
    sw1 i_sw_so_x0v1w_L1_10 (
        .i(bi_x0y0s_L1[9])
        ,.o(_i_sw_so_x0v1w_L1_10__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_10__prog_data)
        );
    sw1 i_sw_so_x0v1w_L1_11 (
        .i(bi_x0y0s_L1[10])
        ,.o(_i_sw_so_x0v1w_L1_11__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_11__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0v1w_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_0__prog_data)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0v1w_L1_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_1__prog_data)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0v1w_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_2__prog_data)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0v1w_L1_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_3__prog_data)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0v1w_L1_4 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_4__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_4__prog_data)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0v1w_L1_5 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_4__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_5__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_5__prog_data)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0v1w_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_5__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_6__prog_data)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0v1w_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_7__prog_data)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0v1w_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_8__prog_data)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0v1w_L1_9 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_9__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_9__prog_data)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0v1w_L1_10 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_9__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_10__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_10__prog_data)
        );
    scanchain_data_d1 i_prog_data_i_sw_so_x0v1w_L1_11 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_10__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_11__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_11__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_11__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign so_x0v1w_L1 = {_i_sw_so_x0v1w_L1_11__o,
        _i_sw_so_x0v1w_L1_10__o,
        _i_sw_so_x0v1w_L1_9__o,
        _i_sw_so_x0v1w_L1_8__o,
        _i_sw_so_x0v1w_L1_7__o,
        _i_sw_so_x0v1w_L1_6__o,
        _i_sw_so_x0v1w_L1_5__o,
        _i_sw_so_x0v1w_L1_4__o,
        _i_sw_so_x0v1w_L1_3__o,
        _i_sw_so_x0v1w_L1_2__o,
        _i_sw_so_x0v1w_L1_1__o,
        _i_sw_so_x0v1w_L1_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_se_W_ex_w (
    input wire [11:0] bi_x0v1n_L1
    , output wire [11:0] so_x0v1w_L1
    , input wire [11:0] bi_x0y0s_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_so_x0v1w_L1_0__o;
    wire [0:0] _i_sw_so_x0v1w_L1_1__o;
    wire [0:0] _i_sw_so_x0v1w_L1_2__o;
    wire [0:0] _i_sw_so_x0v1w_L1_3__o;
    wire [0:0] _i_sw_so_x0v1w_L1_4__o;
    wire [0:0] _i_sw_so_x0v1w_L1_5__o;
    wire [0:0] _i_sw_so_x0v1w_L1_6__o;
    wire [0:0] _i_sw_so_x0v1w_L1_7__o;
    wire [0:0] _i_sw_so_x0v1w_L1_8__o;
    wire [0:0] _i_sw_so_x0v1w_L1_9__o;
    wire [0:0] _i_sw_so_x0v1w_L1_10__o;
    wire [0:0] _i_sw_so_x0v1w_L1_11__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_4__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_4__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_5__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_5__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_6__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_7__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_8__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_9__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_9__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_10__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_10__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_11__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_11__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw2 i_sw_so_x0v1w_L1_0 (
        .i({bi_x0y0s_L1[11],
            bi_x0v1n_L1[1]})
        ,.o(_i_sw_so_x0v1w_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_0__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_1 (
        .i({bi_x0y0s_L1[0],
            bi_x0v1n_L1[2]})
        ,.o(_i_sw_so_x0v1w_L1_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_1__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_2 (
        .i({bi_x0y0s_L1[1],
            bi_x0v1n_L1[3]})
        ,.o(_i_sw_so_x0v1w_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_2__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_3 (
        .i({bi_x0y0s_L1[2],
            bi_x0v1n_L1[4]})
        ,.o(_i_sw_so_x0v1w_L1_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_3__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_4 (
        .i({bi_x0y0s_L1[3],
            bi_x0v1n_L1[5]})
        ,.o(_i_sw_so_x0v1w_L1_4__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_4__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_5 (
        .i({bi_x0y0s_L1[4],
            bi_x0v1n_L1[6]})
        ,.o(_i_sw_so_x0v1w_L1_5__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_5__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_6 (
        .i({bi_x0y0s_L1[5],
            bi_x0v1n_L1[7]})
        ,.o(_i_sw_so_x0v1w_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_6__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_7 (
        .i({bi_x0y0s_L1[6],
            bi_x0v1n_L1[8]})
        ,.o(_i_sw_so_x0v1w_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_7__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_8 (
        .i({bi_x0y0s_L1[7],
            bi_x0v1n_L1[9]})
        ,.o(_i_sw_so_x0v1w_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_8__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_9 (
        .i({bi_x0y0s_L1[8],
            bi_x0v1n_L1[10]})
        ,.o(_i_sw_so_x0v1w_L1_9__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_9__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_10 (
        .i({bi_x0y0s_L1[9],
            bi_x0v1n_L1[11]})
        ,.o(_i_sw_so_x0v1w_L1_10__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_10__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_11 (
        .i({bi_x0y0s_L1[10],
            bi_x0v1n_L1[0]})
        ,.o(_i_sw_so_x0v1w_L1_11__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_11__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_3__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_4 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_4__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_4__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_5 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_4__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_5__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_5__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_5__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_6__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_7__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_8__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_9 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_9__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_9__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_10 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_9__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_10__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_10__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_11 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_10__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_11__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_11__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_11__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign so_x0v1w_L1 = {_i_sw_so_x0v1w_L1_11__o,
        _i_sw_so_x0v1w_L1_10__o,
        _i_sw_so_x0v1w_L1_9__o,
        _i_sw_so_x0v1w_L1_8__o,
        _i_sw_so_x0v1w_L1_7__o,
        _i_sw_so_x0v1w_L1_6__o,
        _i_sw_so_x0v1w_L1_5__o,
        _i_sw_so_x0v1w_L1_4__o,
        _i_sw_so_x0v1w_L1_3__o,
        _i_sw_so_x0v1w_L1_2__o,
        _i_sw_so_x0v1w_L1_1__o,
        _i_sw_so_x0v1w_L1_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_ne_S_ex_sw (
    input wire [11:0] bi_x0y0e_L1
    , output wire [11:0] so_x0y0s_L1
    , input wire [11:0] cu_x0y0s_L1
    , input wire [11:0] cv_x0y0s_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_so_x0y0s_L1_0__o;
    wire [0:0] _i_sw_so_x0y0s_L1_1__o;
    wire [0:0] _i_sw_so_x0y0s_L1_2__o;
    wire [0:0] _i_sw_so_x0y0s_L1_3__o;
    wire [0:0] _i_sw_so_x0y0s_L1_4__o;
    wire [0:0] _i_sw_so_x0y0s_L1_5__o;
    wire [0:0] _i_sw_so_x0y0s_L1_6__o;
    wire [0:0] _i_sw_so_x0y0s_L1_7__o;
    wire [0:0] _i_sw_so_x0y0s_L1_8__o;
    wire [0:0] _i_sw_so_x0y0s_L1_9__o;
    wire [0:0] _i_sw_so_x0y0s_L1_10__o;
    wire [0:0] _i_sw_so_x0y0s_L1_11__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_4__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_4__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_5__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_5__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_6__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_7__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_8__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_9__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_9__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_10__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_10__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0y0s_L1_11__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0y0s_L1_11__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw3 i_sw_so_x0y0s_L1_0 (
        .i({cv_x0y0s_L1[0],
            cu_x0y0s_L1[0],
            bi_x0y0e_L1[11]})
        ,.o(_i_sw_so_x0y0s_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_0__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_1 (
        .i({cv_x0y0s_L1[1],
            cu_x0y0s_L1[1],
            bi_x0y0e_L1[0]})
        ,.o(_i_sw_so_x0y0s_L1_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_1__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_2 (
        .i({cv_x0y0s_L1[2],
            cu_x0y0s_L1[2],
            bi_x0y0e_L1[1]})
        ,.o(_i_sw_so_x0y0s_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_2__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_3 (
        .i({cv_x0y0s_L1[3],
            cu_x0y0s_L1[3],
            bi_x0y0e_L1[2]})
        ,.o(_i_sw_so_x0y0s_L1_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_3__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_4 (
        .i({cv_x0y0s_L1[4],
            cu_x0y0s_L1[4],
            bi_x0y0e_L1[3]})
        ,.o(_i_sw_so_x0y0s_L1_4__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_4__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_5 (
        .i({cv_x0y0s_L1[5],
            cu_x0y0s_L1[5],
            bi_x0y0e_L1[4]})
        ,.o(_i_sw_so_x0y0s_L1_5__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_5__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_6 (
        .i({cv_x0y0s_L1[6],
            cu_x0y0s_L1[6],
            bi_x0y0e_L1[5]})
        ,.o(_i_sw_so_x0y0s_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_6__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_7 (
        .i({cv_x0y0s_L1[7],
            cu_x0y0s_L1[7],
            bi_x0y0e_L1[6]})
        ,.o(_i_sw_so_x0y0s_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_7__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_8 (
        .i({cv_x0y0s_L1[8],
            cu_x0y0s_L1[8],
            bi_x0y0e_L1[7]})
        ,.o(_i_sw_so_x0y0s_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_8__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_9 (
        .i({cv_x0y0s_L1[9],
            cu_x0y0s_L1[9],
            bi_x0y0e_L1[8]})
        ,.o(_i_sw_so_x0y0s_L1_9__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_9__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_10 (
        .i({cv_x0y0s_L1[10],
            cu_x0y0s_L1[10],
            bi_x0y0e_L1[9]})
        ,.o(_i_sw_so_x0y0s_L1_10__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_10__prog_data)
        );
    sw3 i_sw_so_x0y0s_L1_11 (
        .i({cv_x0y0s_L1[11],
            cu_x0y0s_L1[11],
            bi_x0y0e_L1[10]})
        ,.o(_i_sw_so_x0y0s_L1_11__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_11__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_3__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_4 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_4__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_4__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_5 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_4__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_5__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_5__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_5__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_6__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_7__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_8__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_9 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_9__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_9__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_10 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_9__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_10__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_10__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0y0s_L1_11 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_10__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0y0s_L1_11__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0y0s_L1_11__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0y0s_L1_11__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign so_x0y0s_L1 = {_i_sw_so_x0y0s_L1_11__o,
        _i_sw_so_x0y0s_L1_10__o,
        _i_sw_so_x0y0s_L1_9__o,
        _i_sw_so_x0y0s_L1_8__o,
        _i_sw_so_x0y0s_L1_7__o,
        _i_sw_so_x0y0s_L1_6__o,
        _i_sw_so_x0y0s_L1_5__o,
        _i_sw_so_x0y0s_L1_4__o,
        _i_sw_so_x0y0s_L1_3__o,
        _i_sw_so_x0y0s_L1_2__o,
        _i_sw_so_x0y0s_L1_1__o,
        _i_sw_so_x0y0s_L1_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_se_W_ex_sw (
    input wire [11:0] bi_x0v1n_L1
    , output wire [11:0] so_x0v1w_L1
    , input wire [11:0] cu_x0v1w_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_so_x0v1w_L1_0__o;
    wire [0:0] _i_sw_so_x0v1w_L1_1__o;
    wire [0:0] _i_sw_so_x0v1w_L1_2__o;
    wire [0:0] _i_sw_so_x0v1w_L1_3__o;
    wire [0:0] _i_sw_so_x0v1w_L1_4__o;
    wire [0:0] _i_sw_so_x0v1w_L1_5__o;
    wire [0:0] _i_sw_so_x0v1w_L1_6__o;
    wire [0:0] _i_sw_so_x0v1w_L1_7__o;
    wire [0:0] _i_sw_so_x0v1w_L1_8__o;
    wire [0:0] _i_sw_so_x0v1w_L1_9__o;
    wire [0:0] _i_sw_so_x0v1w_L1_10__o;
    wire [0:0] _i_sw_so_x0v1w_L1_11__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_4__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_4__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_5__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_5__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_6__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_7__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_8__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_9__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_9__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_10__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_10__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_x0v1w_L1_11__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_x0v1w_L1_11__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw2 i_sw_so_x0v1w_L1_0 (
        .i({cu_x0v1w_L1[0],
            bi_x0v1n_L1[1]})
        ,.o(_i_sw_so_x0v1w_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_0__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_1 (
        .i({cu_x0v1w_L1[1],
            bi_x0v1n_L1[2]})
        ,.o(_i_sw_so_x0v1w_L1_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_1__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_2 (
        .i({cu_x0v1w_L1[2],
            bi_x0v1n_L1[3]})
        ,.o(_i_sw_so_x0v1w_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_2__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_3 (
        .i({cu_x0v1w_L1[3],
            bi_x0v1n_L1[4]})
        ,.o(_i_sw_so_x0v1w_L1_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_3__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_4 (
        .i({cu_x0v1w_L1[4],
            bi_x0v1n_L1[5]})
        ,.o(_i_sw_so_x0v1w_L1_4__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_4__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_5 (
        .i({cu_x0v1w_L1[5],
            bi_x0v1n_L1[6]})
        ,.o(_i_sw_so_x0v1w_L1_5__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_5__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_6 (
        .i({cu_x0v1w_L1[6],
            bi_x0v1n_L1[7]})
        ,.o(_i_sw_so_x0v1w_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_6__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_7 (
        .i({cu_x0v1w_L1[7],
            bi_x0v1n_L1[8]})
        ,.o(_i_sw_so_x0v1w_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_7__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_8 (
        .i({cu_x0v1w_L1[8],
            bi_x0v1n_L1[9]})
        ,.o(_i_sw_so_x0v1w_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_8__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_9 (
        .i({cu_x0v1w_L1[9],
            bi_x0v1n_L1[10]})
        ,.o(_i_sw_so_x0v1w_L1_9__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_9__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_10 (
        .i({cu_x0v1w_L1[10],
            bi_x0v1n_L1[11]})
        ,.o(_i_sw_so_x0v1w_L1_10__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_10__prog_data)
        );
    sw2 i_sw_so_x0v1w_L1_11 (
        .i({cu_x0v1w_L1[11],
            bi_x0v1n_L1[0]})
        ,.o(_i_sw_so_x0v1w_L1_11__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_11__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_3__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_4 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_4__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_4__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_5 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_4__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_5__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_5__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_5__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_6__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_7__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_8__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_9 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_9__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_9__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_10 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_9__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_10__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_10__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_x0v1w_L1_11 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_10__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_x0v1w_L1_11__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_x0v1w_L1_11__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_x0v1w_L1_11__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign so_x0v1w_L1 = {_i_sw_so_x0v1w_L1_11__o,
        _i_sw_so_x0v1w_L1_10__o,
        _i_sw_so_x0v1w_L1_9__o,
        _i_sw_so_x0v1w_L1_8__o,
        _i_sw_so_x0v1w_L1_7__o,
        _i_sw_so_x0v1w_L1_6__o,
        _i_sw_so_x0v1w_L1_5__o,
        _i_sw_so_x0v1w_L1_4__o,
        _i_sw_so_x0v1w_L1_3__o,
        _i_sw_so_x0v1w_L1_2__o,
        _i_sw_so_x0v1w_L1_1__o,
        _i_sw_so_x0v1w_L1_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_nw_w_ex_nw (
    input wire [11:0] bi_u1y1s_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    );
    
        
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
        
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
        

endmodule
// Automatically generated by PRGA's RTL generator
module t_io_e (
    input wire [11:0] bi_u1y0n_L1
    , input wire [11:0] bi_u1y0s_L1
    , output wire [11:0] cu_u1y0n_L1
    , output wire [11:0] cu_u1y0s_L1
    , input wire [0:0] ipin_x0y0_0
    , output wire [0:0] opin_x0y0_0
    , output wire [0:0] oe_x0y0_0
    , input wire [0:0] ipin_x0y0_1
    , output wire [0:0] opin_x0y0_1
    , output wire [0:0] oe_x0y0_1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_blk_i0__inpad;
    wire [0:0] _i_blk_i0__opin;
    wire [0:0] _i_blk_i0__oe;
    wire [0:0] _i_blk_i0__prog_dout;
    wire [0:0] _i_blk_i0__prog_we_o;
    wire [0:0] _i_blk_i1__inpad;
    wire [0:0] _i_blk_i1__opin;
    wire [0:0] _i_blk_i1__oe;
    wire [0:0] _i_blk_i1__prog_dout;
    wire [0:0] _i_blk_i1__prog_we_o;
    wire [0:0] _i_cbox_w0__bp_x0y0i0_outpad;
    wire [11:0] _i_cbox_w0__cu_u1y0n_L1;
    wire [11:0] _i_cbox_w0__cu_u1y0s_L1;
    wire [0:0] _i_cbox_w0__bp_x0y0i1_outpad;
    wire [0:0] _i_cbox_w0__prog_dout;
    wire [0:0] _i_cbox_w0__prog_we_o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_buf_prog_rst_l1__Q;
    wire [0:0] _i_buf_prog_done_l1__Q;
        
    iob i_blk_i0 (
        .outpad(_i_cbox_w0__bp_x0y0i0_outpad)
        ,.inpad(_i_blk_i0__inpad)
        ,.ipin(ipin_x0y0_0)
        ,.opin(_i_blk_i0__opin)
        ,.oe(_i_blk_i0__oe)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_blk_i0__prog_dout)
        ,.prog_we_o(_i_blk_i0__prog_we_o)
        );
    iob i_blk_i1 (
        .outpad(_i_cbox_w0__bp_x0y0i1_outpad)
        ,.inpad(_i_blk_i1__inpad)
        ,.ipin(ipin_x0y0_1)
        ,.opin(_i_blk_i1__opin)
        ,.oe(_i_blk_i1__oe)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_blk_i0__prog_we_o)
        ,.prog_din(_i_blk_i0__prog_dout)
        ,.prog_dout(_i_blk_i1__prog_dout)
        ,.prog_we_o(_i_blk_i1__prog_we_o)
        );
    cbox_t_io_e_w0 i_cbox_w0 (
        .bp_x0y0i0_outpad(_i_cbox_w0__bp_x0y0i0_outpad)
        ,.bi_u1y0n_L1(bi_u1y0n_L1)
        ,.bi_u1y0s_L1(bi_u1y0s_L1)
        ,.bp_x0y0i0_inpad(_i_blk_i0__inpad)
        ,.cu_u1y0n_L1(_i_cbox_w0__cu_u1y0n_L1)
        ,.cu_u1y0s_L1(_i_cbox_w0__cu_u1y0s_L1)
        ,.bp_x0y0i1_outpad(_i_cbox_w0__bp_x0y0i1_outpad)
        ,.bp_x0y0i1_inpad(_i_blk_i1__inpad)
        ,.prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l1__Q)
        ,.prog_done(_i_buf_prog_done_l1__Q)
        ,.prog_we(_i_blk_i1__prog_we_o)
        ,.prog_din(_i_blk_i1__prog_dout)
        ,.prog_dout(_i_cbox_w0__prog_dout)
        ,.prog_we_o(_i_cbox_w0__prog_we_o)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(_i_buf_prog_rst_l1__Q)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(_i_buf_prog_done_l1__Q)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    prga_simple_buf i_buf_prog_rst_l1 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l1__Q)
        );
    prga_simple_bufr i_buf_prog_done_l1 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l1__Q)
        );
        
    assign cu_u1y0n_L1 = _i_cbox_w0__cu_u1y0n_L1;
    assign cu_u1y0s_L1 = _i_cbox_w0__cu_u1y0s_L1;
    assign opin_x0y0_0 = _i_blk_i0__opin;
    assign oe_x0y0_0 = _i_blk_i0__oe;
    assign opin_x0y0_1 = _i_blk_i1__opin;
    assign oe_x0y0_1 = _i_blk_i1__oe;
    assign prog_dout = _i_cbox_w0__prog_dout;
    assign prog_we_o = _i_cbox_w0__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_nw_w_ex_w (
    input wire [11:0] bi_u1y0n_L1
    , input wire [11:0] bi_u1y1s_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    );
    
        
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
        
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
        

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_sw_N_ex_nw (
    input wire [11:0] bi_u1v1e_L1
    , output wire [11:0] so_u1y0n_L1
    , input wire [11:0] cu_u1y0n_L1
    , input wire [11:0] cv_u1y0n_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_so_u1y0n_L1_0__o;
    wire [0:0] _i_sw_so_u1y0n_L1_1__o;
    wire [0:0] _i_sw_so_u1y0n_L1_2__o;
    wire [0:0] _i_sw_so_u1y0n_L1_3__o;
    wire [0:0] _i_sw_so_u1y0n_L1_4__o;
    wire [0:0] _i_sw_so_u1y0n_L1_5__o;
    wire [0:0] _i_sw_so_u1y0n_L1_6__o;
    wire [0:0] _i_sw_so_u1y0n_L1_7__o;
    wire [0:0] _i_sw_so_u1y0n_L1_8__o;
    wire [0:0] _i_sw_so_u1y0n_L1_9__o;
    wire [0:0] _i_sw_so_u1y0n_L1_10__o;
    wire [0:0] _i_sw_so_u1y0n_L1_11__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_0__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_1__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_2__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_3__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_4__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_4__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_5__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_5__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_6__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_7__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_8__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_9__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_9__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_10__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_10__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_11__prog_dout;
    wire [1:0] _i_prog_data_i_sw_so_u1y0n_L1_11__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw3 i_sw_so_u1y0n_L1_0 (
        .i({cv_u1y0n_L1[0],
            cu_u1y0n_L1[0],
            bi_u1v1e_L1[9]})
        ,.o(_i_sw_so_u1y0n_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_0__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_1 (
        .i({cv_u1y0n_L1[1],
            cu_u1y0n_L1[1],
            bi_u1v1e_L1[10]})
        ,.o(_i_sw_so_u1y0n_L1_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_1__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_2 (
        .i({cv_u1y0n_L1[2],
            cu_u1y0n_L1[2],
            bi_u1v1e_L1[11]})
        ,.o(_i_sw_so_u1y0n_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_2__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_3 (
        .i({cv_u1y0n_L1[3],
            cu_u1y0n_L1[3],
            bi_u1v1e_L1[0]})
        ,.o(_i_sw_so_u1y0n_L1_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_3__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_4 (
        .i({cv_u1y0n_L1[4],
            cu_u1y0n_L1[4],
            bi_u1v1e_L1[1]})
        ,.o(_i_sw_so_u1y0n_L1_4__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_4__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_5 (
        .i({cv_u1y0n_L1[5],
            cu_u1y0n_L1[5],
            bi_u1v1e_L1[2]})
        ,.o(_i_sw_so_u1y0n_L1_5__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_5__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_6 (
        .i({cv_u1y0n_L1[6],
            cu_u1y0n_L1[6],
            bi_u1v1e_L1[3]})
        ,.o(_i_sw_so_u1y0n_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_6__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_7 (
        .i({cv_u1y0n_L1[7],
            cu_u1y0n_L1[7],
            bi_u1v1e_L1[4]})
        ,.o(_i_sw_so_u1y0n_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_7__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_8 (
        .i({cv_u1y0n_L1[8],
            cu_u1y0n_L1[8],
            bi_u1v1e_L1[5]})
        ,.o(_i_sw_so_u1y0n_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_8__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_9 (
        .i({cv_u1y0n_L1[9],
            cu_u1y0n_L1[9],
            bi_u1v1e_L1[6]})
        ,.o(_i_sw_so_u1y0n_L1_9__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_9__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_10 (
        .i({cv_u1y0n_L1[10],
            cu_u1y0n_L1[10],
            bi_u1v1e_L1[7]})
        ,.o(_i_sw_so_u1y0n_L1_10__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_10__prog_data)
        );
    sw3 i_sw_so_u1y0n_L1_11 (
        .i({cv_u1y0n_L1[11],
            cu_u1y0n_L1[11],
            bi_u1v1e_L1[8]})
        ,.o(_i_sw_so_u1y0n_L1_11__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_11__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_0__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_1__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_2__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_3__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_4 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_4__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_4__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_5 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_4__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_5__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_5__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_5__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_6__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_7__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_8__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_9 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_9__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_9__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_10 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_9__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_10__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_10__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_so_u1y0n_L1_11 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_10__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_11__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_11__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_11__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign so_u1y0n_L1 = {_i_sw_so_u1y0n_L1_11__o,
        _i_sw_so_u1y0n_L1_10__o,
        _i_sw_so_u1y0n_L1_9__o,
        _i_sw_so_u1y0n_L1_8__o,
        _i_sw_so_u1y0n_L1_7__o,
        _i_sw_so_u1y0n_L1_6__o,
        _i_sw_so_u1y0n_L1_5__o,
        _i_sw_so_u1y0n_L1_4__o,
        _i_sw_so_u1y0n_L1_3__o,
        _i_sw_so_u1y0n_L1_2__o,
        _i_sw_so_u1y0n_L1_1__o,
        _i_sw_so_u1y0n_L1_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_sw_N_ex_w (
    input wire [11:0] bi_u1v1n_L1
    , output wire [11:0] so_u1y0n_L1
    , input wire [11:0] bi_u1v1e_L1
    , input wire [11:0] cu_u1y0n_L1
    , input wire [11:0] cv_u1y0n_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_so_u1y0n_L1_0__o;
    wire [0:0] _i_sw_so_u1y0n_L1_1__o;
    wire [0:0] _i_sw_so_u1y0n_L1_2__o;
    wire [0:0] _i_sw_so_u1y0n_L1_3__o;
    wire [0:0] _i_sw_so_u1y0n_L1_4__o;
    wire [0:0] _i_sw_so_u1y0n_L1_5__o;
    wire [0:0] _i_sw_so_u1y0n_L1_6__o;
    wire [0:0] _i_sw_so_u1y0n_L1_7__o;
    wire [0:0] _i_sw_so_u1y0n_L1_8__o;
    wire [0:0] _i_sw_so_u1y0n_L1_9__o;
    wire [0:0] _i_sw_so_u1y0n_L1_10__o;
    wire [0:0] _i_sw_so_u1y0n_L1_11__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_0__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_u1y0n_L1_0__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_1__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_u1y0n_L1_1__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_2__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_u1y0n_L1_2__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_3__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_u1y0n_L1_3__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_4__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_u1y0n_L1_4__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_5__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_u1y0n_L1_5__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_6__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_u1y0n_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_7__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_u1y0n_L1_7__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_8__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_u1y0n_L1_8__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_9__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_u1y0n_L1_9__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_10__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_u1y0n_L1_10__prog_data;
    wire [0:0] _i_prog_data_i_sw_so_u1y0n_L1_11__prog_dout;
    wire [2:0] _i_prog_data_i_sw_so_u1y0n_L1_11__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw4 i_sw_so_u1y0n_L1_0 (
        .i({cv_u1y0n_L1[0],
            cu_u1y0n_L1[0],
            bi_u1v1e_L1[9],
            bi_u1v1n_L1[0]})
        ,.o(_i_sw_so_u1y0n_L1_0__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_0__prog_data)
        );
    sw4 i_sw_so_u1y0n_L1_1 (
        .i({cv_u1y0n_L1[1],
            cu_u1y0n_L1[1],
            bi_u1v1e_L1[10],
            bi_u1v1n_L1[1]})
        ,.o(_i_sw_so_u1y0n_L1_1__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_1__prog_data)
        );
    sw4 i_sw_so_u1y0n_L1_2 (
        .i({cv_u1y0n_L1[2],
            cu_u1y0n_L1[2],
            bi_u1v1e_L1[11],
            bi_u1v1n_L1[2]})
        ,.o(_i_sw_so_u1y0n_L1_2__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_2__prog_data)
        );
    sw4 i_sw_so_u1y0n_L1_3 (
        .i({cv_u1y0n_L1[3],
            cu_u1y0n_L1[3],
            bi_u1v1e_L1[0],
            bi_u1v1n_L1[3]})
        ,.o(_i_sw_so_u1y0n_L1_3__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_3__prog_data)
        );
    sw4 i_sw_so_u1y0n_L1_4 (
        .i({cv_u1y0n_L1[4],
            cu_u1y0n_L1[4],
            bi_u1v1e_L1[1],
            bi_u1v1n_L1[4]})
        ,.o(_i_sw_so_u1y0n_L1_4__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_4__prog_data)
        );
    sw4 i_sw_so_u1y0n_L1_5 (
        .i({cv_u1y0n_L1[5],
            cu_u1y0n_L1[5],
            bi_u1v1e_L1[2],
            bi_u1v1n_L1[5]})
        ,.o(_i_sw_so_u1y0n_L1_5__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_5__prog_data)
        );
    sw4 i_sw_so_u1y0n_L1_6 (
        .i({cv_u1y0n_L1[6],
            cu_u1y0n_L1[6],
            bi_u1v1e_L1[3],
            bi_u1v1n_L1[6]})
        ,.o(_i_sw_so_u1y0n_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_6__prog_data)
        );
    sw4 i_sw_so_u1y0n_L1_7 (
        .i({cv_u1y0n_L1[7],
            cu_u1y0n_L1[7],
            bi_u1v1e_L1[4],
            bi_u1v1n_L1[7]})
        ,.o(_i_sw_so_u1y0n_L1_7__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_7__prog_data)
        );
    sw4 i_sw_so_u1y0n_L1_8 (
        .i({cv_u1y0n_L1[8],
            cu_u1y0n_L1[8],
            bi_u1v1e_L1[5],
            bi_u1v1n_L1[8]})
        ,.o(_i_sw_so_u1y0n_L1_8__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_8__prog_data)
        );
    sw4 i_sw_so_u1y0n_L1_9 (
        .i({cv_u1y0n_L1[9],
            cu_u1y0n_L1[9],
            bi_u1v1e_L1[6],
            bi_u1v1n_L1[9]})
        ,.o(_i_sw_so_u1y0n_L1_9__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_9__prog_data)
        );
    sw4 i_sw_so_u1y0n_L1_10 (
        .i({cv_u1y0n_L1[10],
            cu_u1y0n_L1[10],
            bi_u1v1e_L1[7],
            bi_u1v1n_L1[10]})
        ,.o(_i_sw_so_u1y0n_L1_10__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_10__prog_data)
        );
    sw4 i_sw_so_u1y0n_L1_11 (
        .i({cv_u1y0n_L1[11],
            cu_u1y0n_L1[11],
            bi_u1v1e_L1[8],
            bi_u1v1n_L1[11]})
        ,.o(_i_sw_so_u1y0n_L1_11__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_11__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_u1y0n_L1_0 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_0__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_0__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_u1y0n_L1_1 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_0__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_1__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_1__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_u1y0n_L1_2 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_1__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_2__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_2__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_u1y0n_L1_3 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_2__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_3__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_3__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_u1y0n_L1_4 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_3__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_4__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_4__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_u1y0n_L1_5 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_4__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_5__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_5__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_u1y0n_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_5__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_6__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_u1y0n_L1_7 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_7__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_7__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_u1y0n_L1_8 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_7__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_8__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_8__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_u1y0n_L1_9 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_8__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_9__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_9__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_u1y0n_L1_10 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_9__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_10__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_10__prog_data)
        );
    scanchain_data_d3 i_prog_data_i_sw_so_u1y0n_L1_11 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_10__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_so_u1y0n_L1_11__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_so_u1y0n_L1_11__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_so_u1y0n_L1_11__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign so_u1y0n_L1 = {_i_sw_so_u1y0n_L1_11__o,
        _i_sw_so_u1y0n_L1_10__o,
        _i_sw_so_u1y0n_L1_9__o,
        _i_sw_so_u1y0n_L1_8__o,
        _i_sw_so_u1y0n_L1_7__o,
        _i_sw_so_u1y0n_L1_6__o,
        _i_sw_so_u1y0n_L1_5__o,
        _i_sw_so_u1y0n_L1_4__o,
        _i_sw_so_u1y0n_L1_3__o,
        _i_sw_so_u1y0n_L1_2__o,
        _i_sw_so_u1y0n_L1_1__o,
        _i_sw_so_u1y0n_L1_0__o};
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_nw_w_ex_sw (
    input wire [11:0] bi_u1y0n_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    );
    
        
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
        
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
        

endmodule
// Automatically generated by PRGA's RTL generator
module sbox_sw_s_ex_sw (
    input wire [11:0] bi_u1v1e_L1
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    );
    
        
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
        
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
        

endmodule
// Automatically generated by PRGA's RTL generator
module prga_simple_buf (
    input wire [0:0] C,
    input wire [0:0] D,
    output reg [0:0] Q
    );

    always @(posedge C) begin
        Q <= D;
    end

endmodule// Automatically generated by PRGA's RTL generator
module prga_simple_bufr (
    input wire [0:0] C,
    input wire [0:0] R,
    input wire [0:0] D,
    output reg [0:0] Q
    );

    always @(posedge C) begin
        if (R) begin
            Q <= 1'b0;
        end else begin
            Q <= D;
        end
    end

endmodule// Automatically generated by PRGA's RTL generator
module iob (
    input wire [0:0] outpad
    , output wire [0:0] inpad
    , input wire [0:0] ipin
    , output wire [0:0] opin
    , output wire [0:0] oe
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _io__inpad;
    wire [0:0] _io__opin;
    wire [0:0] _io__oe;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_io__prog_dout;
    wire [1:0] _i_prog_data_io__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    iopad io (
        .outpad(outpad)
        ,.inpad(_io__inpad)
        ,.ipin(ipin)
        ,.opin(_io__opin)
        ,.oe(_io__oe)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_io__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d2 i_prog_data_io (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_io__prog_dout)
        ,.prog_data(_i_prog_data_io__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_io__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign inpad = _io__inpad;
    assign opin = _io__opin;
    assign oe = _io__oe;
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module cbox_t_io_w_e0 (
    output wire [0:0] bp_x0y0i0_outpad
    , input wire [11:0] bi_x0y0n_L1
    , input wire [11:0] bi_x0y0s_L1
    , input wire [0:0] bp_x0y0i0_inpad
    , output wire [11:0] cu_x0y0n_L1
    , output wire [11:0] cu_x0y0s_L1
    , output wire [0:0] bp_x0y0i1_outpad
    , input wire [0:0] bp_x0y0i1_inpad
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_bp_x0y0i0_outpad__o;
    wire [0:0] _i_sw_cu_x0y0n_L1_6__o;
    wire [0:0] _i_sw_cu_x0y0s_L1_6__o;
    wire [0:0] _i_sw_bp_x0y0i1_outpad__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_bp_x0y0i0_outpad__prog_dout;
    wire [3:0] _i_prog_data_i_sw_bp_x0y0i0_outpad__prog_data;
    wire [0:0] _i_prog_data_i_sw_cu_x0y0n_L1_6__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cu_x0y0n_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_cu_x0y0s_L1_6__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cu_x0y0s_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_bp_x0y0i1_outpad__prog_dout;
    wire [3:0] _i_prog_data_i_sw_bp_x0y0i1_outpad__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw12 i_sw_bp_x0y0i0_outpad (
        .i({bi_x0y0s_L1[10],
            bi_x0y0n_L1[10],
            bi_x0y0s_L1[8],
            bi_x0y0n_L1[8],
            bi_x0y0s_L1[6],
            bi_x0y0n_L1[6],
            bi_x0y0s_L1[4],
            bi_x0y0n_L1[4],
            bi_x0y0s_L1[2],
            bi_x0y0n_L1[2],
            bi_x0y0s_L1[0],
            bi_x0y0n_L1[0]})
        ,.o(_i_sw_bp_x0y0i0_outpad__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_outpad__prog_data)
        );
    sw2 i_sw_cu_x0y0n_L1_6 (
        .i({bp_x0y0i1_inpad,
            bp_x0y0i0_inpad})
        ,.o(_i_sw_cu_x0y0n_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cu_x0y0n_L1_6__prog_data)
        );
    sw2 i_sw_cu_x0y0s_L1_6 (
        .i({bp_x0y0i1_inpad,
            bp_x0y0i0_inpad})
        ,.o(_i_sw_cu_x0y0s_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cu_x0y0s_L1_6__prog_data)
        );
    sw12 i_sw_bp_x0y0i1_outpad (
        .i({bi_x0y0s_L1[11],
            bi_x0y0n_L1[11],
            bi_x0y0s_L1[9],
            bi_x0y0n_L1[9],
            bi_x0y0s_L1[7],
            bi_x0y0n_L1[7],
            bi_x0y0s_L1[6],
            bi_x0y0n_L1[6],
            bi_x0y0s_L1[3],
            bi_x0y0n_L1[3],
            bi_x0y0s_L1[1],
            bi_x0y0n_L1[1]})
        ,.o(_i_sw_bp_x0y0i1_outpad__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i1_outpad__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d4 i_prog_data_i_sw_bp_x0y0i0_outpad (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_bp_x0y0i0_outpad__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_outpad__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cu_x0y0n_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_bp_x0y0i0_outpad__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cu_x0y0n_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cu_x0y0n_L1_6__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cu_x0y0s_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cu_x0y0n_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cu_x0y0s_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cu_x0y0s_L1_6__prog_data)
        );
    scanchain_data_d4 i_prog_data_i_sw_bp_x0y0i1_outpad (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cu_x0y0s_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_bp_x0y0i1_outpad__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i1_outpad__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_bp_x0y0i1_outpad__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign bp_x0y0i0_outpad = _i_sw_bp_x0y0i0_outpad__o;
    assign cu_x0y0n_L1 = {bp_x0y0i1_inpad,
        bp_x0y0i0_inpad,
        bp_x0y0i1_inpad,
        bp_x0y0i0_inpad,
        bp_x0y0i1_inpad,
        _i_sw_cu_x0y0n_L1_6__o,
        1'bx,
        bp_x0y0i0_inpad,
        bp_x0y0i1_inpad,
        bp_x0y0i0_inpad,
        bp_x0y0i1_inpad,
        bp_x0y0i0_inpad};
    assign cu_x0y0s_L1 = {bp_x0y0i1_inpad,
        bp_x0y0i0_inpad,
        bp_x0y0i1_inpad,
        bp_x0y0i0_inpad,
        bp_x0y0i1_inpad,
        _i_sw_cu_x0y0s_L1_6__o,
        1'bx,
        bp_x0y0i0_inpad,
        bp_x0y0i1_inpad,
        bp_x0y0i0_inpad,
        bp_x0y0i1_inpad,
        bp_x0y0i0_inpad};
    assign bp_x0y0i1_outpad = _i_sw_bp_x0y0i1_outpad__o;
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module sw3 (
    input wire [2:0] i
    , output reg [0:0] o

    , input wire [0:0] prog_done
    , input wire [1:0] prog_data
    );

    always @* begin
        if (~prog_done) begin
            o = 1'b0;
        end else begin
            o = 1'b0;   // if ``prog_data == 0`` or ``prog_data`` out of bound, output 0
            case (prog_data)
                2'd1: o = i[0];
                2'd2: o = i[1];
                2'd3: o = i[2];
            endcase
        end
    end

endmodule// Automatically generated by PRGA's RTL generator
module sw2 (
    input wire [1:0] i
    , output reg [0:0] o

    , input wire [0:0] prog_done
    , input wire [1:0] prog_data
    );

    always @* begin
        if (~prog_done) begin
            o = 1'b0;
        end else begin
            o = 1'b0;   // if ``prog_data == 0`` or ``prog_data`` out of bound, output 0
            case (prog_data)
                2'd1: o = i[0];
                2'd2: o = i[1];
            endcase
        end
    end

endmodule// Automatically generated by PRGA's RTL generator
module scanchain_delim (
    input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done

    , input wire [0:0] prog_we
    , input wire [1 - 1:0] prog_din

    , output reg [0:0] prog_we_o
    , output reg [1 - 1:0] prog_dout
    );

    always @(posedge prog_clk) begin
        if (prog_rst) begin
            prog_we_o <= 1'b0;
            prog_dout <= 1'b0;
        end else if (~prog_done && prog_we) begin
            prog_we_o <= 1'b1;
            prog_dout <= prog_din;
        end else begin
            prog_we_o <= 1'b0;
        end
    end

endmodule// Automatically generated by PRGA's RTL generator
module scanchain_data_d2 (
    input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done

    , input wire [0:0] prog_we
    , input wire [1 - 1:0] prog_din

    , output reg [2 - 1:0] prog_data
    , output wire [1 - 1:0] prog_dout
    );

    localparam CHAIN_BITCOUNT = 2;
    localparam CHAIN_WIDTH = 1;

    wire [CHAIN_BITCOUNT + CHAIN_WIDTH - 1:0] prog_data_next;
    assign prog_data_next = {prog_data, prog_din};

    always @(posedge prog_clk) begin
        if (prog_rst) begin
            prog_data <= {CHAIN_BITCOUNT{1'b0}};
        end else if (~prog_done && prog_we) begin
            prog_data <= prog_data_next[0 +: CHAIN_BITCOUNT];
        end
    end

    assign prog_dout = prog_data_next[CHAIN_BITCOUNT +: CHAIN_WIDTH];

endmodule// Automatically generated by PRGA's RTL generator
module sw1 (
    input wire [0:0] i
    , output reg [0:0] o

    , input wire [0:0] prog_done
    , input wire [0:0] prog_data
    );

    always @* begin
        if (~prog_done) begin
            o = 1'b0;
        end else begin
            o = 1'b0;   // if ``prog_data == 0`` or ``prog_data`` out of bound, output 0
            case (prog_data)
                1'd1: o = i[0];
            endcase
        end
    end

endmodule// Automatically generated by PRGA's RTL generator
module scanchain_data_d1 (
    input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done

    , input wire [0:0] prog_we
    , input wire [1 - 1:0] prog_din

    , output reg [1 - 1:0] prog_data
    , output wire [1 - 1:0] prog_dout
    );

    localparam CHAIN_BITCOUNT = 1;
    localparam CHAIN_WIDTH = 1;

    wire [CHAIN_BITCOUNT + CHAIN_WIDTH - 1:0] prog_data_next;
    assign prog_data_next = {prog_data, prog_din};

    always @(posedge prog_clk) begin
        if (prog_rst) begin
            prog_data <= {CHAIN_BITCOUNT{1'b0}};
        end else if (~prog_done && prog_we) begin
            prog_data <= prog_data_next[0 +: CHAIN_BITCOUNT];
        end
    end

    assign prog_dout = prog_data_next[CHAIN_BITCOUNT +: CHAIN_WIDTH];

endmodule// Automatically generated by PRGA's RTL generator
module sw4 (
    input wire [3:0] i
    , output reg [0:0] o

    , input wire [0:0] prog_done
    , input wire [2:0] prog_data
    );

    always @* begin
        if (~prog_done) begin
            o = 1'b0;
        end else begin
            o = 1'b0;   // if ``prog_data == 0`` or ``prog_data`` out of bound, output 0
            case (prog_data)
                3'd1: o = i[0];
                3'd2: o = i[1];
                3'd3: o = i[2];
                3'd4: o = i[3];
            endcase
        end
    end

endmodule// Automatically generated by PRGA's RTL generator
module scanchain_data_d3 (
    input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done

    , input wire [0:0] prog_we
    , input wire [1 - 1:0] prog_din

    , output reg [3 - 1:0] prog_data
    , output wire [1 - 1:0] prog_dout
    );

    localparam CHAIN_BITCOUNT = 3;
    localparam CHAIN_WIDTH = 1;

    wire [CHAIN_BITCOUNT + CHAIN_WIDTH - 1:0] prog_data_next;
    assign prog_data_next = {prog_data, prog_din};

    always @(posedge prog_clk) begin
        if (prog_rst) begin
            prog_data <= {CHAIN_BITCOUNT{1'b0}};
        end else if (~prog_done && prog_we) begin
            prog_data <= prog_data_next[0 +: CHAIN_BITCOUNT];
        end
    end

    assign prog_dout = prog_data_next[CHAIN_BITCOUNT +: CHAIN_WIDTH];

endmodule// Automatically generated by PRGA's RTL generator
module cbox_t_io_n_s0 (
    output wire [0:0] bp_x0y0i0_outpad
    , input wire [11:0] bi_x0v1e_L1
    , input wire [11:0] bi_x0v1w_L1
    , input wire [0:0] bp_x0y0i0_inpad
    , output wire [11:0] cu_x0v1e_L1
    , output wire [11:0] cu_x0v1w_L1
    , output wire [0:0] bp_x0y0i1_outpad
    , input wire [0:0] bp_x0y0i1_inpad
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_bp_x0y0i0_outpad__o;
    wire [0:0] _i_sw_cu_x0v1e_L1_6__o;
    wire [0:0] _i_sw_cu_x0v1w_L1_6__o;
    wire [0:0] _i_sw_bp_x0y0i1_outpad__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_bp_x0y0i0_outpad__prog_dout;
    wire [3:0] _i_prog_data_i_sw_bp_x0y0i0_outpad__prog_data;
    wire [0:0] _i_prog_data_i_sw_cu_x0v1e_L1_6__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cu_x0v1e_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_cu_x0v1w_L1_6__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cu_x0v1w_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_bp_x0y0i1_outpad__prog_dout;
    wire [3:0] _i_prog_data_i_sw_bp_x0y0i1_outpad__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw12 i_sw_bp_x0y0i0_outpad (
        .i({bi_x0v1w_L1[10],
            bi_x0v1e_L1[10],
            bi_x0v1w_L1[8],
            bi_x0v1e_L1[8],
            bi_x0v1w_L1[6],
            bi_x0v1e_L1[6],
            bi_x0v1w_L1[4],
            bi_x0v1e_L1[4],
            bi_x0v1w_L1[2],
            bi_x0v1e_L1[2],
            bi_x0v1w_L1[0],
            bi_x0v1e_L1[0]})
        ,.o(_i_sw_bp_x0y0i0_outpad__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_outpad__prog_data)
        );
    sw2 i_sw_cu_x0v1e_L1_6 (
        .i({bp_x0y0i1_inpad,
            bp_x0y0i0_inpad})
        ,.o(_i_sw_cu_x0v1e_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cu_x0v1e_L1_6__prog_data)
        );
    sw2 i_sw_cu_x0v1w_L1_6 (
        .i({bp_x0y0i1_inpad,
            bp_x0y0i0_inpad})
        ,.o(_i_sw_cu_x0v1w_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cu_x0v1w_L1_6__prog_data)
        );
    sw12 i_sw_bp_x0y0i1_outpad (
        .i({bi_x0v1w_L1[11],
            bi_x0v1e_L1[11],
            bi_x0v1w_L1[9],
            bi_x0v1e_L1[9],
            bi_x0v1w_L1[7],
            bi_x0v1e_L1[7],
            bi_x0v1w_L1[6],
            bi_x0v1e_L1[6],
            bi_x0v1w_L1[3],
            bi_x0v1e_L1[3],
            bi_x0v1w_L1[1],
            bi_x0v1e_L1[1]})
        ,.o(_i_sw_bp_x0y0i1_outpad__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i1_outpad__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d4 i_prog_data_i_sw_bp_x0y0i0_outpad (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_bp_x0y0i0_outpad__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_outpad__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cu_x0v1e_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_bp_x0y0i0_outpad__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cu_x0v1e_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cu_x0v1e_L1_6__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cu_x0v1w_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cu_x0v1e_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cu_x0v1w_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cu_x0v1w_L1_6__prog_data)
        );
    scanchain_data_d4 i_prog_data_i_sw_bp_x0y0i1_outpad (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cu_x0v1w_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_bp_x0y0i1_outpad__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i1_outpad__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_bp_x0y0i1_outpad__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign bp_x0y0i0_outpad = _i_sw_bp_x0y0i0_outpad__o;
    assign cu_x0v1e_L1 = {bp_x0y0i1_inpad,
        bp_x0y0i0_inpad,
        bp_x0y0i1_inpad,
        bp_x0y0i0_inpad,
        bp_x0y0i1_inpad,
        _i_sw_cu_x0v1e_L1_6__o,
        1'bx,
        bp_x0y0i0_inpad,
        bp_x0y0i1_inpad,
        bp_x0y0i0_inpad,
        bp_x0y0i1_inpad,
        bp_x0y0i0_inpad};
    assign cu_x0v1w_L1 = {bp_x0y0i1_inpad,
        bp_x0y0i0_inpad,
        bp_x0y0i1_inpad,
        bp_x0y0i0_inpad,
        bp_x0y0i1_inpad,
        _i_sw_cu_x0v1w_L1_6__o,
        1'bx,
        bp_x0y0i0_inpad,
        bp_x0y0i1_inpad,
        bp_x0y0i0_inpad,
        bp_x0y0i1_inpad,
        bp_x0y0i0_inpad};
    assign bp_x0y0i1_outpad = _i_sw_bp_x0y0i1_outpad__o;
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module cbox_t_io_e_w0 (
    output wire [0:0] bp_x0y0i0_outpad
    , input wire [11:0] bi_u1y0n_L1
    , input wire [11:0] bi_u1y0s_L1
    , input wire [0:0] bp_x0y0i0_inpad
    , output wire [11:0] cu_u1y0n_L1
    , output wire [11:0] cu_u1y0s_L1
    , output wire [0:0] bp_x0y0i1_outpad
    , input wire [0:0] bp_x0y0i1_inpad
    , input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done
    , input wire [0:0] prog_we
    , input wire [0:0] prog_din
    , output wire [0:0] prog_dout
    , output wire [0:0] prog_we_o
    );
    
        
    wire [0:0] _i_sw_bp_x0y0i0_outpad__o;
    wire [0:0] _i_sw_cu_u1y0n_L1_6__o;
    wire [0:0] _i_sw_cu_u1y0s_L1_6__o;
    wire [0:0] _i_sw_bp_x0y0i1_outpad__o;
    wire [0:0] _i_buf_prog_rst_l0__Q;
    wire [0:0] _i_buf_prog_done_l0__Q;
    wire [0:0] _i_scanchain_head__prog_dout;
    wire [0:0] _i_scanchain_head__prog_we_o;
    wire [0:0] _i_prog_data_i_sw_bp_x0y0i0_outpad__prog_dout;
    wire [3:0] _i_prog_data_i_sw_bp_x0y0i0_outpad__prog_data;
    wire [0:0] _i_prog_data_i_sw_cu_u1y0n_L1_6__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cu_u1y0n_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_cu_u1y0s_L1_6__prog_dout;
    wire [1:0] _i_prog_data_i_sw_cu_u1y0s_L1_6__prog_data;
    wire [0:0] _i_prog_data_i_sw_bp_x0y0i1_outpad__prog_dout;
    wire [3:0] _i_prog_data_i_sw_bp_x0y0i1_outpad__prog_data;
    wire [0:0] _i_scanchain_tail__prog_dout;
    wire [0:0] _i_scanchain_tail__prog_we_o;
        
    sw12 i_sw_bp_x0y0i0_outpad (
        .i({bi_u1y0s_L1[10],
            bi_u1y0n_L1[10],
            bi_u1y0s_L1[8],
            bi_u1y0n_L1[8],
            bi_u1y0s_L1[6],
            bi_u1y0n_L1[6],
            bi_u1y0s_L1[4],
            bi_u1y0n_L1[4],
            bi_u1y0s_L1[2],
            bi_u1y0n_L1[2],
            bi_u1y0s_L1[0],
            bi_u1y0n_L1[0]})
        ,.o(_i_sw_bp_x0y0i0_outpad__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_outpad__prog_data)
        );
    sw2 i_sw_cu_u1y0n_L1_6 (
        .i({bp_x0y0i1_inpad,
            bp_x0y0i0_inpad})
        ,.o(_i_sw_cu_u1y0n_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cu_u1y0n_L1_6__prog_data)
        );
    sw2 i_sw_cu_u1y0s_L1_6 (
        .i({bp_x0y0i1_inpad,
            bp_x0y0i0_inpad})
        ,.o(_i_sw_cu_u1y0s_L1_6__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_cu_u1y0s_L1_6__prog_data)
        );
    sw12 i_sw_bp_x0y0i1_outpad (
        .i({bi_u1y0s_L1[11],
            bi_u1y0n_L1[11],
            bi_u1y0s_L1[9],
            bi_u1y0n_L1[9],
            bi_u1y0s_L1[7],
            bi_u1y0n_L1[7],
            bi_u1y0s_L1[6],
            bi_u1y0n_L1[6],
            bi_u1y0s_L1[3],
            bi_u1y0n_L1[3],
            bi_u1y0s_L1[1],
            bi_u1y0n_L1[1]})
        ,.o(_i_sw_bp_x0y0i1_outpad__o)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i1_outpad__prog_data)
        );
    prga_simple_buf i_buf_prog_rst_l0 (
        .C(prog_clk)
        ,.D(prog_rst)
        ,.Q(_i_buf_prog_rst_l0__Q)
        );
    prga_simple_bufr i_buf_prog_done_l0 (
        .C(prog_clk)
        ,.R(_i_buf_prog_rst_l0__Q)
        ,.D(prog_done)
        ,.Q(_i_buf_prog_done_l0__Q)
        );
    scanchain_delim i_scanchain_head (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(prog_we)
        ,.prog_din(prog_din)
        ,.prog_dout(_i_scanchain_head__prog_dout)
        ,.prog_we_o(_i_scanchain_head__prog_we_o)
        );
    scanchain_data_d4 i_prog_data_i_sw_bp_x0y0i0_outpad (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_scanchain_head__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_bp_x0y0i0_outpad__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i0_outpad__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cu_u1y0n_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_bp_x0y0i0_outpad__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cu_u1y0n_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cu_u1y0n_L1_6__prog_data)
        );
    scanchain_data_d2 i_prog_data_i_sw_cu_u1y0s_L1_6 (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cu_u1y0n_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_cu_u1y0s_L1_6__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_cu_u1y0s_L1_6__prog_data)
        );
    scanchain_data_d4 i_prog_data_i_sw_bp_x0y0i1_outpad (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_cu_u1y0s_L1_6__prog_dout)
        ,.prog_dout(_i_prog_data_i_sw_bp_x0y0i1_outpad__prog_dout)
        ,.prog_data(_i_prog_data_i_sw_bp_x0y0i1_outpad__prog_data)
        );
    scanchain_delim i_scanchain_tail (
        .prog_clk(prog_clk)
        ,.prog_rst(_i_buf_prog_rst_l0__Q)
        ,.prog_done(_i_buf_prog_done_l0__Q)
        ,.prog_we(_i_scanchain_head__prog_we_o)
        ,.prog_din(_i_prog_data_i_sw_bp_x0y0i1_outpad__prog_dout)
        ,.prog_dout(_i_scanchain_tail__prog_dout)
        ,.prog_we_o(_i_scanchain_tail__prog_we_o)
        );
        
    assign bp_x0y0i0_outpad = _i_sw_bp_x0y0i0_outpad__o;
    assign cu_u1y0n_L1 = {bp_x0y0i1_inpad,
        bp_x0y0i0_inpad,
        bp_x0y0i1_inpad,
        bp_x0y0i0_inpad,
        bp_x0y0i1_inpad,
        _i_sw_cu_u1y0n_L1_6__o,
        1'bx,
        bp_x0y0i0_inpad,
        bp_x0y0i1_inpad,
        bp_x0y0i0_inpad,
        bp_x0y0i1_inpad,
        bp_x0y0i0_inpad};
    assign cu_u1y0s_L1 = {bp_x0y0i1_inpad,
        bp_x0y0i0_inpad,
        bp_x0y0i1_inpad,
        bp_x0y0i0_inpad,
        bp_x0y0i1_inpad,
        _i_sw_cu_u1y0s_L1_6__o,
        1'bx,
        bp_x0y0i0_inpad,
        bp_x0y0i1_inpad,
        bp_x0y0i0_inpad,
        bp_x0y0i1_inpad,
        bp_x0y0i0_inpad};
    assign bp_x0y0i1_outpad = _i_sw_bp_x0y0i1_outpad__o;
    assign prog_dout = _i_scanchain_tail__prog_dout;
    assign prog_we_o = _i_scanchain_tail__prog_we_o;

endmodule
// Automatically generated by PRGA's RTL generator
module iopad (
    input wire [0:0] outpad
    , output reg [0:0] inpad

    , input wire [0:0] ipin
    , output reg [0:0] opin
    , output reg [0:0] oe

    , input wire [0:0] prog_done    // programming
    , input wire [1:0] prog_data    // mode:
                                    //  - 00: disabled
                                    //  - 01: input mode
                                    //  - 10: output mode
    );

    localparam  MODE_INPUT      = 2'h1,
                MODE_OUTPUT     = 2'h2;

    always @* begin
        inpad = 1'b0;
        opin = 1'b0;
        oe = 1'b0;

        if (prog_done) begin
            case (prog_data)
                MODE_INPUT: begin
                    inpad = ipin;
                end
                MODE_OUTPUT: begin
                    opin = outpad;
                    oe = 1'b1;
                end
            endcase
        end
    end

endmodule// Automatically generated by PRGA's RTL generator
module sw12 (
    input wire [11:0] i
    , output reg [0:0] o

    , input wire [0:0] prog_done
    , input wire [3:0] prog_data
    );

    always @* begin
        if (~prog_done) begin
            o = 1'b0;
        end else begin
            o = 1'b0;   // if ``prog_data == 0`` or ``prog_data`` out of bound, output 0
            case (prog_data)
                4'd1: o = i[0];
                4'd2: o = i[1];
                4'd3: o = i[2];
                4'd4: o = i[3];
                4'd5: o = i[4];
                4'd6: o = i[5];
                4'd7: o = i[6];
                4'd8: o = i[7];
                4'd9: o = i[8];
                4'd10: o = i[9];
                4'd11: o = i[10];
                4'd12: o = i[11];
            endcase
        end
    end

endmodule// Automatically generated by PRGA's RTL generator
module scanchain_data_d4 (
    input wire [0:0] prog_clk
    , input wire [0:0] prog_rst
    , input wire [0:0] prog_done

    , input wire [0:0] prog_we
    , input wire [1 - 1:0] prog_din

    , output reg [4 - 1:0] prog_data
    , output wire [1 - 1:0] prog_dout
    );

    localparam CHAIN_BITCOUNT = 4;
    localparam CHAIN_WIDTH = 1;

    wire [CHAIN_BITCOUNT + CHAIN_WIDTH - 1:0] prog_data_next;
    assign prog_data_next = {prog_data, prog_din};

    always @(posedge prog_clk) begin
        if (prog_rst) begin
            prog_data <= {CHAIN_BITCOUNT{1'b0}};
        end else if (~prog_done && prog_we) begin
            prog_data <= prog_data_next[0 +: CHAIN_BITCOUNT];
        end
    end

    assign prog_dout = prog_data_next[CHAIN_BITCOUNT +: CHAIN_WIDTH];

endmodule
