VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tile_clb
  CLASS BLOCK ;
  FOREIGN tile_clb ;
  ORIGIN 0.000 0.000 ;
  SIZE 165.600 BY 244.800 ;
  PIN bi_u1y0n_L1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 5.130 4.000 5.410 ;
    END
  END bi_u1y0n_L1[0]
  PIN bi_u1y0n_L1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 209.130 4.000 209.410 ;
    END
  END bi_u1y0n_L1[10]
  PIN bi_u1y0n_L1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 229.530 4.000 229.810 ;
    END
  END bi_u1y0n_L1[11]
  PIN bi_u1y0n_L1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 25.530 4.000 25.810 ;
    END
  END bi_u1y0n_L1[1]
  PIN bi_u1y0n_L1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 45.930 4.000 46.210 ;
    END
  END bi_u1y0n_L1[2]
  PIN bi_u1y0n_L1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 66.330 4.000 66.610 ;
    END
  END bi_u1y0n_L1[3]
  PIN bi_u1y0n_L1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 86.730 4.000 87.010 ;
    END
  END bi_u1y0n_L1[4]
  PIN bi_u1y0n_L1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 107.130 4.000 107.410 ;
    END
  END bi_u1y0n_L1[5]
  PIN bi_u1y0n_L1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 127.530 4.000 127.810 ;
    END
  END bi_u1y0n_L1[6]
  PIN bi_u1y0n_L1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 147.930 4.000 148.210 ;
    END
  END bi_u1y0n_L1[7]
  PIN bi_u1y0n_L1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 168.330 4.000 168.610 ;
    END
  END bi_u1y0n_L1[8]
  PIN bi_u1y0n_L1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 188.730 4.000 189.010 ;
    END
  END bi_u1y0n_L1[9]
  PIN bi_u1y0s_L1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 15.330 4.000 15.610 ;
    END
  END bi_u1y0s_L1[0]
  PIN bi_u1y0s_L1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 219.330 4.000 219.610 ;
    END
  END bi_u1y0s_L1[10]
  PIN bi_u1y0s_L1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 239.730 4.000 240.010 ;
    END
  END bi_u1y0s_L1[11]
  PIN bi_u1y0s_L1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 35.730 4.000 36.010 ;
    END
  END bi_u1y0s_L1[1]
  PIN bi_u1y0s_L1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 56.130 4.000 56.410 ;
    END
  END bi_u1y0s_L1[2]
  PIN bi_u1y0s_L1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 76.530 4.000 76.810 ;
    END
  END bi_u1y0s_L1[3]
  PIN bi_u1y0s_L1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 96.930 4.000 97.210 ;
    END
  END bi_u1y0s_L1[4]
  PIN bi_u1y0s_L1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 117.330 4.000 117.610 ;
    END
  END bi_u1y0s_L1[5]
  PIN bi_u1y0s_L1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 137.730 4.000 138.010 ;
    END
  END bi_u1y0s_L1[6]
  PIN bi_u1y0s_L1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 158.130 4.000 158.410 ;
    END
  END bi_u1y0s_L1[7]
  PIN bi_u1y0s_L1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 178.530 4.000 178.810 ;
    END
  END bi_u1y0s_L1[8]
  PIN bi_u1y0s_L1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000 198.930 4.000 199.210 ;
    END
  END bi_u1y0s_L1[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END clk
  PIN cu_x0y0n_L1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.600 5.130 165.600 5.410 ;
    END
  END cu_x0y0n_L1[0]
  PIN cu_x0y0n_L1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.600 209.130 165.600 209.410 ;
    END
  END cu_x0y0n_L1[10]
  PIN cu_x0y0n_L1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.600 229.530 165.600 229.810 ;
    END
  END cu_x0y0n_L1[11]
  PIN cu_x0y0n_L1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.600 25.530 165.600 25.810 ;
    END
  END cu_x0y0n_L1[1]
  PIN cu_x0y0n_L1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.600 45.930 165.600 46.210 ;
    END
  END cu_x0y0n_L1[2]
  PIN cu_x0y0n_L1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.600 66.330 165.600 66.610 ;
    END
  END cu_x0y0n_L1[3]
  PIN cu_x0y0n_L1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.600 86.730 165.600 87.010 ;
    END
  END cu_x0y0n_L1[4]
  PIN cu_x0y0n_L1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.600 107.130 165.600 107.410 ;
    END
  END cu_x0y0n_L1[5]
  PIN cu_x0y0n_L1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.600 127.530 165.600 127.810 ;
    END
  END cu_x0y0n_L1[6]
  PIN cu_x0y0n_L1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.600 147.930 165.600 148.210 ;
    END
  END cu_x0y0n_L1[7]
  PIN cu_x0y0n_L1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.600 168.330 165.600 168.610 ;
    END
  END cu_x0y0n_L1[8]
  PIN cu_x0y0n_L1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.600 188.730 165.600 189.010 ;
    END
  END cu_x0y0n_L1[9]
  PIN cu_x0y0s_L1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.600 15.330 165.600 15.610 ;
    END
  END cu_x0y0s_L1[0]
  PIN cu_x0y0s_L1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.600 219.330 165.600 219.610 ;
    END
  END cu_x0y0s_L1[10]
  PIN cu_x0y0s_L1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.600 239.730 165.600 240.010 ;
    END
  END cu_x0y0s_L1[11]
  PIN cu_x0y0s_L1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.600 35.730 165.600 36.010 ;
    END
  END cu_x0y0s_L1[1]
  PIN cu_x0y0s_L1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.600 56.130 165.600 56.410 ;
    END
  END cu_x0y0s_L1[2]
  PIN cu_x0y0s_L1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.600 76.530 165.600 76.810 ;
    END
  END cu_x0y0s_L1[3]
  PIN cu_x0y0s_L1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.600 96.930 165.600 97.210 ;
    END
  END cu_x0y0s_L1[4]
  PIN cu_x0y0s_L1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.600 117.330 165.600 117.610 ;
    END
  END cu_x0y0s_L1[5]
  PIN cu_x0y0s_L1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.600 137.730 165.600 138.010 ;
    END
  END cu_x0y0s_L1[6]
  PIN cu_x0y0s_L1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.600 158.130 165.600 158.410 ;
    END
  END cu_x0y0s_L1[7]
  PIN cu_x0y0s_L1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.600 178.530 165.600 178.810 ;
    END
  END cu_x0y0s_L1[8]
  PIN cu_x0y0s_L1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 161.600 198.930 165.600 199.210 ;
    END
  END cu_x0y0s_L1[9]
  PIN prog_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END prog_clk
  PIN prog_din
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END prog_din
  PIN prog_done
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END prog_done
  PIN prog_dout
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 240.800 41.770 244.800 ;
    END
  END prog_dout
  PIN prog_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END prog_rst
  PIN prog_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END prog_we
  PIN prog_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 240.800 124.570 244.800 ;
    END
  END prog_we_o
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 5.520 7.960 160.080 8.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520 73.240 160.080 73.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520 138.520 160.080 139.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520 203.800 160.080 204.400 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 5.520 40.600 160.080 41.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520 105.880 160.080 106.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520 171.160 160.080 171.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.520 236.440 160.080 237.040 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 2.635 160.080 242.165 ;
      LAYER met1 ;
        RECT 3.840 240.290 161.760 242.320 ;
        RECT 4.280 239.450 161.320 240.290 ;
        RECT 3.840 230.090 161.760 239.450 ;
        RECT 4.280 229.250 161.320 230.090 ;
        RECT 3.840 219.890 161.760 229.250 ;
        RECT 4.280 219.050 161.320 219.890 ;
        RECT 3.840 209.690 161.760 219.050 ;
        RECT 4.280 208.850 161.320 209.690 ;
        RECT 3.840 199.490 161.760 208.850 ;
        RECT 4.280 198.650 161.320 199.490 ;
        RECT 3.840 189.290 161.760 198.650 ;
        RECT 4.280 188.450 161.320 189.290 ;
        RECT 3.840 179.090 161.760 188.450 ;
        RECT 4.280 178.250 161.320 179.090 ;
        RECT 3.840 168.890 161.760 178.250 ;
        RECT 4.280 168.050 161.320 168.890 ;
        RECT 3.840 158.690 161.760 168.050 ;
        RECT 4.280 157.850 161.320 158.690 ;
        RECT 3.840 148.490 161.760 157.850 ;
        RECT 4.280 147.650 161.320 148.490 ;
        RECT 3.840 138.290 161.760 147.650 ;
        RECT 4.280 137.450 161.320 138.290 ;
        RECT 3.840 128.090 161.760 137.450 ;
        RECT 4.280 127.250 161.320 128.090 ;
        RECT 3.840 117.890 161.760 127.250 ;
        RECT 4.280 117.050 161.320 117.890 ;
        RECT 3.840 107.690 161.760 117.050 ;
        RECT 4.280 106.850 161.320 107.690 ;
        RECT 3.840 97.490 161.760 106.850 ;
        RECT 4.280 96.650 161.320 97.490 ;
        RECT 3.840 87.290 161.760 96.650 ;
        RECT 4.280 86.450 161.320 87.290 ;
        RECT 3.840 77.090 161.760 86.450 ;
        RECT 4.280 76.250 161.320 77.090 ;
        RECT 3.840 66.890 161.760 76.250 ;
        RECT 4.280 66.050 161.320 66.890 ;
        RECT 3.840 56.690 161.760 66.050 ;
        RECT 4.280 55.850 161.320 56.690 ;
        RECT 3.840 46.490 161.760 55.850 ;
        RECT 4.280 45.650 161.320 46.490 ;
        RECT 3.840 36.290 161.760 45.650 ;
        RECT 4.280 35.450 161.320 36.290 ;
        RECT 3.840 26.090 161.760 35.450 ;
        RECT 4.280 25.250 161.320 26.090 ;
        RECT 3.840 15.890 161.760 25.250 ;
        RECT 4.280 15.050 161.320 15.890 ;
        RECT 3.840 5.690 161.760 15.050 ;
        RECT 4.280 4.850 161.320 5.690 ;
        RECT 3.840 2.080 161.760 4.850 ;
      LAYER met2 ;
        RECT 6.080 240.520 41.210 242.320 ;
        RECT 42.050 240.520 124.010 242.320 ;
        RECT 124.850 240.520 158.600 242.320 ;
        RECT 6.080 4.280 158.600 240.520 ;
        RECT 6.080 2.050 13.610 4.280 ;
        RECT 14.450 2.050 41.210 4.280 ;
        RECT 42.050 2.050 68.810 4.280 ;
        RECT 69.650 2.050 96.410 4.280 ;
        RECT 97.250 2.050 124.010 4.280 ;
        RECT 124.850 2.050 151.610 4.280 ;
        RECT 152.450 2.050 158.600 4.280 ;
  END
END tile_clb
END LIBRARY

