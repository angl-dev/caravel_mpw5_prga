magic
tech sky130A
magscale 1 2
timestamp 1647871756
<< metal1 >>
rect 71774 702992 71780 703044
rect 71832 703032 71838 703044
rect 72970 703032 72976 703044
rect 71832 703004 72976 703032
rect 71832 702992 71838 703004
rect 72970 702992 72976 703004
rect 73028 702992 73034 703044
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 13722 700816 13728 700868
rect 13780 700856 13786 700868
rect 24302 700856 24308 700868
rect 13780 700828 24308 700856
rect 13780 700816 13786 700828
rect 24302 700816 24308 700828
rect 24360 700816 24366 700868
rect 13630 700748 13636 700800
rect 13688 700788 13694 700800
rect 89162 700788 89168 700800
rect 13688 700760 89168 700788
rect 13688 700748 13694 700760
rect 89162 700748 89168 700760
rect 89220 700748 89226 700800
rect 13078 700680 13084 700732
rect 13136 700720 13142 700732
rect 137830 700720 137836 700732
rect 13136 700692 137836 700720
rect 13136 700680 13142 700692
rect 137830 700680 137836 700692
rect 137888 700680 137894 700732
rect 365714 700680 365720 700732
rect 365772 700720 365778 700732
rect 462314 700720 462320 700732
rect 365772 700692 462320 700720
rect 365772 700680 365778 700692
rect 462314 700680 462320 700692
rect 462372 700680 462378 700732
rect 13446 700612 13452 700664
rect 13504 700652 13510 700664
rect 218974 700652 218980 700664
rect 13504 700624 218980 700652
rect 13504 700612 13510 700624
rect 218974 700612 218980 700624
rect 219032 700612 219038 700664
rect 376754 700612 376760 700664
rect 376812 700652 376818 700664
rect 527174 700652 527180 700664
rect 376812 700624 527180 700652
rect 376812 700612 376818 700624
rect 527174 700612 527180 700624
rect 527232 700612 527238 700664
rect 13354 700544 13360 700596
rect 13412 700584 13418 700596
rect 283834 700584 283840 700596
rect 13412 700556 283840 700584
rect 13412 700544 13418 700556
rect 283834 700544 283840 700556
rect 283892 700544 283898 700596
rect 330478 700544 330484 700596
rect 330536 700584 330542 700596
rect 494790 700584 494796 700596
rect 330536 700556 494796 700584
rect 330536 700544 330542 700556
rect 494790 700544 494796 700556
rect 494848 700544 494854 700596
rect 13538 700476 13544 700528
rect 13596 700516 13602 700528
rect 154114 700516 154120 700528
rect 13596 700488 154120 700516
rect 13596 700476 13602 700488
rect 154114 700476 154120 700488
rect 154172 700476 154178 700528
rect 193214 700476 193220 700528
rect 193272 700516 193278 700528
rect 478506 700516 478512 700528
rect 193272 700488 478512 700516
rect 193272 700476 193278 700488
rect 478506 700476 478512 700488
rect 478564 700476 478570 700528
rect 13262 700408 13268 700460
rect 13320 700448 13326 700460
rect 348786 700448 348792 700460
rect 13320 700420 348792 700448
rect 13320 700408 13326 700420
rect 348786 700408 348792 700420
rect 348844 700408 348850 700460
rect 398098 700408 398104 700460
rect 398156 700448 398162 700460
rect 559650 700448 559656 700460
rect 398156 700420 559656 700448
rect 398156 700408 398162 700420
rect 559650 700408 559656 700420
rect 559708 700408 559714 700460
rect 12986 700340 12992 700392
rect 13044 700380 13050 700392
rect 202782 700380 202788 700392
rect 13044 700352 202788 700380
rect 13044 700340 13050 700352
rect 202782 700340 202788 700352
rect 202840 700340 202846 700392
rect 204254 700340 204260 700392
rect 204312 700380 204318 700392
rect 543458 700380 543464 700392
rect 204312 700352 543464 700380
rect 204312 700340 204318 700352
rect 543458 700340 543464 700352
rect 543516 700340 543522 700392
rect 21358 700272 21364 700324
rect 21416 700312 21422 700324
rect 413646 700312 413652 700324
rect 21416 700284 413652 700312
rect 21416 700272 21422 700284
rect 413646 700272 413652 700284
rect 413704 700272 413710 700324
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 387794 696940 387800 696992
rect 387852 696980 387858 696992
rect 580166 696980 580172 696992
rect 387852 696952 580172 696980
rect 387852 696940 387858 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 2774 683680 2780 683732
rect 2832 683720 2838 683732
rect 4798 683720 4804 683732
rect 2832 683692 4804 683720
rect 2832 683680 2838 683692
rect 4798 683680 4804 683692
rect 4856 683680 4862 683732
rect 215294 683136 215300 683188
rect 215352 683176 215358 683188
rect 580166 683176 580172 683188
rect 215352 683148 580172 683176
rect 215352 683136 215358 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 11790 670732 11796 670744
rect 3568 670704 11796 670732
rect 3568 670692 3574 670704
rect 11790 670692 11796 670704
rect 11848 670692 11854 670744
rect 41506 670692 41512 670744
rect 41564 670732 41570 670744
rect 580166 670732 580172 670744
rect 41564 670704 580172 670732
rect 41564 670692 41570 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 14274 659064 14280 659116
rect 14332 659104 14338 659116
rect 266354 659104 266360 659116
rect 14332 659076 266360 659104
rect 14332 659064 14338 659076
rect 266354 659064 266360 659076
rect 266412 659064 266418 659116
rect 14366 658996 14372 659048
rect 14424 659036 14430 659048
rect 331214 659036 331220 659048
rect 14424 659008 331220 659036
rect 14424 658996 14430 659008
rect 331214 658996 331220 659008
rect 331272 658996 331278 659048
rect 14458 658928 14464 658980
rect 14516 658968 14522 658980
rect 397454 658968 397460 658980
rect 14516 658940 397460 658968
rect 14516 658928 14522 658940
rect 397454 658928 397460 658940
rect 397512 658928 397518 658980
rect 442902 657772 442908 657824
rect 442960 657812 442966 657824
rect 536558 657812 536564 657824
rect 442960 657784 536564 657812
rect 442960 657772 442966 657784
rect 536558 657772 536564 657784
rect 536616 657772 536622 657824
rect 13998 657704 14004 657756
rect 14056 657744 14062 657756
rect 169754 657744 169760 657756
rect 14056 657716 169760 657744
rect 14056 657704 14062 657716
rect 169754 657704 169760 657716
rect 169812 657704 169818 657756
rect 237282 657704 237288 657756
rect 237340 657744 237346 657756
rect 464982 657744 464988 657756
rect 237340 657716 464988 657744
rect 237340 657704 237346 657716
rect 464982 657704 464988 657716
rect 465040 657704 465046 657756
rect 486418 657704 486424 657756
rect 486476 657744 486482 657756
rect 539226 657744 539232 657756
rect 486476 657716 539232 657744
rect 486476 657704 486482 657716
rect 539226 657704 539232 657716
rect 539284 657704 539290 657756
rect 14182 657636 14188 657688
rect 14240 657676 14246 657688
rect 299474 657676 299480 657688
rect 14240 657648 299480 657676
rect 14240 657636 14246 657648
rect 299474 657636 299480 657648
rect 299532 657636 299538 657688
rect 475562 657636 475568 657688
rect 475620 657676 475626 657688
rect 536282 657676 536288 657688
rect 475620 657648 536288 657676
rect 475620 657636 475626 657648
rect 536282 657636 536288 657648
rect 536340 657636 536346 657688
rect 20622 657568 20628 657620
rect 20680 657608 20686 657620
rect 330478 657608 330484 657620
rect 20680 657580 330484 657608
rect 20680 657568 20686 657580
rect 330478 657568 330484 657580
rect 330536 657568 330542 657620
rect 421466 657568 421472 657620
rect 421524 657608 421530 657620
rect 492582 657608 492588 657620
rect 421524 657580 492588 657608
rect 421524 657568 421530 657580
rect 492582 657568 492588 657580
rect 492640 657568 492646 657620
rect 497274 657568 497280 657620
rect 497332 657608 497338 657620
rect 539134 657608 539140 657620
rect 497332 657580 539140 657608
rect 497332 657568 497338 657580
rect 539134 657568 539140 657580
rect 539192 657568 539198 657620
rect 31386 657500 31392 657552
rect 31444 657540 31450 657552
rect 398098 657540 398104 657552
rect 31444 657512 398104 657540
rect 31444 657500 31450 657512
rect 398098 657500 398104 657512
rect 398156 657500 398162 657552
rect 453850 657500 453856 657552
rect 453908 657540 453914 657552
rect 534994 657540 535000 657552
rect 453908 657512 535000 657540
rect 453908 657500 453914 657512
rect 534994 657500 535000 657512
rect 535052 657500 535058 657552
rect 464706 657432 464712 657484
rect 464764 657472 464770 657484
rect 536466 657472 536472 657484
rect 464764 657444 536472 657472
rect 464764 657432 464770 657444
rect 536466 657432 536472 657444
rect 536524 657432 536530 657484
rect 302142 657364 302148 657416
rect 302200 657404 302206 657416
rect 536190 657404 536196 657416
rect 302200 657376 536196 657404
rect 302200 657364 302206 657376
rect 536190 657364 536196 657376
rect 536248 657364 536254 657416
rect 291010 657296 291016 657348
rect 291068 657336 291074 657348
rect 536374 657336 536380 657348
rect 291068 657308 536380 657336
rect 291068 657296 291074 657308
rect 536374 657296 536380 657308
rect 536432 657296 536438 657348
rect 118050 657228 118056 657280
rect 118108 657268 118114 657280
rect 365622 657268 365628 657280
rect 118108 657240 365628 657268
rect 118108 657228 118114 657240
rect 365622 657228 365628 657240
rect 365680 657228 365686 657280
rect 399754 657228 399760 657280
rect 399812 657268 399818 657280
rect 535270 657268 535276 657280
rect 399812 657240 535276 657268
rect 399812 657228 399818 657240
rect 535270 657228 535276 657240
rect 535328 657228 535334 657280
rect 280706 657160 280712 657212
rect 280764 657200 280770 657212
rect 540238 657200 540244 657212
rect 280764 657172 540244 657200
rect 280764 657160 280770 657172
rect 540238 657160 540244 657172
rect 540296 657160 540302 657212
rect 269850 657092 269856 657144
rect 269908 657132 269914 657144
rect 540330 657132 540336 657144
rect 269908 657104 540336 657132
rect 269908 657092 269914 657104
rect 540330 657092 540336 657104
rect 540388 657092 540394 657144
rect 248046 657024 248052 657076
rect 248104 657064 248110 657076
rect 540422 657064 540428 657076
rect 248104 657036 540428 657064
rect 248104 657024 248110 657036
rect 540422 657024 540428 657036
rect 540480 657024 540486 657076
rect 128906 656956 128912 657008
rect 128964 656996 128970 657008
rect 430574 656996 430580 657008
rect 128964 656968 430580 656996
rect 128964 656956 128970 656968
rect 430574 656956 430580 656968
rect 430632 656956 430638 657008
rect 432322 656956 432328 657008
rect 432380 656996 432386 657008
rect 535086 656996 535092 657008
rect 432380 656968 535092 656996
rect 432380 656956 432386 656968
rect 535086 656956 535092 656968
rect 535144 656956 535150 657008
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 11882 656928 11888 656940
rect 3476 656900 11888 656928
rect 3476 656888 3482 656900
rect 11882 656888 11888 656900
rect 11940 656888 11946 656940
rect 96522 656888 96528 656940
rect 96580 656928 96586 656940
rect 453942 656928 453948 656940
rect 96580 656900 453948 656928
rect 96580 656888 96586 656900
rect 453942 656888 453948 656900
rect 454000 656888 454006 656940
rect 529842 656888 529848 656940
rect 529900 656928 529906 656940
rect 534718 656928 534724 656940
rect 529900 656900 534724 656928
rect 529900 656888 529906 656900
rect 534718 656888 534724 656900
rect 534776 656888 534782 656940
rect 13170 656276 13176 656328
rect 13228 656316 13234 656328
rect 21358 656316 21364 656328
rect 13228 656288 21364 656316
rect 13228 656276 13234 656288
rect 21358 656276 21364 656288
rect 21416 656276 21422 656328
rect 453942 656276 453948 656328
rect 454000 656316 454006 656328
rect 580810 656316 580816 656328
rect 454000 656288 580816 656316
rect 454000 656276 454006 656288
rect 580810 656276 580816 656288
rect 580868 656276 580874 656328
rect 12894 656208 12900 656260
rect 12952 656248 12958 656260
rect 71774 656248 71780 656260
rect 12952 656220 71780 656248
rect 12952 656208 12958 656220
rect 71774 656208 71780 656220
rect 71832 656208 71838 656260
rect 430574 656208 430580 656260
rect 430632 656248 430638 656260
rect 580534 656248 580540 656260
rect 430632 656220 580540 656248
rect 430632 656208 430638 656220
rect 580534 656208 580540 656220
rect 580592 656208 580598 656260
rect 14090 656140 14096 656192
rect 14148 656180 14154 656192
rect 234614 656180 234620 656192
rect 14148 656152 234620 656180
rect 14148 656140 14154 656152
rect 234614 656140 234620 656152
rect 234672 656140 234678 656192
rect 365622 656140 365628 656192
rect 365680 656180 365686 656192
rect 580718 656180 580724 656192
rect 365680 656152 580724 656180
rect 365680 656140 365686 656152
rect 580718 656140 580724 656152
rect 580776 656140 580782 656192
rect 507670 656072 507676 656124
rect 507728 656112 507734 656124
rect 534902 656112 534908 656124
rect 507728 656084 534908 656112
rect 507728 656072 507734 656084
rect 534902 656072 534908 656084
rect 534960 656072 534966 656124
rect 183186 656004 183192 656056
rect 183244 656044 183250 656056
rect 537478 656044 537484 656056
rect 183244 656016 537484 656044
rect 183244 656004 183250 656016
rect 537478 656004 537484 656016
rect 537536 656004 537542 656056
rect 172330 655936 172336 655988
rect 172388 655976 172394 655988
rect 537662 655976 537668 655988
rect 172388 655948 537668 655976
rect 172388 655936 172394 655948
rect 537662 655936 537668 655948
rect 537720 655936 537726 655988
rect 161290 655868 161296 655920
rect 161348 655908 161354 655920
rect 538950 655908 538956 655920
rect 161348 655880 538956 655908
rect 161348 655868 161354 655880
rect 538950 655868 538956 655880
rect 539008 655868 539014 655920
rect 150250 655800 150256 655852
rect 150308 655840 150314 655852
rect 539042 655840 539048 655852
rect 150308 655812 539048 655840
rect 150308 655800 150314 655812
rect 539042 655800 539048 655812
rect 539100 655800 539106 655852
rect 85482 655732 85488 655784
rect 85540 655772 85546 655784
rect 537754 655772 537760 655784
rect 85540 655744 537760 655772
rect 85540 655732 85546 655744
rect 537754 655732 537760 655744
rect 537812 655732 537818 655784
rect 74350 655664 74356 655716
rect 74408 655704 74414 655716
rect 537938 655704 537944 655716
rect 74408 655676 537944 655704
rect 74408 655664 74414 655676
rect 537938 655664 537944 655676
rect 537996 655664 538002 655716
rect 63954 655596 63960 655648
rect 64012 655636 64018 655648
rect 538030 655636 538036 655648
rect 64012 655608 538036 655636
rect 64012 655596 64018 655608
rect 538030 655596 538036 655608
rect 538088 655596 538094 655648
rect 53098 655528 53104 655580
rect 53156 655568 53162 655580
rect 538122 655568 538128 655580
rect 53156 655540 538128 655568
rect 53156 655528 53162 655540
rect 538122 655528 538128 655540
rect 538180 655528 538186 655580
rect 13814 654848 13820 654900
rect 13872 654888 13878 654900
rect 40034 654888 40040 654900
rect 13872 654860 40040 654888
rect 13872 654848 13878 654860
rect 40034 654848 40040 654860
rect 40092 654848 40098 654900
rect 492582 654848 492588 654900
rect 492640 654888 492646 654900
rect 580902 654888 580908 654900
rect 492640 654860 580908 654888
rect 492640 654848 492646 654860
rect 580902 654848 580908 654860
rect 580960 654848 580966 654900
rect 13906 654780 13912 654832
rect 13964 654820 13970 654832
rect 104894 654820 104900 654832
rect 13964 654792 104900 654820
rect 13964 654780 13970 654792
rect 104894 654780 104900 654792
rect 104952 654780 104958 654832
rect 464982 654780 464988 654832
rect 465040 654820 465046 654832
rect 580166 654820 580172 654832
rect 465040 654792 580172 654820
rect 465040 654780 465046 654792
rect 580166 654780 580172 654792
rect 580224 654780 580230 654832
rect 520366 654712 520372 654764
rect 520424 654752 520430 654764
rect 520424 654724 521654 654752
rect 520424 654712 520430 654724
rect 107378 654644 107384 654696
rect 107436 654684 107442 654696
rect 520182 654684 520188 654696
rect 107436 654656 520188 654684
rect 107436 654644 107442 654656
rect 520182 654644 520188 654656
rect 520240 654644 520246 654696
rect 521626 654684 521654 654724
rect 537846 654684 537852 654696
rect 521626 654656 537852 654684
rect 537846 654644 537852 654656
rect 537904 654644 537910 654696
rect 356514 654576 356520 654628
rect 356572 654616 356578 654628
rect 516778 654616 516784 654628
rect 356572 654588 516784 654616
rect 356572 654576 356578 654588
rect 516778 654576 516784 654588
rect 516836 654576 516842 654628
rect 518158 654576 518164 654628
rect 518216 654616 518222 654628
rect 518216 654588 520320 654616
rect 518216 654576 518222 654588
rect 345658 654508 345664 654560
rect 345716 654548 345722 654560
rect 520182 654548 520188 654560
rect 345716 654520 520188 654548
rect 345716 654508 345722 654520
rect 520182 654508 520188 654520
rect 520240 654508 520246 654560
rect 334802 654440 334808 654492
rect 334860 654480 334866 654492
rect 515214 654480 515220 654492
rect 334860 654452 515220 654480
rect 334860 654440 334866 654452
rect 515214 654440 515220 654452
rect 515272 654440 515278 654492
rect 520292 654480 520320 654588
rect 521608 654576 521614 654628
rect 521666 654616 521672 654628
rect 536098 654616 536104 654628
rect 521666 654588 536104 654616
rect 521666 654576 521672 654588
rect 536098 654576 536104 654588
rect 536156 654576 536162 654628
rect 520366 654508 520372 654560
rect 520424 654548 520430 654560
rect 538858 654548 538864 654560
rect 520424 654520 538864 654548
rect 520424 654508 520430 654520
rect 538858 654508 538864 654520
rect 538916 654508 538922 654560
rect 518268 654452 519032 654480
rect 520292 654452 520688 654480
rect 226242 654372 226248 654424
rect 226300 654412 226306 654424
rect 226300 654384 229094 654412
rect 226300 654372 226306 654384
rect 229066 654208 229094 654384
rect 258994 654372 259000 654424
rect 259052 654412 259058 654424
rect 259052 654384 267734 654412
rect 259052 654372 259058 654384
rect 267706 654276 267734 654384
rect 313090 654372 313096 654424
rect 313148 654412 313154 654424
rect 313148 654384 316034 654412
rect 313148 654372 313154 654384
rect 316006 654344 316034 654384
rect 323946 654372 323952 654424
rect 324004 654412 324010 654424
rect 518066 654412 518072 654424
rect 324004 654384 518072 654412
rect 324004 654372 324010 654384
rect 518066 654372 518072 654384
rect 518124 654372 518130 654424
rect 518158 654372 518164 654424
rect 518216 654372 518222 654424
rect 518176 654344 518204 654372
rect 316006 654316 518204 654344
rect 518268 654276 518296 654452
rect 518710 654372 518716 654424
rect 518768 654372 518774 654424
rect 519004 654412 519032 654452
rect 519004 654384 520504 654412
rect 267706 654248 518296 654276
rect 518728 654208 518756 654372
rect 520476 654276 520504 654384
rect 520660 654344 520688 654452
rect 521608 654440 521614 654492
rect 521666 654480 521672 654492
rect 580258 654480 580264 654492
rect 521666 654452 580264 654480
rect 521666 654440 521672 654452
rect 580258 654440 580264 654452
rect 580316 654440 580322 654492
rect 520734 654372 520740 654424
rect 520792 654412 520798 654424
rect 580350 654412 580356 654424
rect 520792 654384 580356 654412
rect 520792 654372 520798 654384
rect 580350 654372 580356 654384
rect 580408 654372 580414 654424
rect 580442 654344 580448 654356
rect 520660 654316 580448 654344
rect 580442 654304 580448 654316
rect 580500 654304 580506 654356
rect 539318 654276 539324 654288
rect 520476 654248 539324 654276
rect 539318 654236 539324 654248
rect 539376 654236 539382 654288
rect 229066 654180 509234 654208
rect 518728 654180 525104 654208
rect 509206 654140 509234 654180
rect 525076 654140 525104 654180
rect 534810 654140 534816 654152
rect 509206 654112 510614 654140
rect 525076 654112 534816 654140
rect 510586 654004 510614 654112
rect 534810 654100 534816 654112
rect 534868 654100 534874 654152
rect 536650 654004 536656 654016
rect 510586 653976 511994 654004
rect 511966 653868 511994 653976
rect 519004 653976 536656 654004
rect 519004 653868 519032 653976
rect 536650 653964 536656 653976
rect 536708 653964 536714 654016
rect 511966 653840 519032 653868
rect 535270 644376 535276 644428
rect 535328 644416 535334 644428
rect 579982 644416 579988 644428
rect 535328 644388 579988 644416
rect 535328 644376 535334 644388
rect 579982 644376 579988 644388
rect 580040 644376 580046 644428
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 10318 632108 10324 632120
rect 3476 632080 10324 632108
rect 3476 632068 3482 632080
rect 10318 632068 10324 632080
rect 10376 632068 10382 632120
rect 536650 632000 536656 632052
rect 536708 632040 536714 632052
rect 579982 632040 579988 632052
rect 536708 632012 579988 632040
rect 536708 632000 536714 632012
rect 579982 632000 579988 632012
rect 580040 632000 580046 632052
rect 538122 618196 538128 618248
rect 538180 618236 538186 618248
rect 579982 618236 579988 618248
rect 538180 618208 579988 618236
rect 538180 618196 538186 618208
rect 579982 618196 579988 618208
rect 580040 618196 580046 618248
rect 535178 607860 535184 607912
rect 535236 607900 535242 607912
rect 580626 607900 580632 607912
rect 535236 607872 580632 607900
rect 535236 607860 535242 607872
rect 580626 607860 580632 607872
rect 580684 607860 580690 607912
rect 3510 579640 3516 579692
rect 3568 579680 3574 579692
rect 11698 579680 11704 579692
rect 3568 579652 11704 579680
rect 3568 579640 3574 579652
rect 11698 579640 11704 579652
rect 11756 579640 11762 579692
rect 6914 568488 6920 568540
rect 6972 568528 6978 568540
rect 12434 568528 12440 568540
rect 6972 568500 12440 568528
rect 6972 568488 6978 568500
rect 12434 568488 12440 568500
rect 12492 568488 12498 568540
rect 538030 564340 538036 564392
rect 538088 564380 538094 564392
rect 580166 564380 580172 564392
rect 538088 564352 580172 564380
rect 538088 564340 538094 564352
rect 580166 564340 580172 564352
rect 580224 564340 580230 564392
rect 3602 542308 3608 542360
rect 3660 542348 3666 542360
rect 12434 542348 12440 542360
rect 3660 542320 12440 542348
rect 3660 542308 3666 542320
rect 12434 542308 12440 542320
rect 12492 542308 12498 542360
rect 3694 528504 3700 528556
rect 3752 528544 3758 528556
rect 12434 528544 12440 528556
rect 3752 528516 12440 528544
rect 3752 528504 3758 528516
rect 12434 528504 12440 528516
rect 12492 528504 12498 528556
rect 2958 527144 2964 527196
rect 3016 527184 3022 527196
rect 7558 527184 7564 527196
rect 3016 527156 7564 527184
rect 3016 527144 3022 527156
rect 7558 527144 7564 527156
rect 7616 527144 7622 527196
rect 540422 525716 540428 525768
rect 540480 525756 540486 525768
rect 580166 525756 580172 525768
rect 540480 525728 580172 525756
rect 540480 525716 540486 525728
rect 580166 525716 580172 525728
rect 580224 525716 580230 525768
rect 10410 514768 10416 514820
rect 10468 514808 10474 514820
rect 12434 514808 12440 514820
rect 10468 514780 12440 514808
rect 10468 514768 10474 514780
rect 12434 514768 12440 514780
rect 12492 514768 12498 514820
rect 537938 511912 537944 511964
rect 537996 511952 538002 511964
rect 580166 511952 580172 511964
rect 537996 511924 580172 511952
rect 537996 511912 538002 511924
rect 580166 511912 580172 511924
rect 580224 511912 580230 511964
rect 3234 502256 3240 502308
rect 3292 502296 3298 502308
rect 10410 502296 10416 502308
rect 3292 502268 10416 502296
rect 3292 502256 3298 502268
rect 10410 502256 10416 502268
rect 10468 502256 10474 502308
rect 7650 500964 7656 501016
rect 7708 501004 7714 501016
rect 12434 501004 12440 501016
rect 7708 500976 12440 501004
rect 7708 500964 7714 500976
rect 12434 500964 12440 500976
rect 12492 500964 12498 501016
rect 9030 487160 9036 487212
rect 9088 487200 9094 487212
rect 12434 487200 12440 487212
rect 9088 487172 12440 487200
rect 9088 487160 9094 487172
rect 12434 487160 12440 487172
rect 12492 487160 12498 487212
rect 535086 485732 535092 485784
rect 535144 485772 535150 485784
rect 580166 485772 580172 485784
rect 535144 485744 580172 485772
rect 535144 485732 535150 485744
rect 580166 485732 580172 485744
rect 580224 485732 580230 485784
rect 2774 475600 2780 475652
rect 2832 475640 2838 475652
rect 4890 475640 4896 475652
rect 2832 475612 4896 475640
rect 2832 475600 2838 475612
rect 4890 475600 4896 475612
rect 4948 475600 4954 475652
rect 7742 474716 7748 474768
rect 7800 474756 7806 474768
rect 12434 474756 12440 474768
rect 7800 474728 12440 474756
rect 7800 474716 7806 474728
rect 12434 474716 12440 474728
rect 12492 474716 12498 474768
rect 539318 471928 539324 471980
rect 539376 471968 539382 471980
rect 579798 471968 579804 471980
rect 539376 471940 579804 471968
rect 539376 471928 539382 471940
rect 579798 471928 579804 471940
rect 579856 471928 579862 471980
rect 8938 461252 8944 461304
rect 8996 461292 9002 461304
rect 12434 461292 12440 461304
rect 8996 461264 12440 461292
rect 8996 461252 9002 461264
rect 12434 461252 12440 461264
rect 12492 461252 12498 461304
rect 537754 458124 537760 458176
rect 537812 458164 537818 458176
rect 580166 458164 580172 458176
rect 537812 458136 580172 458164
rect 537812 458124 537818 458136
rect 580166 458124 580172 458136
rect 580224 458124 580230 458176
rect 3326 449556 3332 449608
rect 3384 449596 3390 449608
rect 7650 449596 7656 449608
rect 3384 449568 7656 449596
rect 3384 449556 3390 449568
rect 7650 449556 7656 449568
rect 7708 449556 7714 449608
rect 536558 431876 536564 431928
rect 536616 431916 536622 431928
rect 580166 431916 580172 431928
rect 536616 431888 580172 431916
rect 536616 431876 536622 431888
rect 580166 431876 580172 431888
rect 580224 431876 580230 431928
rect 3326 422288 3332 422340
rect 3384 422328 3390 422340
rect 10410 422328 10416 422340
rect 3384 422300 10416 422328
rect 3384 422288 3390 422300
rect 10410 422288 10416 422300
rect 10468 422288 10474 422340
rect 540330 419432 540336 419484
rect 540388 419472 540394 419484
rect 580166 419472 580172 419484
rect 540388 419444 580172 419472
rect 540388 419432 540394 419444
rect 580166 419432 580172 419444
rect 580224 419432 580230 419484
rect 3234 409844 3240 409896
rect 3292 409884 3298 409896
rect 7650 409884 7656 409896
rect 3292 409856 7656 409884
rect 3292 409844 3298 409856
rect 7650 409844 7656 409856
rect 7708 409844 7714 409896
rect 3234 397944 3240 397996
rect 3292 397984 3298 397996
rect 9030 397984 9036 397996
rect 3292 397956 9036 397984
rect 3292 397944 3298 397956
rect 9030 397944 9036 397956
rect 9088 397944 9094 397996
rect 534994 379448 535000 379500
rect 535052 379488 535058 379500
rect 580166 379488 580172 379500
rect 535052 379460 580172 379488
rect 535052 379448 535058 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 3326 371220 3332 371272
rect 3384 371260 3390 371272
rect 11882 371260 11888 371272
rect 3384 371232 11888 371260
rect 3384 371220 3390 371232
rect 11882 371220 11888 371232
rect 11940 371220 11946 371272
rect 540238 365644 540244 365696
rect 540296 365684 540302 365696
rect 580166 365684 580172 365696
rect 540296 365656 580172 365684
rect 540296 365644 540302 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 537846 353200 537852 353252
rect 537904 353240 537910 353252
rect 579614 353240 579620 353252
rect 537904 353212 579620 353240
rect 537904 353200 537910 353212
rect 579614 353200 579620 353212
rect 579672 353200 579678 353252
rect 2958 346332 2964 346384
rect 3016 346372 3022 346384
rect 7742 346372 7748 346384
rect 3016 346344 7748 346372
rect 3016 346332 3022 346344
rect 7742 346332 7748 346344
rect 7800 346332 7806 346384
rect 3418 328380 3424 328432
rect 3476 328420 3482 328432
rect 12434 328420 12440 328432
rect 3476 328392 12440 328420
rect 3476 328380 3482 328392
rect 12434 328380 12440 328392
rect 12492 328380 12498 328432
rect 536466 325592 536472 325644
rect 536524 325632 536530 325644
rect 580166 325632 580172 325644
rect 536524 325604 580172 325632
rect 536524 325592 536530 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 3418 318792 3424 318844
rect 3476 318832 3482 318844
rect 13078 318832 13084 318844
rect 3476 318804 13084 318832
rect 3476 318792 3482 318804
rect 13078 318792 13084 318804
rect 13136 318792 13142 318844
rect 3510 315936 3516 315988
rect 3568 315976 3574 315988
rect 12434 315976 12440 315988
rect 3568 315948 12440 315976
rect 3568 315936 3574 315948
rect 12434 315936 12440 315948
rect 12492 315936 12498 315988
rect 536374 313216 536380 313268
rect 536432 313256 536438 313268
rect 580166 313256 580172 313268
rect 536432 313228 580172 313256
rect 536432 313216 536438 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 3602 302132 3608 302184
rect 3660 302172 3666 302184
rect 12434 302172 12440 302184
rect 3660 302144 12440 302172
rect 3660 302132 3666 302144
rect 12434 302132 12440 302144
rect 12492 302132 12498 302184
rect 3326 293564 3332 293616
rect 3384 293604 3390 293616
rect 8938 293604 8944 293616
rect 3384 293576 8944 293604
rect 3384 293564 3390 293576
rect 8938 293564 8944 293576
rect 8996 293564 9002 293616
rect 3694 288328 3700 288380
rect 3752 288368 3758 288380
rect 12434 288368 12440 288380
rect 3752 288340 12440 288368
rect 3752 288328 3758 288340
rect 12434 288328 12440 288340
rect 12492 288328 12498 288380
rect 7650 275952 7656 276004
rect 7708 275992 7714 276004
rect 12434 275992 12440 276004
rect 7708 275964 12440 275992
rect 7708 275952 7714 275964
rect 12434 275952 12440 275964
rect 12492 275952 12498 276004
rect 536282 273164 536288 273216
rect 536340 273204 536346 273216
rect 580166 273204 580172 273216
rect 536340 273176 580172 273204
rect 536340 273164 536346 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 3786 262148 3792 262200
rect 3844 262188 3850 262200
rect 12434 262188 12440 262200
rect 3844 262160 12440 262188
rect 3844 262148 3850 262160
rect 12434 262148 12440 262160
rect 12492 262148 12498 262200
rect 536190 259360 536196 259412
rect 536248 259400 536254 259412
rect 579798 259400 579804 259412
rect 536248 259372 579804 259400
rect 536248 259360 536254 259372
rect 579798 259360 579804 259372
rect 579856 259360 579862 259412
rect 3418 248344 3424 248396
rect 3476 248384 3482 248396
rect 12434 248384 12440 248396
rect 3476 248356 12440 248384
rect 3476 248344 3482 248356
rect 12434 248344 12440 248356
rect 12492 248344 12498 248396
rect 539226 233180 539232 233232
rect 539284 233220 539290 233232
rect 579982 233220 579988 233232
rect 539284 233192 579988 233220
rect 539284 233180 539290 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 539134 193128 539140 193180
rect 539192 193168 539198 193180
rect 580166 193168 580172 193180
rect 539192 193140 580172 193168
rect 539192 193128 539198 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 539042 166948 539048 167000
rect 539100 166988 539106 167000
rect 580166 166988 580172 167000
rect 539100 166960 580172 166988
rect 539100 166948 539106 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 534902 153144 534908 153196
rect 534960 153184 534966 153196
rect 579798 153184 579804 153196
rect 534960 153156 579804 153184
rect 534960 153144 534966 153156
rect 579798 153144 579804 153156
rect 579856 153144 579862 153196
rect 4798 128256 4804 128308
rect 4856 128296 4862 128308
rect 12434 128296 12440 128308
rect 4856 128268 12440 128296
rect 4856 128256 4862 128268
rect 12434 128256 12440 128268
rect 12492 128256 12498 128308
rect 538950 126896 538956 126948
rect 539008 126936 539014 126948
rect 580166 126936 580172 126948
rect 539008 126908 580172 126936
rect 539008 126896 539014 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 10318 115880 10324 115932
rect 10376 115920 10382 115932
rect 12434 115920 12440 115932
rect 10376 115892 12440 115920
rect 10376 115880 10382 115892
rect 12434 115880 12440 115892
rect 12492 115880 12498 115932
rect 534810 113092 534816 113144
rect 534868 113132 534874 113144
rect 579798 113132 579804 113144
rect 534868 113104 579804 113132
rect 534868 113092 534874 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 538858 100648 538864 100700
rect 538916 100688 538922 100700
rect 580166 100688 580172 100700
rect 538916 100660 580172 100688
rect 538916 100648 538922 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 7558 89632 7564 89684
rect 7616 89672 7622 89684
rect 12434 89672 12440 89684
rect 7616 89644 12440 89672
rect 7616 89632 7622 89644
rect 12434 89632 12440 89644
rect 12492 89632 12498 89684
rect 537662 86912 537668 86964
rect 537720 86952 537726 86964
rect 580166 86952 580172 86964
rect 537720 86924 580172 86952
rect 537720 86912 537726 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 4890 75828 4896 75880
rect 4948 75868 4954 75880
rect 12434 75868 12440 75880
rect 4948 75840 12440 75868
rect 4948 75828 4954 75840
rect 12434 75828 12440 75840
rect 12492 75828 12498 75880
rect 534718 73108 534724 73160
rect 534776 73148 534782 73160
rect 580166 73148 580172 73160
rect 534776 73120 580172 73148
rect 534776 73108 534782 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 10410 62024 10416 62076
rect 10468 62064 10474 62076
rect 12802 62064 12808 62076
rect 10468 62036 12808 62064
rect 10468 62024 10474 62036
rect 12802 62024 12808 62036
rect 12860 62024 12866 62076
rect 536098 60664 536104 60716
rect 536156 60704 536162 60716
rect 580166 60704 580172 60716
rect 536156 60676 580172 60704
rect 536156 60664 536162 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 537478 46860 537484 46912
rect 537536 46900 537542 46912
rect 580166 46900 580172 46912
rect 537536 46872 580172 46900
rect 537536 46860 537542 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 537570 33056 537576 33108
rect 537628 33096 537634 33108
rect 580166 33096 580172 33108
rect 537628 33068 580172 33096
rect 537628 33056 537634 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 537754 20612 537760 20664
rect 537812 20652 537818 20664
rect 579982 20652 579988 20664
rect 537812 20624 579988 20652
rect 537812 20612 537818 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 13722 13744 13728 13796
rect 13780 13784 13786 13796
rect 52086 13784 52092 13796
rect 13780 13756 52092 13784
rect 13780 13744 13786 13756
rect 52086 13744 52092 13756
rect 52144 13744 52150 13796
rect 3510 13676 3516 13728
rect 3568 13716 3574 13728
rect 423490 13716 423496 13728
rect 3568 13688 423496 13716
rect 3568 13676 3574 13688
rect 423490 13676 423496 13688
rect 423548 13676 423554 13728
rect 3694 13608 3700 13660
rect 3752 13648 3758 13660
rect 349154 13648 349160 13660
rect 3752 13620 349160 13648
rect 3752 13608 3758 13620
rect 349154 13608 349160 13620
rect 349212 13608 349218 13660
rect 3602 13540 3608 13592
rect 3660 13580 3666 13592
rect 200574 13580 200580 13592
rect 3660 13552 200580 13580
rect 3660 13540 3666 13552
rect 200574 13540 200580 13552
rect 200632 13540 200638 13592
rect 3418 13472 3424 13524
rect 3476 13512 3482 13524
rect 126330 13512 126336 13524
rect 3476 13484 126336 13512
rect 3476 13472 3482 13484
rect 126330 13472 126336 13484
rect 126388 13472 126394 13524
rect 52086 13064 52092 13116
rect 52144 13104 52150 13116
rect 579614 13104 579620 13116
rect 52144 13076 579620 13104
rect 52144 13064 52150 13076
rect 579614 13064 579620 13076
rect 579672 13064 579678 13116
rect 537846 6808 537852 6860
rect 537904 6848 537910 6860
rect 580166 6848 580172 6860
rect 537904 6820 580172 6848
rect 537904 6808 537910 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
<< via1 >>
rect 71780 702992 71832 703044
rect 72976 702992 73028 703044
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 13728 700816 13780 700868
rect 24308 700816 24360 700868
rect 13636 700748 13688 700800
rect 89168 700748 89220 700800
rect 13084 700680 13136 700732
rect 137836 700680 137888 700732
rect 365720 700680 365772 700732
rect 462320 700680 462372 700732
rect 13452 700612 13504 700664
rect 218980 700612 219032 700664
rect 376760 700612 376812 700664
rect 527180 700612 527232 700664
rect 13360 700544 13412 700596
rect 283840 700544 283892 700596
rect 330484 700544 330536 700596
rect 494796 700544 494848 700596
rect 13544 700476 13596 700528
rect 154120 700476 154172 700528
rect 193220 700476 193272 700528
rect 478512 700476 478564 700528
rect 13268 700408 13320 700460
rect 348792 700408 348844 700460
rect 398104 700408 398156 700460
rect 559656 700408 559708 700460
rect 12992 700340 13044 700392
rect 202788 700340 202840 700392
rect 204260 700340 204312 700392
rect 543464 700340 543516 700392
rect 21364 700272 21416 700324
rect 413652 700272 413704 700324
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 387800 696940 387852 696992
rect 580172 696940 580224 696992
rect 2780 683680 2832 683732
rect 4804 683680 4856 683732
rect 215300 683136 215352 683188
rect 580172 683136 580224 683188
rect 3516 670692 3568 670744
rect 11796 670692 11848 670744
rect 41512 670692 41564 670744
rect 580172 670692 580224 670744
rect 14280 659064 14332 659116
rect 266360 659064 266412 659116
rect 14372 658996 14424 659048
rect 331220 658996 331272 659048
rect 14464 658928 14516 658980
rect 397460 658928 397512 658980
rect 442908 657772 442960 657824
rect 536564 657772 536616 657824
rect 14004 657704 14056 657756
rect 169760 657704 169812 657756
rect 237288 657704 237340 657756
rect 464988 657704 465040 657756
rect 486424 657704 486476 657756
rect 539232 657704 539284 657756
rect 14188 657636 14240 657688
rect 299480 657636 299532 657688
rect 475568 657636 475620 657688
rect 536288 657636 536340 657688
rect 20628 657568 20680 657620
rect 330484 657568 330536 657620
rect 421472 657568 421524 657620
rect 492588 657568 492640 657620
rect 497280 657568 497332 657620
rect 539140 657568 539192 657620
rect 31392 657500 31444 657552
rect 398104 657500 398156 657552
rect 453856 657500 453908 657552
rect 535000 657500 535052 657552
rect 464712 657432 464764 657484
rect 536472 657432 536524 657484
rect 302148 657364 302200 657416
rect 536196 657364 536248 657416
rect 291016 657296 291068 657348
rect 536380 657296 536432 657348
rect 118056 657228 118108 657280
rect 365628 657228 365680 657280
rect 399760 657228 399812 657280
rect 535276 657228 535328 657280
rect 280712 657160 280764 657212
rect 540244 657160 540296 657212
rect 269856 657092 269908 657144
rect 540336 657092 540388 657144
rect 248052 657024 248104 657076
rect 540428 657024 540480 657076
rect 128912 656956 128964 657008
rect 430580 656956 430632 657008
rect 432328 656956 432380 657008
rect 535092 656956 535144 657008
rect 3424 656888 3476 656940
rect 11888 656888 11940 656940
rect 96528 656888 96580 656940
rect 453948 656888 454000 656940
rect 529848 656888 529900 656940
rect 534724 656888 534776 656940
rect 13176 656276 13228 656328
rect 21364 656276 21416 656328
rect 453948 656276 454000 656328
rect 580816 656276 580868 656328
rect 12900 656208 12952 656260
rect 71780 656208 71832 656260
rect 430580 656208 430632 656260
rect 580540 656208 580592 656260
rect 14096 656140 14148 656192
rect 234620 656140 234672 656192
rect 365628 656140 365680 656192
rect 580724 656140 580776 656192
rect 507676 656072 507728 656124
rect 534908 656072 534960 656124
rect 183192 656004 183244 656056
rect 537484 656004 537536 656056
rect 172336 655936 172388 655988
rect 537668 655936 537720 655988
rect 161296 655868 161348 655920
rect 538956 655868 539008 655920
rect 150256 655800 150308 655852
rect 539048 655800 539100 655852
rect 85488 655732 85540 655784
rect 537760 655732 537812 655784
rect 74356 655664 74408 655716
rect 537944 655664 537996 655716
rect 63960 655596 64012 655648
rect 538036 655596 538088 655648
rect 53104 655528 53156 655580
rect 538128 655528 538180 655580
rect 13820 654848 13872 654900
rect 40040 654848 40092 654900
rect 492588 654848 492640 654900
rect 580908 654848 580960 654900
rect 13912 654780 13964 654832
rect 104900 654780 104952 654832
rect 464988 654780 465040 654832
rect 580172 654780 580224 654832
rect 520372 654712 520424 654764
rect 107384 654644 107436 654696
rect 520188 654644 520240 654696
rect 537852 654644 537904 654696
rect 356520 654576 356572 654628
rect 516784 654576 516836 654628
rect 518164 654576 518216 654628
rect 345664 654508 345716 654560
rect 520188 654508 520240 654560
rect 334808 654440 334860 654492
rect 515220 654440 515272 654492
rect 521614 654576 521666 654628
rect 536104 654576 536156 654628
rect 520372 654508 520424 654560
rect 538864 654508 538916 654560
rect 226248 654372 226300 654424
rect 259000 654372 259052 654424
rect 313096 654372 313148 654424
rect 323952 654372 324004 654424
rect 518072 654372 518124 654424
rect 518164 654372 518216 654424
rect 518716 654372 518768 654424
rect 521614 654440 521666 654492
rect 580264 654440 580316 654492
rect 520740 654372 520792 654424
rect 580356 654372 580408 654424
rect 580448 654304 580500 654356
rect 539324 654236 539376 654288
rect 534816 654100 534868 654152
rect 536656 653964 536708 654016
rect 535276 644376 535328 644428
rect 579988 644376 580040 644428
rect 3424 632068 3476 632120
rect 10324 632068 10376 632120
rect 536656 632000 536708 632052
rect 579988 632000 580040 632052
rect 538128 618196 538180 618248
rect 579988 618196 580040 618248
rect 535184 607860 535236 607912
rect 580632 607860 580684 607912
rect 3516 579640 3568 579692
rect 11704 579640 11756 579692
rect 6920 568488 6972 568540
rect 12440 568488 12492 568540
rect 538036 564340 538088 564392
rect 580172 564340 580224 564392
rect 3608 542308 3660 542360
rect 12440 542308 12492 542360
rect 3700 528504 3752 528556
rect 12440 528504 12492 528556
rect 2964 527144 3016 527196
rect 7564 527144 7616 527196
rect 540428 525716 540480 525768
rect 580172 525716 580224 525768
rect 10416 514768 10468 514820
rect 12440 514768 12492 514820
rect 537944 511912 537996 511964
rect 580172 511912 580224 511964
rect 3240 502256 3292 502308
rect 10416 502256 10468 502308
rect 7656 500964 7708 501016
rect 12440 500964 12492 501016
rect 9036 487160 9088 487212
rect 12440 487160 12492 487212
rect 535092 485732 535144 485784
rect 580172 485732 580224 485784
rect 2780 475600 2832 475652
rect 4896 475600 4948 475652
rect 7748 474716 7800 474768
rect 12440 474716 12492 474768
rect 539324 471928 539376 471980
rect 579804 471928 579856 471980
rect 8944 461252 8996 461304
rect 12440 461252 12492 461304
rect 537760 458124 537812 458176
rect 580172 458124 580224 458176
rect 3332 449556 3384 449608
rect 7656 449556 7708 449608
rect 536564 431876 536616 431928
rect 580172 431876 580224 431928
rect 3332 422288 3384 422340
rect 10416 422288 10468 422340
rect 540336 419432 540388 419484
rect 580172 419432 580224 419484
rect 3240 409844 3292 409896
rect 7656 409844 7708 409896
rect 3240 397944 3292 397996
rect 9036 397944 9088 397996
rect 535000 379448 535052 379500
rect 580172 379448 580224 379500
rect 3332 371220 3384 371272
rect 11888 371220 11940 371272
rect 540244 365644 540296 365696
rect 580172 365644 580224 365696
rect 537852 353200 537904 353252
rect 579620 353200 579672 353252
rect 2964 346332 3016 346384
rect 7748 346332 7800 346384
rect 3424 328380 3476 328432
rect 12440 328380 12492 328432
rect 536472 325592 536524 325644
rect 580172 325592 580224 325644
rect 3424 318792 3476 318844
rect 13084 318792 13136 318844
rect 3516 315936 3568 315988
rect 12440 315936 12492 315988
rect 536380 313216 536432 313268
rect 580172 313216 580224 313268
rect 3608 302132 3660 302184
rect 12440 302132 12492 302184
rect 3332 293564 3384 293616
rect 8944 293564 8996 293616
rect 3700 288328 3752 288380
rect 12440 288328 12492 288380
rect 7656 275952 7708 276004
rect 12440 275952 12492 276004
rect 536288 273164 536340 273216
rect 580172 273164 580224 273216
rect 3792 262148 3844 262200
rect 12440 262148 12492 262200
rect 536196 259360 536248 259412
rect 579804 259360 579856 259412
rect 3424 248344 3476 248396
rect 12440 248344 12492 248396
rect 539232 233180 539284 233232
rect 579988 233180 580040 233232
rect 539140 193128 539192 193180
rect 580172 193128 580224 193180
rect 539048 166948 539100 167000
rect 580172 166948 580224 167000
rect 534908 153144 534960 153196
rect 579804 153144 579856 153196
rect 4804 128256 4856 128308
rect 12440 128256 12492 128308
rect 538956 126896 539008 126948
rect 580172 126896 580224 126948
rect 10324 115880 10376 115932
rect 12440 115880 12492 115932
rect 534816 113092 534868 113144
rect 579804 113092 579856 113144
rect 538864 100648 538916 100700
rect 580172 100648 580224 100700
rect 7564 89632 7616 89684
rect 12440 89632 12492 89684
rect 537668 86912 537720 86964
rect 580172 86912 580224 86964
rect 4896 75828 4948 75880
rect 12440 75828 12492 75880
rect 534724 73108 534776 73160
rect 580172 73108 580224 73160
rect 10416 62024 10468 62076
rect 12808 62024 12860 62076
rect 536104 60664 536156 60716
rect 580172 60664 580224 60716
rect 537484 46860 537536 46912
rect 580172 46860 580224 46912
rect 537576 33056 537628 33108
rect 580172 33056 580224 33108
rect 537760 20612 537812 20664
rect 579988 20612 580040 20664
rect 13728 13744 13780 13796
rect 52092 13744 52144 13796
rect 3516 13676 3568 13728
rect 423496 13676 423548 13728
rect 3700 13608 3752 13660
rect 349160 13608 349212 13660
rect 3608 13540 3660 13592
rect 200580 13540 200632 13592
rect 3424 13472 3476 13524
rect 126336 13472 126388 13524
rect 52092 13064 52144 13116
rect 579620 13064 579672 13116
rect 537852 6808 537904 6860
rect 580172 6808 580224 6860
<< metal2 >>
rect 6932 703582 7972 703610
rect 2778 684312 2834 684321
rect 2778 684247 2834 684256
rect 2792 683738 2820 684247
rect 2780 683732 2832 683738
rect 2780 683674 2832 683680
rect 4804 683732 4856 683738
rect 4804 683674 4856 683680
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3422 619168 3478 619177
rect 3422 619103 3478 619112
rect 2962 527912 3018 527921
rect 2962 527847 3018 527856
rect 2976 527202 3004 527847
rect 2964 527196 3016 527202
rect 2964 527138 3016 527144
rect 3240 502308 3292 502314
rect 3240 502250 3292 502256
rect 3252 501809 3280 502250
rect 3238 501800 3294 501809
rect 3238 501735 3294 501744
rect 2778 475688 2834 475697
rect 2778 475623 2780 475632
rect 2832 475623 2834 475632
rect 2780 475594 2832 475600
rect 3332 449608 3384 449614
rect 3330 449576 3332 449585
rect 3384 449576 3386 449585
rect 3330 449511 3386 449520
rect 3330 423600 3386 423609
rect 3330 423535 3386 423544
rect 3344 422346 3372 423535
rect 3332 422340 3384 422346
rect 3332 422282 3384 422288
rect 3238 410544 3294 410553
rect 3238 410479 3294 410488
rect 3252 409902 3280 410479
rect 3240 409896 3292 409902
rect 3240 409838 3292 409844
rect 3240 397996 3292 398002
rect 3240 397938 3292 397944
rect 3252 397497 3280 397938
rect 3238 397488 3294 397497
rect 3238 397423 3294 397432
rect 3330 371376 3386 371385
rect 3330 371311 3386 371320
rect 3344 371278 3372 371311
rect 3332 371272 3384 371278
rect 3332 371214 3384 371220
rect 2964 346384 3016 346390
rect 2964 346326 3016 346332
rect 2976 345409 3004 346326
rect 2962 345400 3018 345409
rect 2962 345335 3018 345344
rect 3436 328438 3464 619103
rect 3606 606112 3662 606121
rect 3606 606047 3662 606056
rect 3514 580000 3570 580009
rect 3514 579935 3570 579944
rect 3528 579698 3556 579935
rect 3516 579692 3568 579698
rect 3516 579634 3568 579640
rect 3514 566944 3570 566953
rect 3514 566879 3570 566888
rect 3424 328432 3476 328438
rect 3424 328374 3476 328380
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 318850 3464 319223
rect 3424 318844 3476 318850
rect 3424 318786 3476 318792
rect 3528 315994 3556 566879
rect 3620 542366 3648 606047
rect 3698 553888 3754 553897
rect 3698 553823 3754 553832
rect 3608 542360 3660 542366
rect 3608 542302 3660 542308
rect 3712 528562 3740 553823
rect 3700 528556 3752 528562
rect 3700 528498 3752 528504
rect 3606 514856 3662 514865
rect 3606 514791 3662 514800
rect 3516 315988 3568 315994
rect 3516 315930 3568 315936
rect 3422 306232 3478 306241
rect 3422 306167 3478 306176
rect 3332 293616 3384 293622
rect 3332 293558 3384 293564
rect 3344 293185 3372 293558
rect 3330 293176 3386 293185
rect 3330 293111 3386 293120
rect 3436 248402 3464 306167
rect 3620 302190 3648 514791
rect 3698 462632 3754 462641
rect 3698 462567 3754 462576
rect 3608 302184 3660 302190
rect 3608 302126 3660 302132
rect 3712 288386 3740 462567
rect 3790 358456 3846 358465
rect 3790 358391 3846 358400
rect 3700 288380 3752 288386
rect 3700 288322 3752 288328
rect 3804 262206 3832 358391
rect 3792 262200 3844 262206
rect 3792 262142 3844 262148
rect 3424 248396 3476 248402
rect 3424 248338 3476 248344
rect 3422 214976 3478 214985
rect 3422 214911 3478 214920
rect 3436 13530 3464 214911
rect 3514 162888 3570 162897
rect 3514 162823 3570 162832
rect 3528 13734 3556 162823
rect 4816 128314 4844 683674
rect 6932 568546 6960 703582
rect 7944 703474 7972 703582
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 703474 8156 703520
rect 7944 703446 8156 703474
rect 24320 700874 24348 703520
rect 13728 700868 13780 700874
rect 13728 700810 13780 700816
rect 24308 700868 24360 700874
rect 24308 700810 24360 700816
rect 13636 700800 13688 700806
rect 13636 700742 13688 700748
rect 13084 700732 13136 700738
rect 13084 700674 13136 700680
rect 12992 700392 13044 700398
rect 12992 700334 13044 700340
rect 11796 670744 11848 670750
rect 11796 670686 11848 670692
rect 10324 632120 10376 632126
rect 10324 632062 10376 632068
rect 6920 568540 6972 568546
rect 6920 568482 6972 568488
rect 7564 527196 7616 527202
rect 7564 527138 7616 527144
rect 4896 475652 4948 475658
rect 4896 475594 4948 475600
rect 4804 128308 4856 128314
rect 4804 128250 4856 128256
rect 3606 110664 3662 110673
rect 3606 110599 3662 110608
rect 3516 13728 3568 13734
rect 3516 13670 3568 13676
rect 3620 13598 3648 110599
rect 4908 75886 4936 475594
rect 7576 89690 7604 527138
rect 7656 501016 7708 501022
rect 7656 500958 7708 500964
rect 7668 449614 7696 500958
rect 9036 487212 9088 487218
rect 9036 487154 9088 487160
rect 7748 474768 7800 474774
rect 7748 474710 7800 474716
rect 7656 449608 7708 449614
rect 7656 449550 7708 449556
rect 7656 409896 7708 409902
rect 7656 409838 7708 409844
rect 7668 276010 7696 409838
rect 7760 346390 7788 474710
rect 8944 461304 8996 461310
rect 8944 461246 8996 461252
rect 7748 346384 7800 346390
rect 7748 346326 7800 346332
rect 8956 293622 8984 461246
rect 9048 398002 9076 487154
rect 9036 397996 9088 398002
rect 9036 397938 9088 397944
rect 8944 293616 8996 293622
rect 8944 293558 8996 293564
rect 7656 276004 7708 276010
rect 7656 275946 7708 275952
rect 10336 115938 10364 632062
rect 11704 579692 11756 579698
rect 11704 579634 11756 579640
rect 10416 514820 10468 514826
rect 10416 514762 10468 514768
rect 10428 502314 10456 514762
rect 10416 502308 10468 502314
rect 10416 502250 10468 502256
rect 10416 422340 10468 422346
rect 10416 422282 10468 422288
rect 10324 115932 10376 115938
rect 10324 115874 10376 115880
rect 7564 89684 7616 89690
rect 7564 89626 7616 89632
rect 4896 75880 4948 75886
rect 4896 75822 4948 75828
rect 3698 71632 3754 71641
rect 3698 71567 3754 71576
rect 3712 13666 3740 71567
rect 10428 62082 10456 422282
rect 11716 102105 11744 579634
rect 11808 342145 11836 670686
rect 11888 656940 11940 656946
rect 11888 656882 11940 656888
rect 11900 555529 11928 656882
rect 12900 656260 12952 656266
rect 12900 656202 12952 656208
rect 12912 582185 12940 656202
rect 13004 608569 13032 700334
rect 12990 608560 13046 608569
rect 12990 608495 13046 608504
rect 13096 595513 13124 700674
rect 13452 700664 13504 700670
rect 13452 700606 13504 700612
rect 13360 700596 13412 700602
rect 13360 700538 13412 700544
rect 13268 700460 13320 700466
rect 13268 700402 13320 700408
rect 13176 656328 13228 656334
rect 13176 656270 13228 656276
rect 13082 595504 13138 595513
rect 13082 595439 13138 595448
rect 12898 582176 12954 582185
rect 12898 582111 12954 582120
rect 12438 568576 12494 568585
rect 12438 568511 12440 568520
rect 12492 568511 12494 568520
rect 12440 568482 12492 568488
rect 11886 555520 11942 555529
rect 11886 555455 11942 555464
rect 12440 542360 12492 542366
rect 12440 542302 12492 542308
rect 12452 542065 12480 542302
rect 12438 542056 12494 542065
rect 12438 541991 12494 542000
rect 12440 528556 12492 528562
rect 12440 528498 12492 528504
rect 12452 528193 12480 528498
rect 12438 528184 12494 528193
rect 12438 528119 12494 528128
rect 12438 514856 12494 514865
rect 12438 514791 12440 514800
rect 12492 514791 12494 514800
rect 12440 514762 12492 514768
rect 12438 501120 12494 501129
rect 12438 501055 12494 501064
rect 12452 501022 12480 501055
rect 12440 501016 12492 501022
rect 12440 500958 12492 500964
rect 12438 487792 12494 487801
rect 12438 487727 12494 487736
rect 12452 487218 12480 487727
rect 12440 487212 12492 487218
rect 12440 487154 12492 487160
rect 12438 474872 12494 474881
rect 12438 474807 12494 474816
rect 12452 474774 12480 474807
rect 12440 474768 12492 474774
rect 12440 474710 12492 474716
rect 12438 461408 12494 461417
rect 12438 461343 12494 461352
rect 12452 461310 12480 461343
rect 12440 461304 12492 461310
rect 12440 461246 12492 461252
rect 13188 435577 13216 656270
rect 13174 435568 13230 435577
rect 13174 435503 13230 435512
rect 13280 421977 13308 700402
rect 13266 421968 13322 421977
rect 13266 421903 13322 421912
rect 13372 408241 13400 700538
rect 13358 408232 13414 408241
rect 13358 408167 13414 408176
rect 13464 395593 13492 700606
rect 13544 700528 13596 700534
rect 13544 700470 13596 700476
rect 13450 395584 13506 395593
rect 13450 395519 13506 395528
rect 13556 382265 13584 700470
rect 13542 382256 13598 382265
rect 13542 382191 13598 382200
rect 11888 371272 11940 371278
rect 11888 371214 11940 371220
rect 11794 342136 11850 342145
rect 11794 342071 11850 342080
rect 11702 102096 11758 102105
rect 11702 102031 11758 102040
rect 10416 62076 10468 62082
rect 10416 62018 10468 62024
rect 11900 48929 11928 371214
rect 13648 368257 13676 700742
rect 13634 368248 13690 368257
rect 13634 368183 13690 368192
rect 13740 355609 13768 700810
rect 21364 700324 21416 700330
rect 21364 700266 21416 700272
rect 14280 659116 14332 659122
rect 14280 659058 14332 659064
rect 14004 657756 14056 657762
rect 14004 657698 14056 657704
rect 13820 654900 13872 654906
rect 13820 654842 13872 654848
rect 13726 355600 13782 355609
rect 13726 355535 13782 355544
rect 12440 328432 12492 328438
rect 12440 328374 12492 328380
rect 12452 328137 12480 328374
rect 12438 328128 12494 328137
rect 12438 328063 12494 328072
rect 13084 318844 13136 318850
rect 13084 318786 13136 318792
rect 12440 315988 12492 315994
rect 12440 315930 12492 315936
rect 12452 315489 12480 315930
rect 12438 315480 12494 315489
rect 12438 315415 12494 315424
rect 12440 302184 12492 302190
rect 12440 302126 12492 302132
rect 12452 301889 12480 302126
rect 12438 301880 12494 301889
rect 12438 301815 12494 301824
rect 12440 288380 12492 288386
rect 12440 288322 12492 288328
rect 12452 288153 12480 288322
rect 12438 288144 12494 288153
rect 12438 288079 12494 288088
rect 12440 276004 12492 276010
rect 12440 275946 12492 275952
rect 12452 275505 12480 275946
rect 12438 275496 12494 275505
rect 12438 275431 12494 275440
rect 12440 262200 12492 262206
rect 12440 262142 12492 262148
rect 12452 261905 12480 262142
rect 12438 261896 12494 261905
rect 12438 261831 12494 261840
rect 12440 248396 12492 248402
rect 12440 248338 12492 248344
rect 12452 248169 12480 248338
rect 12438 248160 12494 248169
rect 12438 248095 12494 248104
rect 12440 128308 12492 128314
rect 12440 128250 12492 128256
rect 12452 128217 12480 128250
rect 12438 128208 12494 128217
rect 12438 128143 12494 128152
rect 12440 115932 12492 115938
rect 12440 115874 12492 115880
rect 12452 115569 12480 115874
rect 12438 115560 12494 115569
rect 12438 115495 12494 115504
rect 12440 89684 12492 89690
rect 12440 89626 12492 89632
rect 12452 88913 12480 89626
rect 12438 88904 12494 88913
rect 12438 88839 12494 88848
rect 12440 75880 12492 75886
rect 12440 75822 12492 75828
rect 12452 75449 12480 75822
rect 12438 75440 12494 75449
rect 12438 75375 12494 75384
rect 12808 62076 12860 62082
rect 12808 62018 12860 62024
rect 12820 61985 12848 62018
rect 12806 61976 12862 61985
rect 12806 61911 12862 61920
rect 11886 48920 11942 48929
rect 11886 48855 11942 48864
rect 13096 35465 13124 318786
rect 13832 141953 13860 654842
rect 13912 654832 13964 654838
rect 13912 654774 13964 654780
rect 13924 155553 13952 654774
rect 14016 168201 14044 657698
rect 14188 657688 14240 657694
rect 14188 657630 14240 657636
rect 14096 656192 14148 656198
rect 14096 656134 14148 656140
rect 14108 182073 14136 656134
rect 14200 195537 14228 657630
rect 14292 622169 14320 659058
rect 14372 659048 14424 659054
rect 14372 658990 14424 658996
rect 14384 635497 14412 658990
rect 14464 658980 14516 658986
rect 14464 658922 14516 658928
rect 14476 648553 14504 658922
rect 20628 657620 20680 657626
rect 20628 657562 20680 657568
rect 20640 654922 20668 657562
rect 21376 656334 21404 700266
rect 31392 657552 31444 657558
rect 31392 657494 31444 657500
rect 21364 656328 21416 656334
rect 21364 656270 21416 656276
rect 31404 654922 31432 657494
rect 20378 654894 20668 654922
rect 31142 654894 31432 654922
rect 40052 654906 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 703050 73016 703520
rect 71780 703044 71832 703050
rect 71780 702986 71832 702992
rect 72976 703044 73028 703050
rect 72976 702986 73028 702992
rect 41512 670744 41564 670750
rect 41512 670686 41564 670692
rect 41524 654922 41552 670686
rect 71792 656266 71820 702986
rect 89180 700806 89208 703520
rect 89168 700800 89220 700806
rect 89168 700742 89220 700748
rect 96528 656940 96580 656946
rect 96528 656882 96580 656888
rect 71780 656260 71832 656266
rect 71780 656202 71832 656208
rect 85488 655784 85540 655790
rect 85488 655726 85540 655732
rect 74356 655716 74408 655722
rect 74356 655658 74408 655664
rect 63960 655648 64012 655654
rect 63960 655590 64012 655596
rect 53104 655580 53156 655586
rect 53104 655522 53156 655528
rect 53116 654922 53144 655522
rect 63972 654922 64000 655590
rect 40040 654900 40092 654906
rect 41524 654894 41998 654922
rect 52854 654894 53144 654922
rect 63710 654894 64000 654922
rect 74368 654922 74396 655658
rect 85500 654922 85528 655726
rect 96540 654922 96568 656882
rect 74368 654894 74474 654922
rect 85330 654894 85528 654922
rect 96186 654894 96568 654922
rect 40040 654842 40092 654848
rect 104912 654838 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 137848 700738 137876 703520
rect 137836 700732 137888 700738
rect 137836 700674 137888 700680
rect 154132 700534 154160 703520
rect 170324 702434 170352 703520
rect 169772 702406 170352 702434
rect 154120 700528 154172 700534
rect 154120 700470 154172 700476
rect 169772 657762 169800 702406
rect 193220 700528 193272 700534
rect 193220 700470 193272 700476
rect 193232 673454 193260 700470
rect 202800 700398 202828 703520
rect 218992 700670 219020 703520
rect 218980 700664 219032 700670
rect 218980 700606 219032 700612
rect 202788 700392 202840 700398
rect 202788 700334 202840 700340
rect 204260 700392 204312 700398
rect 204260 700334 204312 700340
rect 193232 673426 193352 673454
rect 169760 657756 169812 657762
rect 169760 657698 169812 657704
rect 118056 657280 118108 657286
rect 118056 657222 118108 657228
rect 118068 654922 118096 657222
rect 128912 657008 128964 657014
rect 128912 656950 128964 656956
rect 139766 656976 139822 656985
rect 128924 654922 128952 656950
rect 139766 656911 139822 656920
rect 139780 654922 139808 656911
rect 183192 656056 183244 656062
rect 183192 655998 183244 656004
rect 172336 655988 172388 655994
rect 172336 655930 172388 655936
rect 161296 655920 161348 655926
rect 161296 655862 161348 655868
rect 150256 655852 150308 655858
rect 150256 655794 150308 655800
rect 117806 654894 118096 654922
rect 128662 654894 128952 654922
rect 139518 654894 139808 654922
rect 150268 654922 150296 655794
rect 161308 654922 161336 655862
rect 172348 654922 172376 655930
rect 183204 654922 183232 655998
rect 150268 654894 150374 654922
rect 161138 654894 161336 654922
rect 171994 654894 172376 654922
rect 182850 654894 183232 654922
rect 193324 654922 193352 673426
rect 204272 654922 204300 700334
rect 215300 683188 215352 683194
rect 215300 683130 215352 683136
rect 215312 673454 215340 683130
rect 215312 673426 215432 673454
rect 215404 654922 215432 673426
rect 234632 656198 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 697610 267688 703520
rect 283852 700602 283880 703520
rect 283840 700596 283892 700602
rect 283840 700538 283892 700544
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 266372 659122 266400 697546
rect 266360 659116 266412 659122
rect 266360 659058 266412 659064
rect 237288 657756 237340 657762
rect 237288 657698 237340 657704
rect 234620 656192 234672 656198
rect 234620 656134 234672 656140
rect 237300 654922 237328 657698
rect 299492 657694 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 330484 700596 330536 700602
rect 330484 700538 330536 700544
rect 299480 657688 299532 657694
rect 299480 657630 299532 657636
rect 330496 657626 330524 700538
rect 331232 659054 331260 702986
rect 348804 700466 348832 703520
rect 364996 700505 365024 703520
rect 365720 700732 365772 700738
rect 365720 700674 365772 700680
rect 364982 700496 365038 700505
rect 348792 700460 348844 700466
rect 364982 700431 365038 700440
rect 348792 700402 348844 700408
rect 365732 673454 365760 700674
rect 376760 700664 376812 700670
rect 376760 700606 376812 700612
rect 376772 673454 376800 700606
rect 387800 696992 387852 696998
rect 387800 696934 387852 696940
rect 387812 673454 387840 696934
rect 365732 673426 366680 673454
rect 376772 673426 377352 673454
rect 387812 673426 388208 673454
rect 331220 659048 331272 659054
rect 331220 658990 331272 658996
rect 330484 657620 330536 657626
rect 330484 657562 330536 657568
rect 302148 657416 302200 657422
rect 302148 657358 302200 657364
rect 291016 657348 291068 657354
rect 291016 657290 291068 657296
rect 280712 657212 280764 657218
rect 280712 657154 280764 657160
rect 269856 657144 269908 657150
rect 269856 657086 269908 657092
rect 248052 657076 248104 657082
rect 248052 657018 248104 657024
rect 248064 654922 248092 657018
rect 269868 654922 269896 657086
rect 280724 654922 280752 657154
rect 193324 654894 193706 654922
rect 204272 654894 204470 654922
rect 215326 654894 215432 654922
rect 237038 654894 237328 654922
rect 247802 654894 248092 654922
rect 269514 654894 269896 654922
rect 280370 654894 280752 654922
rect 291028 654922 291056 657290
rect 302160 654922 302188 657358
rect 365628 657280 365680 657286
rect 365628 657222 365680 657228
rect 365640 656198 365668 657222
rect 365628 656192 365680 656198
rect 365628 656134 365680 656140
rect 291028 654894 291134 654922
rect 301990 654894 302188 654922
rect 366652 654922 366680 673426
rect 377324 654922 377352 673426
rect 388180 654922 388208 673426
rect 397472 658986 397500 703520
rect 398104 700460 398156 700466
rect 398104 700402 398156 700408
rect 397460 658980 397512 658986
rect 397460 658922 397512 658928
rect 398116 657558 398144 700402
rect 413664 700330 413692 703520
rect 429856 700369 429884 703520
rect 462332 700738 462360 703520
rect 462320 700732 462372 700738
rect 462320 700674 462372 700680
rect 478524 700534 478552 703520
rect 494808 700602 494836 703520
rect 527192 700670 527220 703520
rect 527180 700664 527232 700670
rect 527180 700606 527232 700612
rect 494796 700596 494848 700602
rect 494796 700538 494848 700544
rect 478512 700528 478564 700534
rect 478512 700470 478564 700476
rect 543476 700398 543504 703520
rect 559668 700466 559696 703520
rect 559656 700460 559708 700466
rect 559656 700402 559708 700408
rect 543464 700392 543516 700398
rect 429842 700360 429898 700369
rect 413652 700324 413704 700330
rect 543464 700334 543516 700340
rect 429842 700295 429898 700304
rect 413652 700266 413704 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 442908 657824 442960 657830
rect 442908 657766 442960 657772
rect 536564 657824 536616 657830
rect 536564 657766 536616 657772
rect 421472 657620 421524 657626
rect 421472 657562 421524 657568
rect 398104 657552 398156 657558
rect 398104 657494 398156 657500
rect 399760 657280 399812 657286
rect 399760 657222 399812 657228
rect 399772 654922 399800 657222
rect 410614 657112 410670 657121
rect 410614 657047 410670 657056
rect 410628 654922 410656 657047
rect 421484 654922 421512 657562
rect 430580 657008 430632 657014
rect 430580 656950 430632 656956
rect 432328 657008 432380 657014
rect 432328 656950 432380 656956
rect 430592 656266 430620 656950
rect 430580 656260 430632 656266
rect 430580 656202 430632 656208
rect 432340 654922 432368 656950
rect 442920 654922 442948 657766
rect 464988 657756 465040 657762
rect 464988 657698 465040 657704
rect 486424 657756 486476 657762
rect 486424 657698 486476 657704
rect 453856 657552 453908 657558
rect 453856 657494 453908 657500
rect 453868 654922 453896 657494
rect 464712 657484 464764 657490
rect 464712 657426 464764 657432
rect 453948 656940 454000 656946
rect 453948 656882 454000 656888
rect 453960 656334 453988 656882
rect 453948 656328 454000 656334
rect 453948 656270 454000 656276
rect 464724 654922 464752 657426
rect 366652 654894 367034 654922
rect 377324 654894 377798 654922
rect 388180 654894 388654 654922
rect 399510 654894 399800 654922
rect 410366 654894 410656 654922
rect 421130 654894 421512 654922
rect 431986 654894 432368 654922
rect 442842 654894 442948 654922
rect 453698 654894 453896 654922
rect 464462 654894 464752 654922
rect 465000 654838 465028 657698
rect 475568 657688 475620 657694
rect 475568 657630 475620 657636
rect 475580 654922 475608 657630
rect 486436 654922 486464 657698
rect 536288 657688 536340 657694
rect 536288 657630 536340 657636
rect 492588 657620 492640 657626
rect 492588 657562 492640 657568
rect 497280 657620 497332 657626
rect 497280 657562 497332 657568
rect 475318 654894 475608 654922
rect 486174 654894 486464 654922
rect 492600 654906 492628 657562
rect 497292 654922 497320 657562
rect 535000 657552 535052 657558
rect 535000 657494 535052 657500
rect 529848 656940 529900 656946
rect 529848 656882 529900 656888
rect 534724 656940 534776 656946
rect 534724 656882 534776 656888
rect 507676 656124 507728 656130
rect 507676 656066 507728 656072
rect 492588 654900 492640 654906
rect 497030 654894 497320 654922
rect 507688 654922 507716 656066
rect 529860 654922 529888 656882
rect 507688 654894 507794 654922
rect 529506 654894 529888 654922
rect 492588 654842 492640 654848
rect 104900 654832 104952 654838
rect 104900 654774 104952 654780
rect 464988 654832 465040 654838
rect 464988 654774 465040 654780
rect 520372 654764 520424 654770
rect 520372 654706 520424 654712
rect 107384 654696 107436 654702
rect 107042 654644 107384 654650
rect 520188 654696 520240 654702
rect 516782 654664 516838 654673
rect 107042 654638 107436 654644
rect 107042 654622 107424 654638
rect 356178 654634 356560 654650
rect 356178 654628 356572 654634
rect 356178 654622 356520 654628
rect 520384 654650 520412 654706
rect 520240 654644 520412 654650
rect 520188 654638 520412 654644
rect 516782 654599 516784 654608
rect 356520 654570 356572 654576
rect 516836 654599 516838 654608
rect 518164 654628 518216 654634
rect 516784 654570 516836 654576
rect 520200 654622 520412 654638
rect 521474 654664 521530 654673
rect 521530 654634 521654 654650
rect 521530 654628 521666 654634
rect 521530 654622 521614 654628
rect 521474 654599 521530 654608
rect 518164 654570 518216 654576
rect 521614 654570 521666 654576
rect 345664 654560 345716 654566
rect 334466 654498 334848 654514
rect 345322 654508 345664 654514
rect 345322 654502 345716 654508
rect 515218 654528 515274 654537
rect 334466 654492 334860 654498
rect 334466 654486 334808 654492
rect 345322 654486 345704 654502
rect 515218 654463 515220 654472
rect 334808 654434 334860 654440
rect 515272 654463 515274 654472
rect 515220 654434 515272 654440
rect 518176 654430 518204 654570
rect 520188 654560 520240 654566
rect 520372 654560 520424 654566
rect 520240 654508 520372 654514
rect 520188 654502 520424 654508
rect 521474 654528 521530 654537
rect 520200 654486 520412 654502
rect 521530 654498 521654 654514
rect 521530 654492 521666 654498
rect 521530 654486 521614 654492
rect 521474 654463 521530 654472
rect 521614 654434 521666 654440
rect 226248 654424 226300 654430
rect 226182 654372 226248 654378
rect 259000 654424 259052 654430
rect 226182 654366 226300 654372
rect 258658 654372 259000 654378
rect 313096 654424 313148 654430
rect 258658 654366 259052 654372
rect 312846 654372 313096 654378
rect 323952 654424 324004 654430
rect 312846 654366 313148 654372
rect 323702 654372 323952 654378
rect 518072 654424 518124 654430
rect 323702 654366 324004 654372
rect 518070 654392 518072 654401
rect 518164 654424 518216 654430
rect 518124 654392 518126 654401
rect 226182 654350 226288 654366
rect 258658 654350 259040 654366
rect 312846 654350 313136 654366
rect 323702 654350 323992 654366
rect 518716 654424 518768 654430
rect 518164 654366 518216 654372
rect 518650 654372 518716 654378
rect 520740 654424 520792 654430
rect 518650 654366 518768 654372
rect 520738 654392 520740 654401
rect 520792 654392 520794 654401
rect 518650 654350 518756 654366
rect 518070 654327 518126 654336
rect 520738 654327 520794 654336
rect 14462 648544 14518 648553
rect 14462 648479 14518 648488
rect 14370 635488 14426 635497
rect 14370 635423 14426 635432
rect 14278 622160 14334 622169
rect 14278 622095 14334 622104
rect 14186 195528 14242 195537
rect 14186 195463 14242 195472
rect 14094 182064 14150 182073
rect 14094 181999 14150 182008
rect 14002 168192 14058 168201
rect 14002 168127 14058 168136
rect 13910 155544 13966 155553
rect 13910 155479 13966 155488
rect 13818 141944 13874 141953
rect 13818 141879 13874 141888
rect 534736 73166 534764 656882
rect 534908 656124 534960 656130
rect 534908 656066 534960 656072
rect 534816 654152 534868 654158
rect 534816 654094 534868 654100
rect 534828 113150 534856 654094
rect 534920 153202 534948 656066
rect 535012 379506 535040 657494
rect 536196 657416 536248 657422
rect 536196 657358 536248 657364
rect 535276 657280 535328 657286
rect 535276 657222 535328 657228
rect 535092 657008 535144 657014
rect 535092 656950 535144 656956
rect 535182 656976 535238 656985
rect 535104 485790 535132 656950
rect 535182 656911 535238 656920
rect 535196 607918 535224 656911
rect 535288 644434 535316 657222
rect 536104 654628 536156 654634
rect 536104 654570 536156 654576
rect 535276 644428 535328 644434
rect 535276 644370 535328 644376
rect 535184 607912 535236 607918
rect 535184 607854 535236 607860
rect 535092 485784 535144 485790
rect 535092 485726 535144 485732
rect 535000 379500 535052 379506
rect 535000 379442 535052 379448
rect 534908 153196 534960 153202
rect 534908 153138 534960 153144
rect 534816 113144 534868 113150
rect 534816 113086 534868 113092
rect 534724 73160 534776 73166
rect 534724 73102 534776 73108
rect 536116 60722 536144 654570
rect 536208 259418 536236 657358
rect 536300 273222 536328 657630
rect 536472 657484 536524 657490
rect 536472 657426 536524 657432
rect 536380 657348 536432 657354
rect 536380 657290 536432 657296
rect 536392 313274 536420 657290
rect 536484 325650 536512 657426
rect 536576 431934 536604 657766
rect 539232 657756 539284 657762
rect 539232 657698 539284 657704
rect 539140 657620 539192 657626
rect 539140 657562 539192 657568
rect 537484 656056 537536 656062
rect 537484 655998 537536 656004
rect 536656 654016 536708 654022
rect 536656 653958 536708 653964
rect 536668 632058 536696 653958
rect 536656 632052 536708 632058
rect 536656 631994 536708 632000
rect 536564 431928 536616 431934
rect 536564 431870 536616 431876
rect 536472 325644 536524 325650
rect 536472 325586 536524 325592
rect 536380 313268 536432 313274
rect 536380 313210 536432 313216
rect 536288 273216 536340 273222
rect 536288 273158 536340 273164
rect 536196 259412 536248 259418
rect 536196 259354 536248 259360
rect 536104 60716 536156 60722
rect 536104 60658 536156 60664
rect 537496 46918 537524 655998
rect 537668 655988 537720 655994
rect 537668 655930 537720 655936
rect 537574 635216 537630 635225
rect 537574 635151 537630 635160
rect 537484 46912 537536 46918
rect 537484 46854 537536 46860
rect 13082 35456 13138 35465
rect 13082 35391 13138 35400
rect 537588 33114 537616 635151
rect 537680 86970 537708 655930
rect 538956 655920 539008 655926
rect 538956 655862 539008 655868
rect 537760 655784 537812 655790
rect 537760 655726 537812 655732
rect 537772 458182 537800 655726
rect 537944 655716 537996 655722
rect 537944 655658 537996 655664
rect 537852 654696 537904 654702
rect 537852 654638 537904 654644
rect 537760 458176 537812 458182
rect 537760 458118 537812 458124
rect 537758 421152 537814 421161
rect 537758 421087 537814 421096
rect 537668 86964 537720 86970
rect 537668 86906 537720 86912
rect 537576 33108 537628 33114
rect 537576 33050 537628 33056
rect 13726 21176 13782 21185
rect 13726 21111 13782 21120
rect 13740 13802 13768 21111
rect 537772 20670 537800 421087
rect 537864 353258 537892 654638
rect 537956 511970 537984 655658
rect 538036 655648 538088 655654
rect 538036 655590 538088 655596
rect 538048 564398 538076 655590
rect 538128 655580 538180 655586
rect 538128 655522 538180 655528
rect 538140 618254 538168 655522
rect 538864 654560 538916 654566
rect 538864 654502 538916 654508
rect 538128 618248 538180 618254
rect 538128 618190 538180 618196
rect 538036 564392 538088 564398
rect 538036 564334 538088 564340
rect 537944 511964 537996 511970
rect 537944 511906 537996 511912
rect 537852 353252 537904 353258
rect 537852 353194 537904 353200
rect 537850 207768 537906 207777
rect 537850 207703 537906 207712
rect 537760 20664 537812 20670
rect 537760 20606 537812 20612
rect 52104 13802 52132 15028
rect 13728 13796 13780 13802
rect 13728 13738 13780 13744
rect 52092 13796 52144 13802
rect 52092 13738 52144 13744
rect 3700 13660 3752 13666
rect 3700 13602 3752 13608
rect 3608 13592 3660 13598
rect 3608 13534 3660 13540
rect 3424 13524 3476 13530
rect 3424 13466 3476 13472
rect 52104 13122 52132 13738
rect 126348 13530 126376 15028
rect 200592 13598 200620 15028
rect 349172 13666 349200 15028
rect 423508 13734 423536 15028
rect 423496 13728 423548 13734
rect 423496 13670 423548 13676
rect 349160 13660 349212 13666
rect 349160 13602 349212 13608
rect 200580 13592 200632 13598
rect 200580 13534 200632 13540
rect 126336 13524 126388 13530
rect 126336 13466 126388 13472
rect 52092 13116 52144 13122
rect 52092 13058 52144 13064
rect 537864 6866 537892 207703
rect 538876 100706 538904 654502
rect 538968 126954 538996 655862
rect 539048 655852 539100 655858
rect 539048 655794 539100 655800
rect 539060 167006 539088 655794
rect 539152 193186 539180 657562
rect 539244 233238 539272 657698
rect 540244 657212 540296 657218
rect 540244 657154 540296 657160
rect 539324 654288 539376 654294
rect 539324 654230 539376 654236
rect 539336 471986 539364 654230
rect 539324 471980 539376 471986
rect 539324 471922 539376 471928
rect 540256 365702 540284 657154
rect 540336 657144 540388 657150
rect 540336 657086 540388 657092
rect 540348 419490 540376 657086
rect 540428 657076 540480 657082
rect 540428 657018 540480 657024
rect 540440 525774 540468 657018
rect 580816 656328 580868 656334
rect 580816 656270 580868 656276
rect 580540 656260 580592 656266
rect 580540 656202 580592 656208
rect 580172 654832 580224 654838
rect 580172 654774 580224 654780
rect 580078 653440 580134 653449
rect 580078 653375 580134 653384
rect 579988 644428 580040 644434
rect 579988 644370 580040 644376
rect 580000 644065 580028 644370
rect 579986 644056 580042 644065
rect 579986 643991 580042 644000
rect 579988 632052 580040 632058
rect 579988 631994 580040 632000
rect 580000 630873 580028 631994
rect 579986 630864 580042 630873
rect 579986 630799 580042 630808
rect 579988 618248 580040 618254
rect 579988 618190 580040 618196
rect 580000 617545 580028 618190
rect 579986 617536 580042 617545
rect 579986 617471 580042 617480
rect 580092 591025 580120 653375
rect 580078 591016 580134 591025
rect 580078 590951 580134 590960
rect 580184 577697 580212 654774
rect 580264 654492 580316 654498
rect 580264 654434 580316 654440
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580172 564392 580224 564398
rect 580170 564360 580172 564369
rect 580224 564360 580226 564369
rect 580170 564295 580226 564304
rect 540428 525768 540480 525774
rect 540428 525710 540480 525716
rect 580172 525768 580224 525774
rect 580172 525710 580224 525716
rect 580184 524521 580212 525710
rect 580170 524512 580226 524521
rect 580170 524447 580226 524456
rect 580172 511964 580224 511970
rect 580172 511906 580224 511912
rect 580184 511329 580212 511906
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580172 485784 580224 485790
rect 580172 485726 580224 485732
rect 580184 484673 580212 485726
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 579804 471980 579856 471986
rect 579804 471922 579856 471928
rect 579816 471481 579844 471922
rect 579802 471472 579858 471481
rect 579802 471407 579858 471416
rect 580172 458176 580224 458182
rect 580170 458144 580172 458153
rect 580224 458144 580226 458153
rect 580170 458079 580226 458088
rect 580172 431928 580224 431934
rect 580172 431870 580224 431876
rect 580184 431633 580212 431870
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 540336 419484 540388 419490
rect 540336 419426 540388 419432
rect 580172 419484 580224 419490
rect 580172 419426 580224 419432
rect 580184 418305 580212 419426
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 540244 365696 540296 365702
rect 540244 365638 540296 365644
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 579620 353252 579672 353258
rect 579620 353194 579672 353200
rect 579632 351937 579660 353194
rect 579618 351928 579674 351937
rect 579618 351863 579674 351872
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 579804 259412 579856 259418
rect 579804 259354 579856 259360
rect 579816 258913 579844 259354
rect 579802 258904 579858 258913
rect 579802 258839 579858 258848
rect 539232 233232 539284 233238
rect 539232 233174 539284 233180
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 539140 193180 539192 193186
rect 539140 193122 539192 193128
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 539048 167000 539100 167006
rect 539048 166942 539100 166948
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 579804 153196 579856 153202
rect 579804 153138 579856 153144
rect 579816 152697 579844 153138
rect 579802 152688 579858 152697
rect 579802 152623 579858 152632
rect 580276 139369 580304 654434
rect 580356 654424 580408 654430
rect 580356 654366 580408 654372
rect 580368 179217 580396 654366
rect 580448 654356 580500 654362
rect 580448 654298 580500 654304
rect 580460 219065 580488 654298
rect 580552 245585 580580 656202
rect 580724 656192 580776 656198
rect 580724 656134 580776 656140
rect 580632 607912 580684 607918
rect 580632 607854 580684 607860
rect 580538 245576 580594 245585
rect 580538 245511 580594 245520
rect 580446 219056 580502 219065
rect 580446 218991 580502 219000
rect 580644 205737 580672 607854
rect 580736 298761 580764 656134
rect 580828 404977 580856 656270
rect 580908 654900 580960 654906
rect 580908 654842 580960 654848
rect 580920 537849 580948 654842
rect 580906 537840 580962 537849
rect 580906 537775 580962 537784
rect 580814 404968 580870 404977
rect 580814 404903 580870 404912
rect 580722 298752 580778 298761
rect 580722 298687 580778 298696
rect 580630 205728 580686 205737
rect 580630 205663 580686 205672
rect 580354 179208 580410 179217
rect 580354 179143 580410 179152
rect 580262 139360 580318 139369
rect 580262 139295 580318 139304
rect 538956 126948 539008 126954
rect 538956 126890 539008 126896
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 538864 100700 538916 100706
rect 538864 100642 538916 100648
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 579620 13116 579672 13122
rect 579620 13058 579672 13064
rect 537852 6860 537904 6866
rect 537852 6802 537904 6808
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579632 354 579660 13058
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 579774 354 579886 480
rect 579632 326 579886 354
rect 579774 -960 579886 326
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 2778 684256 2834 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3422 619112 3478 619168
rect 2962 527856 3018 527912
rect 3238 501744 3294 501800
rect 2778 475652 2834 475688
rect 2778 475632 2780 475652
rect 2780 475632 2832 475652
rect 2832 475632 2834 475652
rect 3330 449556 3332 449576
rect 3332 449556 3384 449576
rect 3384 449556 3386 449576
rect 3330 449520 3386 449556
rect 3330 423544 3386 423600
rect 3238 410488 3294 410544
rect 3238 397432 3294 397488
rect 3330 371320 3386 371376
rect 2962 345344 3018 345400
rect 3606 606056 3662 606112
rect 3514 579944 3570 580000
rect 3514 566888 3570 566944
rect 3422 319232 3478 319288
rect 3698 553832 3754 553888
rect 3606 514800 3662 514856
rect 3422 306176 3478 306232
rect 3330 293120 3386 293176
rect 3698 462576 3754 462632
rect 3790 358400 3846 358456
rect 3422 214920 3478 214976
rect 3514 162832 3570 162888
rect 3606 110608 3662 110664
rect 3698 71576 3754 71632
rect 12990 608504 13046 608560
rect 13082 595448 13138 595504
rect 12898 582120 12954 582176
rect 12438 568540 12494 568576
rect 12438 568520 12440 568540
rect 12440 568520 12492 568540
rect 12492 568520 12494 568540
rect 11886 555464 11942 555520
rect 12438 542000 12494 542056
rect 12438 528128 12494 528184
rect 12438 514820 12494 514856
rect 12438 514800 12440 514820
rect 12440 514800 12492 514820
rect 12492 514800 12494 514820
rect 12438 501064 12494 501120
rect 12438 487736 12494 487792
rect 12438 474816 12494 474872
rect 12438 461352 12494 461408
rect 13174 435512 13230 435568
rect 13266 421912 13322 421968
rect 13358 408176 13414 408232
rect 13450 395528 13506 395584
rect 13542 382200 13598 382256
rect 11794 342080 11850 342136
rect 11702 102040 11758 102096
rect 13634 368192 13690 368248
rect 13726 355544 13782 355600
rect 12438 328072 12494 328128
rect 12438 315424 12494 315480
rect 12438 301824 12494 301880
rect 12438 288088 12494 288144
rect 12438 275440 12494 275496
rect 12438 261840 12494 261896
rect 12438 248104 12494 248160
rect 12438 128152 12494 128208
rect 12438 115504 12494 115560
rect 12438 88848 12494 88904
rect 12438 75384 12494 75440
rect 12806 61920 12862 61976
rect 11886 48864 11942 48920
rect 139766 656920 139822 656976
rect 364982 700440 365038 700496
rect 429842 700304 429898 700360
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 410614 657056 410670 657112
rect 516782 654628 516838 654664
rect 516782 654608 516784 654628
rect 516784 654608 516836 654628
rect 516836 654608 516838 654628
rect 521474 654608 521530 654664
rect 515218 654492 515274 654528
rect 515218 654472 515220 654492
rect 515220 654472 515272 654492
rect 515272 654472 515274 654492
rect 521474 654472 521530 654528
rect 518070 654372 518072 654392
rect 518072 654372 518124 654392
rect 518124 654372 518126 654392
rect 518070 654336 518126 654372
rect 520738 654372 520740 654392
rect 520740 654372 520792 654392
rect 520792 654372 520794 654392
rect 520738 654336 520794 654372
rect 14462 648488 14518 648544
rect 14370 635432 14426 635488
rect 14278 622104 14334 622160
rect 14186 195472 14242 195528
rect 14094 182008 14150 182064
rect 14002 168136 14058 168192
rect 13910 155488 13966 155544
rect 13818 141888 13874 141944
rect 535182 656920 535238 656976
rect 537574 635160 537630 635216
rect 13082 35400 13138 35456
rect 537758 421096 537814 421152
rect 13726 21120 13782 21176
rect 537850 207712 537906 207768
rect 580078 653384 580134 653440
rect 579986 644000 580042 644056
rect 579986 630808 580042 630864
rect 579986 617480 580042 617536
rect 580078 590960 580134 591016
rect 580170 577632 580226 577688
rect 580170 564340 580172 564360
rect 580172 564340 580224 564360
rect 580224 564340 580226 564360
rect 580170 564304 580226 564340
rect 580170 524456 580226 524512
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579802 471416 579858 471472
rect 580170 458124 580172 458144
rect 580172 458124 580224 458144
rect 580224 458124 580226 458144
rect 580170 458088 580226 458124
rect 580170 431568 580226 431624
rect 580170 418240 580226 418296
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 579618 351872 579674 351928
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580170 272176 580226 272232
rect 579802 258848 579858 258904
rect 579986 232328 580042 232384
rect 580170 192480 580226 192536
rect 580170 165824 580226 165880
rect 579802 152632 579858 152688
rect 580538 245520 580594 245576
rect 580446 219000 580502 219056
rect 580906 537784 580962 537840
rect 580814 404912 580870 404968
rect 580722 298696 580778 298752
rect 580630 205672 580686 205728
rect 580354 179152 580410 179208
rect 580262 139304 580318 139360
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect 13670 700436 13676 700500
rect 13740 700498 13746 700500
rect 364977 700498 365043 700501
rect 13740 700496 365043 700498
rect 13740 700440 364982 700496
rect 365038 700440 365043 700496
rect 13740 700438 365043 700440
rect 13740 700436 13746 700438
rect 364977 700435 365043 700438
rect 12750 700300 12756 700364
rect 12820 700362 12826 700364
rect 429837 700362 429903 700365
rect 12820 700360 429903 700362
rect 12820 700304 429842 700360
rect 429898 700304 429903 700360
rect 12820 700302 429903 700304
rect 12820 700300 12826 700302
rect 429837 700299 429903 700302
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 2773 684314 2839 684317
rect -960 684312 2839 684314
rect -960 684256 2778 684312
rect 2834 684256 2839 684312
rect -960 684254 2839 684256
rect -960 684164 480 684254
rect 2773 684251 2839 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect 410609 657114 410675 657117
rect 469622 657114 469628 657116
rect 410609 657112 469628 657114
rect 410609 657056 410614 657112
rect 410670 657056 469628 657112
rect 410609 657054 469628 657056
rect 410609 657051 410675 657054
rect 469622 657052 469628 657054
rect 469692 657052 469698 657116
rect 139761 656978 139827 656981
rect 535177 656978 535243 656981
rect 139761 656976 535243 656978
rect 139761 656920 139766 656976
rect 139822 656920 535182 656976
rect 535238 656920 535243 656976
rect 139761 656918 535243 656920
rect 139761 656915 139827 656918
rect 535177 656915 535243 656918
rect 516777 654666 516843 654669
rect 521469 654666 521535 654669
rect 516777 654664 521535 654666
rect 516777 654608 516782 654664
rect 516838 654608 521474 654664
rect 521530 654608 521535 654664
rect 516777 654606 521535 654608
rect 516777 654603 516843 654606
rect 521469 654603 521535 654606
rect 515213 654530 515279 654533
rect 521469 654530 521535 654533
rect 515213 654528 521535 654530
rect 515213 654472 515218 654528
rect 515274 654472 521474 654528
rect 521530 654472 521535 654528
rect 515213 654470 521535 654472
rect 515213 654467 515279 654470
rect 521469 654467 521535 654470
rect 518065 654394 518131 654397
rect 520733 654394 520799 654397
rect 518065 654392 520799 654394
rect 518065 654336 518070 654392
rect 518126 654336 520738 654392
rect 520794 654336 520799 654392
rect 518065 654334 520799 654336
rect 518065 654331 518131 654334
rect 520733 654331 520799 654334
rect 469622 653380 469628 653444
rect 469692 653442 469698 653444
rect 580073 653442 580139 653445
rect 469692 653440 580139 653442
rect 469692 653384 580078 653440
rect 580134 653384 580139 653440
rect 469692 653382 580139 653384
rect 469692 653380 469698 653382
rect 580073 653379 580139 653382
rect 14457 648546 14523 648549
rect 14457 648544 15210 648546
rect 14457 648488 14462 648544
rect 14518 648488 15210 648544
rect 14457 648486 15210 648488
rect 14457 648483 14523 648486
rect 15150 648244 15210 648486
rect -960 644996 480 645236
rect 579981 644058 580047 644061
rect 583520 644058 584960 644148
rect 579981 644056 584960 644058
rect 579981 644000 579986 644056
rect 580042 644000 584960 644056
rect 579981 643998 584960 644000
rect 579981 643995 580047 643998
rect 583520 643908 584960 643998
rect 14365 635490 14431 635493
rect 14365 635488 15210 635490
rect 14365 635432 14370 635488
rect 14426 635432 15210 635488
rect 14365 635430 15210 635432
rect 14365 635427 14431 635430
rect 15150 634916 15210 635430
rect 537569 635218 537635 635221
rect 534582 635216 537635 635218
rect 534582 635160 537574 635216
rect 537630 635160 537635 635216
rect 534582 635158 537635 635160
rect 534582 634916 534642 635158
rect 537569 635155 537635 635158
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 579981 630866 580047 630869
rect 583520 630866 584960 630956
rect 579981 630864 584960 630866
rect 579981 630808 579986 630864
rect 580042 630808 584960 630864
rect 579981 630806 584960 630808
rect 579981 630803 580047 630806
rect 583520 630716 584960 630806
rect 14273 622162 14339 622165
rect 14273 622160 15210 622162
rect 14273 622104 14278 622160
rect 14334 622104 15210 622160
rect 14273 622102 15210 622104
rect 14273 622099 14339 622102
rect 15150 621588 15210 622102
rect -960 619170 480 619260
rect 3417 619170 3483 619173
rect -960 619168 3483 619170
rect -960 619112 3422 619168
rect 3478 619112 3483 619168
rect -960 619110 3483 619112
rect -960 619020 480 619110
rect 3417 619107 3483 619110
rect 579981 617538 580047 617541
rect 583520 617538 584960 617628
rect 579981 617536 584960 617538
rect 579981 617480 579986 617536
rect 580042 617480 584960 617536
rect 579981 617478 584960 617480
rect 579981 617475 580047 617478
rect 583520 617388 584960 617478
rect 12985 608562 13051 608565
rect 12985 608560 15210 608562
rect 12985 608504 12990 608560
rect 13046 608504 15210 608560
rect 12985 608502 15210 608504
rect 12985 608499 13051 608502
rect 15150 608260 15210 608502
rect -960 606114 480 606204
rect 3601 606114 3667 606117
rect -960 606112 3667 606114
rect -960 606056 3606 606112
rect 3662 606056 3667 606112
rect -960 606054 3667 606056
rect -960 605964 480 606054
rect 3601 606051 3667 606054
rect 583520 604060 584960 604300
rect 13077 595506 13143 595509
rect 13077 595504 15210 595506
rect 13077 595448 13082 595504
rect 13138 595448 15210 595504
rect 13077 595446 15210 595448
rect 13077 595443 13143 595446
rect 15150 594932 15210 595446
rect -960 592908 480 593148
rect 580073 591018 580139 591021
rect 583520 591018 584960 591108
rect 580073 591016 584960 591018
rect 580073 590960 580078 591016
rect 580134 590960 584960 591016
rect 580073 590958 584960 590960
rect 580073 590955 580139 590958
rect 583520 590868 584960 590958
rect 12893 582178 12959 582181
rect 12893 582176 15210 582178
rect 12893 582120 12898 582176
rect 12954 582120 15210 582176
rect 12893 582118 15210 582120
rect 12893 582115 12959 582118
rect 15150 581604 15210 582118
rect -960 580002 480 580092
rect 3509 580002 3575 580005
rect -960 580000 3575 580002
rect -960 579944 3514 580000
rect 3570 579944 3575 580000
rect -960 579942 3575 579944
rect -960 579852 480 579942
rect 3509 579939 3575 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect 12433 568578 12499 568581
rect 12433 568576 15394 568578
rect 12433 568520 12438 568576
rect 12494 568520 15394 568576
rect 12433 568518 15394 568520
rect 12433 568515 12499 568518
rect 15334 568276 15394 568518
rect -960 566946 480 567036
rect 3509 566946 3575 566949
rect -960 566944 3575 566946
rect -960 566888 3514 566944
rect 3570 566888 3575 566944
rect -960 566886 3575 566888
rect -960 566796 480 566886
rect 3509 566883 3575 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect 11881 555522 11947 555525
rect 11881 555520 15210 555522
rect 11881 555464 11886 555520
rect 11942 555464 15210 555520
rect 11881 555462 15210 555464
rect 11881 555459 11947 555462
rect 15150 554948 15210 555462
rect -960 553890 480 553980
rect 3693 553890 3759 553893
rect -960 553888 3759 553890
rect -960 553832 3698 553888
rect 3754 553832 3759 553888
rect -960 553830 3759 553832
rect -960 553740 480 553830
rect 3693 553827 3759 553830
rect 583520 551020 584960 551260
rect 12433 542058 12499 542061
rect 12433 542056 15210 542058
rect 12433 542000 12438 542056
rect 12494 542000 15210 542056
rect 12433 541998 15210 542000
rect 12433 541995 12499 541998
rect 15150 541620 15210 541998
rect -960 540684 480 540924
rect 580901 537842 580967 537845
rect 583520 537842 584960 537932
rect 580901 537840 584960 537842
rect 580901 537784 580906 537840
rect 580962 537784 584960 537840
rect 580901 537782 584960 537784
rect 580901 537779 580967 537782
rect 583520 537692 584960 537782
rect 12433 528186 12499 528189
rect 15150 528186 15210 528292
rect 12433 528184 15210 528186
rect 12433 528128 12438 528184
rect 12494 528128 15210 528184
rect 12433 528126 15210 528128
rect 12433 528123 12499 528126
rect -960 527914 480 528004
rect 2957 527914 3023 527917
rect -960 527912 3023 527914
rect -960 527856 2962 527912
rect 3018 527856 3023 527912
rect -960 527854 3023 527856
rect -960 527764 480 527854
rect 2957 527851 3023 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3601 514858 3667 514861
rect -960 514856 3667 514858
rect -960 514800 3606 514856
rect 3662 514800 3667 514856
rect -960 514798 3667 514800
rect -960 514708 480 514798
rect 3601 514795 3667 514798
rect 12433 514858 12499 514861
rect 15150 514858 15210 514964
rect 12433 514856 15210 514858
rect 12433 514800 12438 514856
rect 12494 514800 15210 514856
rect 12433 514798 15210 514800
rect 12433 514795 12499 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3233 501802 3299 501805
rect -960 501800 3299 501802
rect -960 501744 3238 501800
rect 3294 501744 3299 501800
rect -960 501742 3299 501744
rect -960 501652 480 501742
rect 3233 501739 3299 501742
rect 12433 501122 12499 501125
rect 15150 501122 15210 501636
rect 12433 501120 15210 501122
rect 12433 501064 12438 501120
rect 12494 501064 15210 501120
rect 12433 501062 15210 501064
rect 12433 501059 12499 501062
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 12433 487794 12499 487797
rect 15150 487794 15210 488308
rect 12433 487792 15210 487794
rect 12433 487736 12438 487792
rect 12494 487736 15210 487792
rect 12433 487734 15210 487736
rect 12433 487731 12499 487734
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 2773 475690 2839 475693
rect -960 475688 2839 475690
rect -960 475632 2778 475688
rect 2834 475632 2839 475688
rect -960 475630 2839 475632
rect -960 475540 480 475630
rect 2773 475627 2839 475630
rect 12433 474874 12499 474877
rect 15150 474874 15210 474980
rect 12433 474872 15210 474874
rect 12433 474816 12438 474872
rect 12494 474816 15210 474872
rect 12433 474814 15210 474816
rect 12433 474811 12499 474814
rect 579797 471474 579863 471477
rect 583520 471474 584960 471564
rect 579797 471472 584960 471474
rect 579797 471416 579802 471472
rect 579858 471416 584960 471472
rect 579797 471414 584960 471416
rect 579797 471411 579863 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3693 462634 3759 462637
rect -960 462632 3759 462634
rect -960 462576 3698 462632
rect 3754 462576 3759 462632
rect -960 462574 3759 462576
rect -960 462484 480 462574
rect 3693 462571 3759 462574
rect 12433 461410 12499 461413
rect 15150 461410 15210 461652
rect 12433 461408 15210 461410
rect 12433 461352 12438 461408
rect 12494 461352 15210 461408
rect 12433 461350 15210 461352
rect 12433 461347 12499 461350
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 13169 435570 13235 435573
rect 13169 435568 15210 435570
rect 13169 435512 13174 435568
rect 13230 435512 15210 435568
rect 13169 435510 15210 435512
rect 13169 435507 13235 435510
rect 15150 434996 15210 435510
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3325 423602 3391 423605
rect -960 423600 3391 423602
rect -960 423544 3330 423600
rect 3386 423544 3391 423600
rect -960 423542 3391 423544
rect -960 423452 480 423542
rect 3325 423539 3391 423542
rect 13261 421970 13327 421973
rect 13261 421968 15210 421970
rect 13261 421912 13266 421968
rect 13322 421912 15210 421968
rect 13261 421910 15210 421912
rect 13261 421907 13327 421910
rect 15150 421668 15210 421910
rect 534766 421154 534826 421668
rect 537753 421154 537819 421157
rect 534766 421152 537819 421154
rect 534766 421096 537758 421152
rect 537814 421096 537819 421152
rect 534766 421094 537819 421096
rect 537753 421091 537819 421094
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3233 410546 3299 410549
rect -960 410544 3299 410546
rect -960 410488 3238 410544
rect 3294 410488 3299 410544
rect -960 410486 3299 410488
rect -960 410396 480 410486
rect 3233 410483 3299 410486
rect 13353 408234 13419 408237
rect 15150 408234 15210 408340
rect 13353 408232 15210 408234
rect 13353 408176 13358 408232
rect 13414 408176 15210 408232
rect 13353 408174 15210 408176
rect 13353 408171 13419 408174
rect 580809 404970 580875 404973
rect 583520 404970 584960 405060
rect 580809 404968 584960 404970
rect 580809 404912 580814 404968
rect 580870 404912 584960 404968
rect 580809 404910 584960 404912
rect 580809 404907 580875 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3233 397490 3299 397493
rect -960 397488 3299 397490
rect -960 397432 3238 397488
rect 3294 397432 3299 397488
rect -960 397430 3299 397432
rect -960 397340 480 397430
rect 3233 397427 3299 397430
rect 13445 395586 13511 395589
rect 13445 395584 15210 395586
rect 13445 395528 13450 395584
rect 13506 395528 15210 395584
rect 13445 395526 15210 395528
rect 13445 395523 13511 395526
rect 15150 395012 15210 395526
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 13537 382258 13603 382261
rect 13537 382256 15210 382258
rect 13537 382200 13542 382256
rect 13598 382200 15210 382256
rect 13537 382198 15210 382200
rect 13537 382195 13603 382198
rect 15150 381684 15210 382198
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3325 371378 3391 371381
rect -960 371376 3391 371378
rect -960 371320 3330 371376
rect 3386 371320 3391 371376
rect -960 371318 3391 371320
rect -960 371228 480 371318
rect 3325 371315 3391 371318
rect 13629 368250 13695 368253
rect 15150 368250 15210 368356
rect 13629 368248 15210 368250
rect 13629 368192 13634 368248
rect 13690 368192 15210 368248
rect 13629 368190 15210 368192
rect 13629 368187 13695 368190
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3785 358458 3851 358461
rect -960 358456 3851 358458
rect -960 358400 3790 358456
rect 3846 358400 3851 358456
rect -960 358398 3851 358400
rect -960 358308 480 358398
rect 3785 358395 3851 358398
rect 13721 355602 13787 355605
rect 13721 355600 15210 355602
rect 13721 355544 13726 355600
rect 13782 355544 15210 355600
rect 13721 355542 15210 355544
rect 13721 355539 13787 355542
rect 15150 355028 15210 355542
rect 579613 351930 579679 351933
rect 583520 351930 584960 352020
rect 579613 351928 584960 351930
rect 579613 351872 579618 351928
rect 579674 351872 584960 351928
rect 579613 351870 584960 351872
rect 579613 351867 579679 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 2957 345402 3023 345405
rect -960 345400 3023 345402
rect -960 345344 2962 345400
rect 3018 345344 3023 345400
rect -960 345342 3023 345344
rect -960 345252 480 345342
rect 2957 345339 3023 345342
rect 11789 342138 11855 342141
rect 11789 342136 15210 342138
rect 11789 342080 11794 342136
rect 11850 342080 15210 342136
rect 11789 342078 15210 342080
rect 11789 342075 11855 342078
rect 15150 341700 15210 342078
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 12433 328130 12499 328133
rect 15150 328130 15210 328236
rect 12433 328128 15210 328130
rect 12433 328072 12438 328128
rect 12494 328072 15210 328128
rect 12433 328070 15210 328072
rect 12433 328067 12499 328070
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 12433 315482 12499 315485
rect 12433 315480 15210 315482
rect 12433 315424 12438 315480
rect 12494 315424 15210 315480
rect 12433 315422 15210 315424
rect 12433 315419 12499 315422
rect 15150 314908 15210 315422
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 12433 301882 12499 301885
rect 12433 301880 15210 301882
rect 12433 301824 12438 301880
rect 12494 301824 15210 301880
rect 12433 301822 15210 301824
rect 12433 301819 12499 301822
rect 15150 301580 15210 301822
rect 580717 298754 580783 298757
rect 583520 298754 584960 298844
rect 580717 298752 584960 298754
rect 580717 298696 580722 298752
rect 580778 298696 584960 298752
rect 580717 298694 584960 298696
rect 580717 298691 580783 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3325 293178 3391 293181
rect -960 293176 3391 293178
rect -960 293120 3330 293176
rect 3386 293120 3391 293176
rect -960 293118 3391 293120
rect -960 293028 480 293118
rect 3325 293115 3391 293118
rect 12433 288146 12499 288149
rect 15150 288146 15210 288252
rect 12433 288144 15210 288146
rect 12433 288088 12438 288144
rect 12494 288088 15210 288144
rect 12433 288086 15210 288088
rect 12433 288083 12499 288086
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 12433 275498 12499 275501
rect 12433 275496 15210 275498
rect 12433 275440 12438 275496
rect 12494 275440 15210 275496
rect 12433 275438 15210 275440
rect 12433 275435 12499 275438
rect 15150 274924 15210 275438
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267052 480 267292
rect 12433 261898 12499 261901
rect 12433 261896 15210 261898
rect 12433 261840 12438 261896
rect 12494 261840 15210 261896
rect 12433 261838 15210 261840
rect 12433 261835 12499 261838
rect 15150 261596 15210 261838
rect 579797 258906 579863 258909
rect 583520 258906 584960 258996
rect 579797 258904 584960 258906
rect 579797 258848 579802 258904
rect 579858 258848 584960 258904
rect 579797 258846 584960 258848
rect 579797 258843 579863 258846
rect 583520 258756 584960 258846
rect -960 253996 480 254236
rect 12433 248162 12499 248165
rect 15150 248162 15210 248268
rect 12433 248160 15210 248162
rect 12433 248104 12438 248160
rect 12494 248104 15210 248160
rect 12433 248102 15210 248104
rect 12433 248099 12499 248102
rect 580533 245578 580599 245581
rect 583520 245578 584960 245668
rect 580533 245576 584960 245578
rect 580533 245520 580538 245576
rect 580594 245520 584960 245576
rect 580533 245518 584960 245520
rect 580533 245515 580599 245518
rect 583520 245428 584960 245518
rect -960 240940 480 241180
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 12750 222124 12756 222188
rect 12820 222186 12826 222188
rect 12820 222126 15210 222186
rect 12820 222124 12826 222126
rect 15150 221612 15210 222126
rect 580441 219058 580507 219061
rect 583520 219058 584960 219148
rect 580441 219056 584960 219058
rect 580441 219000 580446 219056
rect 580502 219000 584960 219056
rect 580441 218998 584960 219000
rect 580441 218995 580507 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3417 214978 3483 214981
rect -960 214976 3483 214978
rect -960 214920 3422 214976
rect 3478 214920 3483 214976
rect -960 214918 3483 214920
rect -960 214828 480 214918
rect 3417 214915 3483 214918
rect 13670 208116 13676 208180
rect 13740 208178 13746 208180
rect 15150 208178 15210 208284
rect 13740 208118 15210 208178
rect 13740 208116 13746 208118
rect 534766 207770 534826 208284
rect 537845 207770 537911 207773
rect 534766 207768 537911 207770
rect 534766 207712 537850 207768
rect 537906 207712 537911 207768
rect 534766 207710 537911 207712
rect 537845 207707 537911 207710
rect 580625 205730 580691 205733
rect 583520 205730 584960 205820
rect 580625 205728 584960 205730
rect 580625 205672 580630 205728
rect 580686 205672 584960 205728
rect 580625 205670 584960 205672
rect 580625 205667 580691 205670
rect 583520 205580 584960 205670
rect -960 201772 480 202012
rect 14181 195530 14247 195533
rect 14181 195528 15210 195530
rect 14181 195472 14186 195528
rect 14242 195472 15210 195528
rect 14181 195470 15210 195472
rect 14181 195467 14247 195470
rect 15150 194956 15210 195470
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188716 480 188956
rect 14089 182066 14155 182069
rect 14089 182064 15210 182066
rect 14089 182008 14094 182064
rect 14150 182008 15210 182064
rect 14089 182006 15210 182008
rect 14089 182003 14155 182006
rect 15150 181628 15210 182006
rect 580349 179210 580415 179213
rect 583520 179210 584960 179300
rect 580349 179208 584960 179210
rect 580349 179152 580354 179208
rect 580410 179152 584960 179208
rect 580349 179150 584960 179152
rect 580349 179147 580415 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 13997 168194 14063 168197
rect 15150 168194 15210 168300
rect 13997 168192 15210 168194
rect 13997 168136 14002 168192
rect 14058 168136 15210 168192
rect 13997 168134 15210 168136
rect 13997 168131 14063 168134
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3509 162890 3575 162893
rect -960 162888 3575 162890
rect -960 162832 3514 162888
rect 3570 162832 3575 162888
rect -960 162830 3575 162832
rect -960 162740 480 162830
rect 3509 162827 3575 162830
rect 13905 155546 13971 155549
rect 13905 155544 15210 155546
rect 13905 155488 13910 155544
rect 13966 155488 15210 155544
rect 13905 155486 15210 155488
rect 13905 155483 13971 155486
rect 15150 154972 15210 155486
rect 579797 152690 579863 152693
rect 583520 152690 584960 152780
rect 579797 152688 584960 152690
rect 579797 152632 579802 152688
rect 579858 152632 584960 152688
rect 579797 152630 584960 152632
rect 579797 152627 579863 152630
rect 583520 152540 584960 152630
rect -960 149684 480 149924
rect 13813 141946 13879 141949
rect 13813 141944 15210 141946
rect 13813 141888 13818 141944
rect 13874 141888 15210 141944
rect 13813 141886 15210 141888
rect 13813 141883 13879 141886
rect 15150 141644 15210 141886
rect 580257 139362 580323 139365
rect 583520 139362 584960 139452
rect 580257 139360 584960 139362
rect 580257 139304 580262 139360
rect 580318 139304 584960 139360
rect 580257 139302 584960 139304
rect 580257 139299 580323 139302
rect 583520 139212 584960 139302
rect -960 136628 480 136868
rect 12433 128210 12499 128213
rect 15150 128210 15210 128316
rect 12433 128208 15210 128210
rect 12433 128152 12438 128208
rect 12494 128152 15210 128208
rect 12433 128150 15210 128152
rect 12433 128147 12499 128150
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 12433 115562 12499 115565
rect 12433 115560 15210 115562
rect 12433 115504 12438 115560
rect 12494 115504 15210 115560
rect 12433 115502 15210 115504
rect 12433 115499 12499 115502
rect 15150 114988 15210 115502
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3601 110666 3667 110669
rect -960 110664 3667 110666
rect -960 110608 3606 110664
rect 3662 110608 3667 110664
rect -960 110606 3667 110608
rect -960 110516 480 110606
rect 3601 110603 3667 110606
rect 11697 102098 11763 102101
rect 11697 102096 15210 102098
rect 11697 102040 11702 102096
rect 11758 102040 15210 102096
rect 11697 102038 15210 102040
rect 11697 102035 11763 102038
rect 15150 101660 15210 102038
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97460 480 97700
rect 12433 88906 12499 88909
rect 12433 88904 15210 88906
rect 12433 88848 12438 88904
rect 12494 88848 15210 88904
rect 12433 88846 15210 88848
rect 12433 88843 12499 88846
rect 15150 88332 15210 88846
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84540 480 84780
rect 12433 75442 12499 75445
rect 12433 75440 15210 75442
rect 12433 75384 12438 75440
rect 12494 75384 15210 75440
rect 12433 75382 15210 75384
rect 12433 75379 12499 75382
rect 15150 75004 15210 75382
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3693 71634 3759 71637
rect -960 71632 3759 71634
rect -960 71576 3698 71632
rect 3754 71576 3759 71632
rect -960 71574 3759 71576
rect -960 71484 480 71574
rect 3693 71571 3759 71574
rect 12801 61978 12867 61981
rect 12801 61976 15210 61978
rect 12801 61920 12806 61976
rect 12862 61920 15210 61976
rect 12801 61918 15210 61920
rect 12801 61915 12867 61918
rect 15150 61676 15210 61918
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58428 480 58668
rect 11881 48922 11947 48925
rect 11881 48920 15210 48922
rect 11881 48864 11886 48920
rect 11942 48864 15210 48920
rect 11881 48862 15210 48864
rect 11881 48859 11947 48862
rect 15150 48348 15210 48862
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45372 480 45612
rect 13077 35458 13143 35461
rect 13077 35456 15210 35458
rect 13077 35400 13082 35456
rect 13138 35400 15210 35456
rect 13077 35398 15210 35400
rect 13077 35395 13143 35398
rect 15150 35020 15210 35398
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32316 480 32556
rect 13721 21178 13787 21181
rect 15150 21178 15210 21692
rect 13721 21176 15210 21178
rect 13721 21120 13726 21176
rect 13782 21120 15210 21176
rect 13721 21118 15210 21120
rect 13721 21115 13787 21118
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect -960 19260 480 19500
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6340 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 583520 6476 584960 6566
<< via3 >>
rect 13676 700436 13740 700500
rect 12756 700300 12820 700364
rect 469628 657052 469692 657116
rect 469628 653380 469692 653444
rect 12756 222124 12820 222188
rect 13676 208116 13740 208180
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 12755 700364 12821 700365
rect 12755 700300 12756 700364
rect 12820 700300 12821 700364
rect 12755 700299 12821 700300
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 12758 222189 12818 700299
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 13675 700500 13741 700501
rect 13675 700436 13676 700500
rect 13740 700436 13741 700500
rect 13675 700435 13741 700436
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 657000 13574 662058
rect 12755 222188 12821 222189
rect 12755 222124 12756 222188
rect 12820 222124 12821 222188
rect 12755 222123 12821 222124
rect 13678 208181 13738 700435
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 657000 20414 668898
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 657000 24134 672618
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 657000 27854 676338
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 657000 31574 680058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 657000 38414 686898
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 657000 42134 690618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 657000 45854 658338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 657000 49574 662058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 657000 56414 668898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 657000 60134 672618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 657000 63854 676338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 657000 67574 680058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 657000 74414 686898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 657000 78134 690618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 657000 81854 658338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 657000 85574 662058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 657000 92414 668898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 657000 96134 672618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 657000 99854 676338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 657000 103574 680058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 657000 110414 686898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 657000 114134 690618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 657000 117854 658338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 657000 121574 662058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 657000 128414 668898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 657000 132134 672618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 657000 135854 676338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 657000 139574 680058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 657000 146414 686898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 657000 150134 690618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 657000 153854 658338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 657000 157574 662058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 657000 164414 668898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 657000 168134 672618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 657000 171854 676338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 657000 175574 680058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 657000 182414 686898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 657000 186134 690618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 657000 189854 658338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 657000 193574 662058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 657000 200414 668898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 657000 204134 672618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 657000 207854 676338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 657000 211574 680058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 657000 218414 686898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 657000 222134 690618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 657000 225854 658338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 657000 229574 662058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 657000 236414 668898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 657000 240134 672618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 657000 243854 676338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 657000 247574 680058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 657000 254414 686898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 657000 258134 690618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 657000 261854 658338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 657000 265574 662058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 657000 272414 668898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 657000 276134 672618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 657000 279854 676338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 657000 283574 680058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 657000 290414 686898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 657000 294134 690618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 657000 297854 658338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 657000 301574 662058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 657000 308414 668898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 657000 312134 672618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 657000 315854 676338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 657000 319574 680058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 657000 326414 686898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 657000 330134 690618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 657000 333854 658338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 657000 337574 662058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 657000 344414 668898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 657000 348134 672618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 657000 351854 676338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 657000 355574 680058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 657000 362414 686898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 657000 366134 690618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 657000 369854 658338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 657000 373574 662058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 657000 380414 668898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 657000 384134 672618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 657000 387854 676338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 657000 391574 680058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 657000 398414 686898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 657000 402134 690618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 657000 405854 658338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 657000 409574 662058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 657000 416414 668898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 657000 420134 672618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 657000 423854 676338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 657000 427574 680058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 657000 434414 686898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 657000 438134 690618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 657000 441854 658338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 657000 445574 662058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 657000 452414 668898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 657000 456134 672618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 657000 459854 676338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 657000 463574 680058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469627 657116 469693 657117
rect 469627 657052 469628 657116
rect 469692 657052 469693 657116
rect 469627 657051 469693 657052
rect 469630 653445 469690 657051
rect 469794 657000 470414 686898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 657000 474134 690618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 657000 477854 658338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 657000 481574 662058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 657000 488414 668898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 657000 492134 672618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 657000 495854 676338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 657000 499574 680058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 657000 506414 686898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 657000 510134 690618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 657000 513854 658338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 657000 517574 662058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 657000 524414 668898
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 657000 528134 672618
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 657000 531854 676338
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 657000 535574 680058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 469627 653444 469693 653445
rect 469627 653380 469628 653444
rect 469692 653380 469693 653444
rect 469627 653379 469693 653380
rect 19208 651454 19528 651486
rect 19208 651218 19250 651454
rect 19486 651218 19528 651454
rect 19208 651134 19528 651218
rect 19208 650898 19250 651134
rect 19486 650898 19528 651134
rect 19208 650866 19528 650898
rect 49928 651454 50248 651486
rect 49928 651218 49970 651454
rect 50206 651218 50248 651454
rect 49928 651134 50248 651218
rect 49928 650898 49970 651134
rect 50206 650898 50248 651134
rect 49928 650866 50248 650898
rect 80648 651454 80968 651486
rect 80648 651218 80690 651454
rect 80926 651218 80968 651454
rect 80648 651134 80968 651218
rect 80648 650898 80690 651134
rect 80926 650898 80968 651134
rect 80648 650866 80968 650898
rect 111368 651454 111688 651486
rect 111368 651218 111410 651454
rect 111646 651218 111688 651454
rect 111368 651134 111688 651218
rect 111368 650898 111410 651134
rect 111646 650898 111688 651134
rect 111368 650866 111688 650898
rect 142088 651454 142408 651486
rect 142088 651218 142130 651454
rect 142366 651218 142408 651454
rect 142088 651134 142408 651218
rect 142088 650898 142130 651134
rect 142366 650898 142408 651134
rect 142088 650866 142408 650898
rect 172808 651454 173128 651486
rect 172808 651218 172850 651454
rect 173086 651218 173128 651454
rect 172808 651134 173128 651218
rect 172808 650898 172850 651134
rect 173086 650898 173128 651134
rect 172808 650866 173128 650898
rect 203528 651454 203848 651486
rect 203528 651218 203570 651454
rect 203806 651218 203848 651454
rect 203528 651134 203848 651218
rect 203528 650898 203570 651134
rect 203806 650898 203848 651134
rect 203528 650866 203848 650898
rect 234248 651454 234568 651486
rect 234248 651218 234290 651454
rect 234526 651218 234568 651454
rect 234248 651134 234568 651218
rect 234248 650898 234290 651134
rect 234526 650898 234568 651134
rect 234248 650866 234568 650898
rect 264968 651454 265288 651486
rect 264968 651218 265010 651454
rect 265246 651218 265288 651454
rect 264968 651134 265288 651218
rect 264968 650898 265010 651134
rect 265246 650898 265288 651134
rect 264968 650866 265288 650898
rect 295688 651454 296008 651486
rect 295688 651218 295730 651454
rect 295966 651218 296008 651454
rect 295688 651134 296008 651218
rect 295688 650898 295730 651134
rect 295966 650898 296008 651134
rect 295688 650866 296008 650898
rect 326408 651454 326728 651486
rect 326408 651218 326450 651454
rect 326686 651218 326728 651454
rect 326408 651134 326728 651218
rect 326408 650898 326450 651134
rect 326686 650898 326728 651134
rect 326408 650866 326728 650898
rect 357128 651454 357448 651486
rect 357128 651218 357170 651454
rect 357406 651218 357448 651454
rect 357128 651134 357448 651218
rect 357128 650898 357170 651134
rect 357406 650898 357448 651134
rect 357128 650866 357448 650898
rect 387848 651454 388168 651486
rect 387848 651218 387890 651454
rect 388126 651218 388168 651454
rect 387848 651134 388168 651218
rect 387848 650898 387890 651134
rect 388126 650898 388168 651134
rect 387848 650866 388168 650898
rect 418568 651454 418888 651486
rect 418568 651218 418610 651454
rect 418846 651218 418888 651454
rect 418568 651134 418888 651218
rect 418568 650898 418610 651134
rect 418846 650898 418888 651134
rect 418568 650866 418888 650898
rect 449288 651454 449608 651486
rect 449288 651218 449330 651454
rect 449566 651218 449608 651454
rect 449288 651134 449608 651218
rect 449288 650898 449330 651134
rect 449566 650898 449608 651134
rect 449288 650866 449608 650898
rect 480008 651454 480328 651486
rect 480008 651218 480050 651454
rect 480286 651218 480328 651454
rect 480008 651134 480328 651218
rect 480008 650898 480050 651134
rect 480286 650898 480328 651134
rect 480008 650866 480328 650898
rect 510728 651454 511048 651486
rect 510728 651218 510770 651454
rect 511006 651218 511048 651454
rect 510728 651134 511048 651218
rect 510728 650898 510770 651134
rect 511006 650898 511048 651134
rect 510728 650866 511048 650898
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 34568 633454 34888 633486
rect 34568 633218 34610 633454
rect 34846 633218 34888 633454
rect 34568 633134 34888 633218
rect 34568 632898 34610 633134
rect 34846 632898 34888 633134
rect 34568 632866 34888 632898
rect 65288 633454 65608 633486
rect 65288 633218 65330 633454
rect 65566 633218 65608 633454
rect 65288 633134 65608 633218
rect 65288 632898 65330 633134
rect 65566 632898 65608 633134
rect 65288 632866 65608 632898
rect 96008 633454 96328 633486
rect 96008 633218 96050 633454
rect 96286 633218 96328 633454
rect 96008 633134 96328 633218
rect 96008 632898 96050 633134
rect 96286 632898 96328 633134
rect 96008 632866 96328 632898
rect 126728 633454 127048 633486
rect 126728 633218 126770 633454
rect 127006 633218 127048 633454
rect 126728 633134 127048 633218
rect 126728 632898 126770 633134
rect 127006 632898 127048 633134
rect 126728 632866 127048 632898
rect 157448 633454 157768 633486
rect 157448 633218 157490 633454
rect 157726 633218 157768 633454
rect 157448 633134 157768 633218
rect 157448 632898 157490 633134
rect 157726 632898 157768 633134
rect 157448 632866 157768 632898
rect 188168 633454 188488 633486
rect 188168 633218 188210 633454
rect 188446 633218 188488 633454
rect 188168 633134 188488 633218
rect 188168 632898 188210 633134
rect 188446 632898 188488 633134
rect 188168 632866 188488 632898
rect 218888 633454 219208 633486
rect 218888 633218 218930 633454
rect 219166 633218 219208 633454
rect 218888 633134 219208 633218
rect 218888 632898 218930 633134
rect 219166 632898 219208 633134
rect 218888 632866 219208 632898
rect 249608 633454 249928 633486
rect 249608 633218 249650 633454
rect 249886 633218 249928 633454
rect 249608 633134 249928 633218
rect 249608 632898 249650 633134
rect 249886 632898 249928 633134
rect 249608 632866 249928 632898
rect 280328 633454 280648 633486
rect 280328 633218 280370 633454
rect 280606 633218 280648 633454
rect 280328 633134 280648 633218
rect 280328 632898 280370 633134
rect 280606 632898 280648 633134
rect 280328 632866 280648 632898
rect 311048 633454 311368 633486
rect 311048 633218 311090 633454
rect 311326 633218 311368 633454
rect 311048 633134 311368 633218
rect 311048 632898 311090 633134
rect 311326 632898 311368 633134
rect 311048 632866 311368 632898
rect 341768 633454 342088 633486
rect 341768 633218 341810 633454
rect 342046 633218 342088 633454
rect 341768 633134 342088 633218
rect 341768 632898 341810 633134
rect 342046 632898 342088 633134
rect 341768 632866 342088 632898
rect 372488 633454 372808 633486
rect 372488 633218 372530 633454
rect 372766 633218 372808 633454
rect 372488 633134 372808 633218
rect 372488 632898 372530 633134
rect 372766 632898 372808 633134
rect 372488 632866 372808 632898
rect 403208 633454 403528 633486
rect 403208 633218 403250 633454
rect 403486 633218 403528 633454
rect 403208 633134 403528 633218
rect 403208 632898 403250 633134
rect 403486 632898 403528 633134
rect 403208 632866 403528 632898
rect 433928 633454 434248 633486
rect 433928 633218 433970 633454
rect 434206 633218 434248 633454
rect 433928 633134 434248 633218
rect 433928 632898 433970 633134
rect 434206 632898 434248 633134
rect 433928 632866 434248 632898
rect 464648 633454 464968 633486
rect 464648 633218 464690 633454
rect 464926 633218 464968 633454
rect 464648 633134 464968 633218
rect 464648 632898 464690 633134
rect 464926 632898 464968 633134
rect 464648 632866 464968 632898
rect 495368 633454 495688 633486
rect 495368 633218 495410 633454
rect 495646 633218 495688 633454
rect 495368 633134 495688 633218
rect 495368 632898 495410 633134
rect 495646 632898 495688 633134
rect 495368 632866 495688 632898
rect 526088 633454 526408 633486
rect 526088 633218 526130 633454
rect 526366 633218 526408 633454
rect 526088 633134 526408 633218
rect 526088 632898 526130 633134
rect 526366 632898 526408 633134
rect 526088 632866 526408 632898
rect 19208 615454 19528 615486
rect 19208 615218 19250 615454
rect 19486 615218 19528 615454
rect 19208 615134 19528 615218
rect 19208 614898 19250 615134
rect 19486 614898 19528 615134
rect 19208 614866 19528 614898
rect 49928 615454 50248 615486
rect 49928 615218 49970 615454
rect 50206 615218 50248 615454
rect 49928 615134 50248 615218
rect 49928 614898 49970 615134
rect 50206 614898 50248 615134
rect 49928 614866 50248 614898
rect 80648 615454 80968 615486
rect 80648 615218 80690 615454
rect 80926 615218 80968 615454
rect 80648 615134 80968 615218
rect 80648 614898 80690 615134
rect 80926 614898 80968 615134
rect 80648 614866 80968 614898
rect 111368 615454 111688 615486
rect 111368 615218 111410 615454
rect 111646 615218 111688 615454
rect 111368 615134 111688 615218
rect 111368 614898 111410 615134
rect 111646 614898 111688 615134
rect 111368 614866 111688 614898
rect 142088 615454 142408 615486
rect 142088 615218 142130 615454
rect 142366 615218 142408 615454
rect 142088 615134 142408 615218
rect 142088 614898 142130 615134
rect 142366 614898 142408 615134
rect 142088 614866 142408 614898
rect 172808 615454 173128 615486
rect 172808 615218 172850 615454
rect 173086 615218 173128 615454
rect 172808 615134 173128 615218
rect 172808 614898 172850 615134
rect 173086 614898 173128 615134
rect 172808 614866 173128 614898
rect 203528 615454 203848 615486
rect 203528 615218 203570 615454
rect 203806 615218 203848 615454
rect 203528 615134 203848 615218
rect 203528 614898 203570 615134
rect 203806 614898 203848 615134
rect 203528 614866 203848 614898
rect 234248 615454 234568 615486
rect 234248 615218 234290 615454
rect 234526 615218 234568 615454
rect 234248 615134 234568 615218
rect 234248 614898 234290 615134
rect 234526 614898 234568 615134
rect 234248 614866 234568 614898
rect 264968 615454 265288 615486
rect 264968 615218 265010 615454
rect 265246 615218 265288 615454
rect 264968 615134 265288 615218
rect 264968 614898 265010 615134
rect 265246 614898 265288 615134
rect 264968 614866 265288 614898
rect 295688 615454 296008 615486
rect 295688 615218 295730 615454
rect 295966 615218 296008 615454
rect 295688 615134 296008 615218
rect 295688 614898 295730 615134
rect 295966 614898 296008 615134
rect 295688 614866 296008 614898
rect 326408 615454 326728 615486
rect 326408 615218 326450 615454
rect 326686 615218 326728 615454
rect 326408 615134 326728 615218
rect 326408 614898 326450 615134
rect 326686 614898 326728 615134
rect 326408 614866 326728 614898
rect 357128 615454 357448 615486
rect 357128 615218 357170 615454
rect 357406 615218 357448 615454
rect 357128 615134 357448 615218
rect 357128 614898 357170 615134
rect 357406 614898 357448 615134
rect 357128 614866 357448 614898
rect 387848 615454 388168 615486
rect 387848 615218 387890 615454
rect 388126 615218 388168 615454
rect 387848 615134 388168 615218
rect 387848 614898 387890 615134
rect 388126 614898 388168 615134
rect 387848 614866 388168 614898
rect 418568 615454 418888 615486
rect 418568 615218 418610 615454
rect 418846 615218 418888 615454
rect 418568 615134 418888 615218
rect 418568 614898 418610 615134
rect 418846 614898 418888 615134
rect 418568 614866 418888 614898
rect 449288 615454 449608 615486
rect 449288 615218 449330 615454
rect 449566 615218 449608 615454
rect 449288 615134 449608 615218
rect 449288 614898 449330 615134
rect 449566 614898 449608 615134
rect 449288 614866 449608 614898
rect 480008 615454 480328 615486
rect 480008 615218 480050 615454
rect 480286 615218 480328 615454
rect 480008 615134 480328 615218
rect 480008 614898 480050 615134
rect 480286 614898 480328 615134
rect 480008 614866 480328 614898
rect 510728 615454 511048 615486
rect 510728 615218 510770 615454
rect 511006 615218 511048 615454
rect 510728 615134 511048 615218
rect 510728 614898 510770 615134
rect 511006 614898 511048 615134
rect 510728 614866 511048 614898
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 34568 597454 34888 597486
rect 34568 597218 34610 597454
rect 34846 597218 34888 597454
rect 34568 597134 34888 597218
rect 34568 596898 34610 597134
rect 34846 596898 34888 597134
rect 34568 596866 34888 596898
rect 65288 597454 65608 597486
rect 65288 597218 65330 597454
rect 65566 597218 65608 597454
rect 65288 597134 65608 597218
rect 65288 596898 65330 597134
rect 65566 596898 65608 597134
rect 65288 596866 65608 596898
rect 96008 597454 96328 597486
rect 96008 597218 96050 597454
rect 96286 597218 96328 597454
rect 96008 597134 96328 597218
rect 96008 596898 96050 597134
rect 96286 596898 96328 597134
rect 96008 596866 96328 596898
rect 126728 597454 127048 597486
rect 126728 597218 126770 597454
rect 127006 597218 127048 597454
rect 126728 597134 127048 597218
rect 126728 596898 126770 597134
rect 127006 596898 127048 597134
rect 126728 596866 127048 596898
rect 157448 597454 157768 597486
rect 157448 597218 157490 597454
rect 157726 597218 157768 597454
rect 157448 597134 157768 597218
rect 157448 596898 157490 597134
rect 157726 596898 157768 597134
rect 157448 596866 157768 596898
rect 188168 597454 188488 597486
rect 188168 597218 188210 597454
rect 188446 597218 188488 597454
rect 188168 597134 188488 597218
rect 188168 596898 188210 597134
rect 188446 596898 188488 597134
rect 188168 596866 188488 596898
rect 218888 597454 219208 597486
rect 218888 597218 218930 597454
rect 219166 597218 219208 597454
rect 218888 597134 219208 597218
rect 218888 596898 218930 597134
rect 219166 596898 219208 597134
rect 218888 596866 219208 596898
rect 249608 597454 249928 597486
rect 249608 597218 249650 597454
rect 249886 597218 249928 597454
rect 249608 597134 249928 597218
rect 249608 596898 249650 597134
rect 249886 596898 249928 597134
rect 249608 596866 249928 596898
rect 280328 597454 280648 597486
rect 280328 597218 280370 597454
rect 280606 597218 280648 597454
rect 280328 597134 280648 597218
rect 280328 596898 280370 597134
rect 280606 596898 280648 597134
rect 280328 596866 280648 596898
rect 311048 597454 311368 597486
rect 311048 597218 311090 597454
rect 311326 597218 311368 597454
rect 311048 597134 311368 597218
rect 311048 596898 311090 597134
rect 311326 596898 311368 597134
rect 311048 596866 311368 596898
rect 341768 597454 342088 597486
rect 341768 597218 341810 597454
rect 342046 597218 342088 597454
rect 341768 597134 342088 597218
rect 341768 596898 341810 597134
rect 342046 596898 342088 597134
rect 341768 596866 342088 596898
rect 372488 597454 372808 597486
rect 372488 597218 372530 597454
rect 372766 597218 372808 597454
rect 372488 597134 372808 597218
rect 372488 596898 372530 597134
rect 372766 596898 372808 597134
rect 372488 596866 372808 596898
rect 403208 597454 403528 597486
rect 403208 597218 403250 597454
rect 403486 597218 403528 597454
rect 403208 597134 403528 597218
rect 403208 596898 403250 597134
rect 403486 596898 403528 597134
rect 403208 596866 403528 596898
rect 433928 597454 434248 597486
rect 433928 597218 433970 597454
rect 434206 597218 434248 597454
rect 433928 597134 434248 597218
rect 433928 596898 433970 597134
rect 434206 596898 434248 597134
rect 433928 596866 434248 596898
rect 464648 597454 464968 597486
rect 464648 597218 464690 597454
rect 464926 597218 464968 597454
rect 464648 597134 464968 597218
rect 464648 596898 464690 597134
rect 464926 596898 464968 597134
rect 464648 596866 464968 596898
rect 495368 597454 495688 597486
rect 495368 597218 495410 597454
rect 495646 597218 495688 597454
rect 495368 597134 495688 597218
rect 495368 596898 495410 597134
rect 495646 596898 495688 597134
rect 495368 596866 495688 596898
rect 526088 597454 526408 597486
rect 526088 597218 526130 597454
rect 526366 597218 526408 597454
rect 526088 597134 526408 597218
rect 526088 596898 526130 597134
rect 526366 596898 526408 597134
rect 526088 596866 526408 596898
rect 19208 579454 19528 579486
rect 19208 579218 19250 579454
rect 19486 579218 19528 579454
rect 19208 579134 19528 579218
rect 19208 578898 19250 579134
rect 19486 578898 19528 579134
rect 19208 578866 19528 578898
rect 49928 579454 50248 579486
rect 49928 579218 49970 579454
rect 50206 579218 50248 579454
rect 49928 579134 50248 579218
rect 49928 578898 49970 579134
rect 50206 578898 50248 579134
rect 49928 578866 50248 578898
rect 80648 579454 80968 579486
rect 80648 579218 80690 579454
rect 80926 579218 80968 579454
rect 80648 579134 80968 579218
rect 80648 578898 80690 579134
rect 80926 578898 80968 579134
rect 80648 578866 80968 578898
rect 111368 579454 111688 579486
rect 111368 579218 111410 579454
rect 111646 579218 111688 579454
rect 111368 579134 111688 579218
rect 111368 578898 111410 579134
rect 111646 578898 111688 579134
rect 111368 578866 111688 578898
rect 142088 579454 142408 579486
rect 142088 579218 142130 579454
rect 142366 579218 142408 579454
rect 142088 579134 142408 579218
rect 142088 578898 142130 579134
rect 142366 578898 142408 579134
rect 142088 578866 142408 578898
rect 172808 579454 173128 579486
rect 172808 579218 172850 579454
rect 173086 579218 173128 579454
rect 172808 579134 173128 579218
rect 172808 578898 172850 579134
rect 173086 578898 173128 579134
rect 172808 578866 173128 578898
rect 203528 579454 203848 579486
rect 203528 579218 203570 579454
rect 203806 579218 203848 579454
rect 203528 579134 203848 579218
rect 203528 578898 203570 579134
rect 203806 578898 203848 579134
rect 203528 578866 203848 578898
rect 234248 579454 234568 579486
rect 234248 579218 234290 579454
rect 234526 579218 234568 579454
rect 234248 579134 234568 579218
rect 234248 578898 234290 579134
rect 234526 578898 234568 579134
rect 234248 578866 234568 578898
rect 264968 579454 265288 579486
rect 264968 579218 265010 579454
rect 265246 579218 265288 579454
rect 264968 579134 265288 579218
rect 264968 578898 265010 579134
rect 265246 578898 265288 579134
rect 264968 578866 265288 578898
rect 295688 579454 296008 579486
rect 295688 579218 295730 579454
rect 295966 579218 296008 579454
rect 295688 579134 296008 579218
rect 295688 578898 295730 579134
rect 295966 578898 296008 579134
rect 295688 578866 296008 578898
rect 326408 579454 326728 579486
rect 326408 579218 326450 579454
rect 326686 579218 326728 579454
rect 326408 579134 326728 579218
rect 326408 578898 326450 579134
rect 326686 578898 326728 579134
rect 326408 578866 326728 578898
rect 357128 579454 357448 579486
rect 357128 579218 357170 579454
rect 357406 579218 357448 579454
rect 357128 579134 357448 579218
rect 357128 578898 357170 579134
rect 357406 578898 357448 579134
rect 357128 578866 357448 578898
rect 387848 579454 388168 579486
rect 387848 579218 387890 579454
rect 388126 579218 388168 579454
rect 387848 579134 388168 579218
rect 387848 578898 387890 579134
rect 388126 578898 388168 579134
rect 387848 578866 388168 578898
rect 418568 579454 418888 579486
rect 418568 579218 418610 579454
rect 418846 579218 418888 579454
rect 418568 579134 418888 579218
rect 418568 578898 418610 579134
rect 418846 578898 418888 579134
rect 418568 578866 418888 578898
rect 449288 579454 449608 579486
rect 449288 579218 449330 579454
rect 449566 579218 449608 579454
rect 449288 579134 449608 579218
rect 449288 578898 449330 579134
rect 449566 578898 449608 579134
rect 449288 578866 449608 578898
rect 480008 579454 480328 579486
rect 480008 579218 480050 579454
rect 480286 579218 480328 579454
rect 480008 579134 480328 579218
rect 480008 578898 480050 579134
rect 480286 578898 480328 579134
rect 480008 578866 480328 578898
rect 510728 579454 511048 579486
rect 510728 579218 510770 579454
rect 511006 579218 511048 579454
rect 510728 579134 511048 579218
rect 510728 578898 510770 579134
rect 511006 578898 511048 579134
rect 510728 578866 511048 578898
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 34568 561454 34888 561486
rect 34568 561218 34610 561454
rect 34846 561218 34888 561454
rect 34568 561134 34888 561218
rect 34568 560898 34610 561134
rect 34846 560898 34888 561134
rect 34568 560866 34888 560898
rect 65288 561454 65608 561486
rect 65288 561218 65330 561454
rect 65566 561218 65608 561454
rect 65288 561134 65608 561218
rect 65288 560898 65330 561134
rect 65566 560898 65608 561134
rect 65288 560866 65608 560898
rect 96008 561454 96328 561486
rect 96008 561218 96050 561454
rect 96286 561218 96328 561454
rect 96008 561134 96328 561218
rect 96008 560898 96050 561134
rect 96286 560898 96328 561134
rect 96008 560866 96328 560898
rect 126728 561454 127048 561486
rect 126728 561218 126770 561454
rect 127006 561218 127048 561454
rect 126728 561134 127048 561218
rect 126728 560898 126770 561134
rect 127006 560898 127048 561134
rect 126728 560866 127048 560898
rect 157448 561454 157768 561486
rect 157448 561218 157490 561454
rect 157726 561218 157768 561454
rect 157448 561134 157768 561218
rect 157448 560898 157490 561134
rect 157726 560898 157768 561134
rect 157448 560866 157768 560898
rect 188168 561454 188488 561486
rect 188168 561218 188210 561454
rect 188446 561218 188488 561454
rect 188168 561134 188488 561218
rect 188168 560898 188210 561134
rect 188446 560898 188488 561134
rect 188168 560866 188488 560898
rect 218888 561454 219208 561486
rect 218888 561218 218930 561454
rect 219166 561218 219208 561454
rect 218888 561134 219208 561218
rect 218888 560898 218930 561134
rect 219166 560898 219208 561134
rect 218888 560866 219208 560898
rect 249608 561454 249928 561486
rect 249608 561218 249650 561454
rect 249886 561218 249928 561454
rect 249608 561134 249928 561218
rect 249608 560898 249650 561134
rect 249886 560898 249928 561134
rect 249608 560866 249928 560898
rect 280328 561454 280648 561486
rect 280328 561218 280370 561454
rect 280606 561218 280648 561454
rect 280328 561134 280648 561218
rect 280328 560898 280370 561134
rect 280606 560898 280648 561134
rect 280328 560866 280648 560898
rect 311048 561454 311368 561486
rect 311048 561218 311090 561454
rect 311326 561218 311368 561454
rect 311048 561134 311368 561218
rect 311048 560898 311090 561134
rect 311326 560898 311368 561134
rect 311048 560866 311368 560898
rect 341768 561454 342088 561486
rect 341768 561218 341810 561454
rect 342046 561218 342088 561454
rect 341768 561134 342088 561218
rect 341768 560898 341810 561134
rect 342046 560898 342088 561134
rect 341768 560866 342088 560898
rect 372488 561454 372808 561486
rect 372488 561218 372530 561454
rect 372766 561218 372808 561454
rect 372488 561134 372808 561218
rect 372488 560898 372530 561134
rect 372766 560898 372808 561134
rect 372488 560866 372808 560898
rect 403208 561454 403528 561486
rect 403208 561218 403250 561454
rect 403486 561218 403528 561454
rect 403208 561134 403528 561218
rect 403208 560898 403250 561134
rect 403486 560898 403528 561134
rect 403208 560866 403528 560898
rect 433928 561454 434248 561486
rect 433928 561218 433970 561454
rect 434206 561218 434248 561454
rect 433928 561134 434248 561218
rect 433928 560898 433970 561134
rect 434206 560898 434248 561134
rect 433928 560866 434248 560898
rect 464648 561454 464968 561486
rect 464648 561218 464690 561454
rect 464926 561218 464968 561454
rect 464648 561134 464968 561218
rect 464648 560898 464690 561134
rect 464926 560898 464968 561134
rect 464648 560866 464968 560898
rect 495368 561454 495688 561486
rect 495368 561218 495410 561454
rect 495646 561218 495688 561454
rect 495368 561134 495688 561218
rect 495368 560898 495410 561134
rect 495646 560898 495688 561134
rect 495368 560866 495688 560898
rect 526088 561454 526408 561486
rect 526088 561218 526130 561454
rect 526366 561218 526408 561454
rect 526088 561134 526408 561218
rect 526088 560898 526130 561134
rect 526366 560898 526408 561134
rect 526088 560866 526408 560898
rect 19208 543454 19528 543486
rect 19208 543218 19250 543454
rect 19486 543218 19528 543454
rect 19208 543134 19528 543218
rect 19208 542898 19250 543134
rect 19486 542898 19528 543134
rect 19208 542866 19528 542898
rect 49928 543454 50248 543486
rect 49928 543218 49970 543454
rect 50206 543218 50248 543454
rect 49928 543134 50248 543218
rect 49928 542898 49970 543134
rect 50206 542898 50248 543134
rect 49928 542866 50248 542898
rect 80648 543454 80968 543486
rect 80648 543218 80690 543454
rect 80926 543218 80968 543454
rect 80648 543134 80968 543218
rect 80648 542898 80690 543134
rect 80926 542898 80968 543134
rect 80648 542866 80968 542898
rect 111368 543454 111688 543486
rect 111368 543218 111410 543454
rect 111646 543218 111688 543454
rect 111368 543134 111688 543218
rect 111368 542898 111410 543134
rect 111646 542898 111688 543134
rect 111368 542866 111688 542898
rect 142088 543454 142408 543486
rect 142088 543218 142130 543454
rect 142366 543218 142408 543454
rect 142088 543134 142408 543218
rect 142088 542898 142130 543134
rect 142366 542898 142408 543134
rect 142088 542866 142408 542898
rect 172808 543454 173128 543486
rect 172808 543218 172850 543454
rect 173086 543218 173128 543454
rect 172808 543134 173128 543218
rect 172808 542898 172850 543134
rect 173086 542898 173128 543134
rect 172808 542866 173128 542898
rect 203528 543454 203848 543486
rect 203528 543218 203570 543454
rect 203806 543218 203848 543454
rect 203528 543134 203848 543218
rect 203528 542898 203570 543134
rect 203806 542898 203848 543134
rect 203528 542866 203848 542898
rect 234248 543454 234568 543486
rect 234248 543218 234290 543454
rect 234526 543218 234568 543454
rect 234248 543134 234568 543218
rect 234248 542898 234290 543134
rect 234526 542898 234568 543134
rect 234248 542866 234568 542898
rect 264968 543454 265288 543486
rect 264968 543218 265010 543454
rect 265246 543218 265288 543454
rect 264968 543134 265288 543218
rect 264968 542898 265010 543134
rect 265246 542898 265288 543134
rect 264968 542866 265288 542898
rect 295688 543454 296008 543486
rect 295688 543218 295730 543454
rect 295966 543218 296008 543454
rect 295688 543134 296008 543218
rect 295688 542898 295730 543134
rect 295966 542898 296008 543134
rect 295688 542866 296008 542898
rect 326408 543454 326728 543486
rect 326408 543218 326450 543454
rect 326686 543218 326728 543454
rect 326408 543134 326728 543218
rect 326408 542898 326450 543134
rect 326686 542898 326728 543134
rect 326408 542866 326728 542898
rect 357128 543454 357448 543486
rect 357128 543218 357170 543454
rect 357406 543218 357448 543454
rect 357128 543134 357448 543218
rect 357128 542898 357170 543134
rect 357406 542898 357448 543134
rect 357128 542866 357448 542898
rect 387848 543454 388168 543486
rect 387848 543218 387890 543454
rect 388126 543218 388168 543454
rect 387848 543134 388168 543218
rect 387848 542898 387890 543134
rect 388126 542898 388168 543134
rect 387848 542866 388168 542898
rect 418568 543454 418888 543486
rect 418568 543218 418610 543454
rect 418846 543218 418888 543454
rect 418568 543134 418888 543218
rect 418568 542898 418610 543134
rect 418846 542898 418888 543134
rect 418568 542866 418888 542898
rect 449288 543454 449608 543486
rect 449288 543218 449330 543454
rect 449566 543218 449608 543454
rect 449288 543134 449608 543218
rect 449288 542898 449330 543134
rect 449566 542898 449608 543134
rect 449288 542866 449608 542898
rect 480008 543454 480328 543486
rect 480008 543218 480050 543454
rect 480286 543218 480328 543454
rect 480008 543134 480328 543218
rect 480008 542898 480050 543134
rect 480286 542898 480328 543134
rect 480008 542866 480328 542898
rect 510728 543454 511048 543486
rect 510728 543218 510770 543454
rect 511006 543218 511048 543454
rect 510728 543134 511048 543218
rect 510728 542898 510770 543134
rect 511006 542898 511048 543134
rect 510728 542866 511048 542898
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 34568 525454 34888 525486
rect 34568 525218 34610 525454
rect 34846 525218 34888 525454
rect 34568 525134 34888 525218
rect 34568 524898 34610 525134
rect 34846 524898 34888 525134
rect 34568 524866 34888 524898
rect 65288 525454 65608 525486
rect 65288 525218 65330 525454
rect 65566 525218 65608 525454
rect 65288 525134 65608 525218
rect 65288 524898 65330 525134
rect 65566 524898 65608 525134
rect 65288 524866 65608 524898
rect 96008 525454 96328 525486
rect 96008 525218 96050 525454
rect 96286 525218 96328 525454
rect 96008 525134 96328 525218
rect 96008 524898 96050 525134
rect 96286 524898 96328 525134
rect 96008 524866 96328 524898
rect 126728 525454 127048 525486
rect 126728 525218 126770 525454
rect 127006 525218 127048 525454
rect 126728 525134 127048 525218
rect 126728 524898 126770 525134
rect 127006 524898 127048 525134
rect 126728 524866 127048 524898
rect 157448 525454 157768 525486
rect 157448 525218 157490 525454
rect 157726 525218 157768 525454
rect 157448 525134 157768 525218
rect 157448 524898 157490 525134
rect 157726 524898 157768 525134
rect 157448 524866 157768 524898
rect 188168 525454 188488 525486
rect 188168 525218 188210 525454
rect 188446 525218 188488 525454
rect 188168 525134 188488 525218
rect 188168 524898 188210 525134
rect 188446 524898 188488 525134
rect 188168 524866 188488 524898
rect 218888 525454 219208 525486
rect 218888 525218 218930 525454
rect 219166 525218 219208 525454
rect 218888 525134 219208 525218
rect 218888 524898 218930 525134
rect 219166 524898 219208 525134
rect 218888 524866 219208 524898
rect 249608 525454 249928 525486
rect 249608 525218 249650 525454
rect 249886 525218 249928 525454
rect 249608 525134 249928 525218
rect 249608 524898 249650 525134
rect 249886 524898 249928 525134
rect 249608 524866 249928 524898
rect 280328 525454 280648 525486
rect 280328 525218 280370 525454
rect 280606 525218 280648 525454
rect 280328 525134 280648 525218
rect 280328 524898 280370 525134
rect 280606 524898 280648 525134
rect 280328 524866 280648 524898
rect 311048 525454 311368 525486
rect 311048 525218 311090 525454
rect 311326 525218 311368 525454
rect 311048 525134 311368 525218
rect 311048 524898 311090 525134
rect 311326 524898 311368 525134
rect 311048 524866 311368 524898
rect 341768 525454 342088 525486
rect 341768 525218 341810 525454
rect 342046 525218 342088 525454
rect 341768 525134 342088 525218
rect 341768 524898 341810 525134
rect 342046 524898 342088 525134
rect 341768 524866 342088 524898
rect 372488 525454 372808 525486
rect 372488 525218 372530 525454
rect 372766 525218 372808 525454
rect 372488 525134 372808 525218
rect 372488 524898 372530 525134
rect 372766 524898 372808 525134
rect 372488 524866 372808 524898
rect 403208 525454 403528 525486
rect 403208 525218 403250 525454
rect 403486 525218 403528 525454
rect 403208 525134 403528 525218
rect 403208 524898 403250 525134
rect 403486 524898 403528 525134
rect 403208 524866 403528 524898
rect 433928 525454 434248 525486
rect 433928 525218 433970 525454
rect 434206 525218 434248 525454
rect 433928 525134 434248 525218
rect 433928 524898 433970 525134
rect 434206 524898 434248 525134
rect 433928 524866 434248 524898
rect 464648 525454 464968 525486
rect 464648 525218 464690 525454
rect 464926 525218 464968 525454
rect 464648 525134 464968 525218
rect 464648 524898 464690 525134
rect 464926 524898 464968 525134
rect 464648 524866 464968 524898
rect 495368 525454 495688 525486
rect 495368 525218 495410 525454
rect 495646 525218 495688 525454
rect 495368 525134 495688 525218
rect 495368 524898 495410 525134
rect 495646 524898 495688 525134
rect 495368 524866 495688 524898
rect 526088 525454 526408 525486
rect 526088 525218 526130 525454
rect 526366 525218 526408 525454
rect 526088 525134 526408 525218
rect 526088 524898 526130 525134
rect 526366 524898 526408 525134
rect 526088 524866 526408 524898
rect 19208 507454 19528 507486
rect 19208 507218 19250 507454
rect 19486 507218 19528 507454
rect 19208 507134 19528 507218
rect 19208 506898 19250 507134
rect 19486 506898 19528 507134
rect 19208 506866 19528 506898
rect 49928 507454 50248 507486
rect 49928 507218 49970 507454
rect 50206 507218 50248 507454
rect 49928 507134 50248 507218
rect 49928 506898 49970 507134
rect 50206 506898 50248 507134
rect 49928 506866 50248 506898
rect 80648 507454 80968 507486
rect 80648 507218 80690 507454
rect 80926 507218 80968 507454
rect 80648 507134 80968 507218
rect 80648 506898 80690 507134
rect 80926 506898 80968 507134
rect 80648 506866 80968 506898
rect 111368 507454 111688 507486
rect 111368 507218 111410 507454
rect 111646 507218 111688 507454
rect 111368 507134 111688 507218
rect 111368 506898 111410 507134
rect 111646 506898 111688 507134
rect 111368 506866 111688 506898
rect 142088 507454 142408 507486
rect 142088 507218 142130 507454
rect 142366 507218 142408 507454
rect 142088 507134 142408 507218
rect 142088 506898 142130 507134
rect 142366 506898 142408 507134
rect 142088 506866 142408 506898
rect 172808 507454 173128 507486
rect 172808 507218 172850 507454
rect 173086 507218 173128 507454
rect 172808 507134 173128 507218
rect 172808 506898 172850 507134
rect 173086 506898 173128 507134
rect 172808 506866 173128 506898
rect 203528 507454 203848 507486
rect 203528 507218 203570 507454
rect 203806 507218 203848 507454
rect 203528 507134 203848 507218
rect 203528 506898 203570 507134
rect 203806 506898 203848 507134
rect 203528 506866 203848 506898
rect 234248 507454 234568 507486
rect 234248 507218 234290 507454
rect 234526 507218 234568 507454
rect 234248 507134 234568 507218
rect 234248 506898 234290 507134
rect 234526 506898 234568 507134
rect 234248 506866 234568 506898
rect 264968 507454 265288 507486
rect 264968 507218 265010 507454
rect 265246 507218 265288 507454
rect 264968 507134 265288 507218
rect 264968 506898 265010 507134
rect 265246 506898 265288 507134
rect 264968 506866 265288 506898
rect 295688 507454 296008 507486
rect 295688 507218 295730 507454
rect 295966 507218 296008 507454
rect 295688 507134 296008 507218
rect 295688 506898 295730 507134
rect 295966 506898 296008 507134
rect 295688 506866 296008 506898
rect 326408 507454 326728 507486
rect 326408 507218 326450 507454
rect 326686 507218 326728 507454
rect 326408 507134 326728 507218
rect 326408 506898 326450 507134
rect 326686 506898 326728 507134
rect 326408 506866 326728 506898
rect 357128 507454 357448 507486
rect 357128 507218 357170 507454
rect 357406 507218 357448 507454
rect 357128 507134 357448 507218
rect 357128 506898 357170 507134
rect 357406 506898 357448 507134
rect 357128 506866 357448 506898
rect 387848 507454 388168 507486
rect 387848 507218 387890 507454
rect 388126 507218 388168 507454
rect 387848 507134 388168 507218
rect 387848 506898 387890 507134
rect 388126 506898 388168 507134
rect 387848 506866 388168 506898
rect 418568 507454 418888 507486
rect 418568 507218 418610 507454
rect 418846 507218 418888 507454
rect 418568 507134 418888 507218
rect 418568 506898 418610 507134
rect 418846 506898 418888 507134
rect 418568 506866 418888 506898
rect 449288 507454 449608 507486
rect 449288 507218 449330 507454
rect 449566 507218 449608 507454
rect 449288 507134 449608 507218
rect 449288 506898 449330 507134
rect 449566 506898 449608 507134
rect 449288 506866 449608 506898
rect 480008 507454 480328 507486
rect 480008 507218 480050 507454
rect 480286 507218 480328 507454
rect 480008 507134 480328 507218
rect 480008 506898 480050 507134
rect 480286 506898 480328 507134
rect 480008 506866 480328 506898
rect 510728 507454 511048 507486
rect 510728 507218 510770 507454
rect 511006 507218 511048 507454
rect 510728 507134 511048 507218
rect 510728 506898 510770 507134
rect 511006 506898 511048 507134
rect 510728 506866 511048 506898
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 34568 489454 34888 489486
rect 34568 489218 34610 489454
rect 34846 489218 34888 489454
rect 34568 489134 34888 489218
rect 34568 488898 34610 489134
rect 34846 488898 34888 489134
rect 34568 488866 34888 488898
rect 65288 489454 65608 489486
rect 65288 489218 65330 489454
rect 65566 489218 65608 489454
rect 65288 489134 65608 489218
rect 65288 488898 65330 489134
rect 65566 488898 65608 489134
rect 65288 488866 65608 488898
rect 96008 489454 96328 489486
rect 96008 489218 96050 489454
rect 96286 489218 96328 489454
rect 96008 489134 96328 489218
rect 96008 488898 96050 489134
rect 96286 488898 96328 489134
rect 96008 488866 96328 488898
rect 126728 489454 127048 489486
rect 126728 489218 126770 489454
rect 127006 489218 127048 489454
rect 126728 489134 127048 489218
rect 126728 488898 126770 489134
rect 127006 488898 127048 489134
rect 126728 488866 127048 488898
rect 157448 489454 157768 489486
rect 157448 489218 157490 489454
rect 157726 489218 157768 489454
rect 157448 489134 157768 489218
rect 157448 488898 157490 489134
rect 157726 488898 157768 489134
rect 157448 488866 157768 488898
rect 188168 489454 188488 489486
rect 188168 489218 188210 489454
rect 188446 489218 188488 489454
rect 188168 489134 188488 489218
rect 188168 488898 188210 489134
rect 188446 488898 188488 489134
rect 188168 488866 188488 488898
rect 218888 489454 219208 489486
rect 218888 489218 218930 489454
rect 219166 489218 219208 489454
rect 218888 489134 219208 489218
rect 218888 488898 218930 489134
rect 219166 488898 219208 489134
rect 218888 488866 219208 488898
rect 249608 489454 249928 489486
rect 249608 489218 249650 489454
rect 249886 489218 249928 489454
rect 249608 489134 249928 489218
rect 249608 488898 249650 489134
rect 249886 488898 249928 489134
rect 249608 488866 249928 488898
rect 280328 489454 280648 489486
rect 280328 489218 280370 489454
rect 280606 489218 280648 489454
rect 280328 489134 280648 489218
rect 280328 488898 280370 489134
rect 280606 488898 280648 489134
rect 280328 488866 280648 488898
rect 311048 489454 311368 489486
rect 311048 489218 311090 489454
rect 311326 489218 311368 489454
rect 311048 489134 311368 489218
rect 311048 488898 311090 489134
rect 311326 488898 311368 489134
rect 311048 488866 311368 488898
rect 341768 489454 342088 489486
rect 341768 489218 341810 489454
rect 342046 489218 342088 489454
rect 341768 489134 342088 489218
rect 341768 488898 341810 489134
rect 342046 488898 342088 489134
rect 341768 488866 342088 488898
rect 372488 489454 372808 489486
rect 372488 489218 372530 489454
rect 372766 489218 372808 489454
rect 372488 489134 372808 489218
rect 372488 488898 372530 489134
rect 372766 488898 372808 489134
rect 372488 488866 372808 488898
rect 403208 489454 403528 489486
rect 403208 489218 403250 489454
rect 403486 489218 403528 489454
rect 403208 489134 403528 489218
rect 403208 488898 403250 489134
rect 403486 488898 403528 489134
rect 403208 488866 403528 488898
rect 433928 489454 434248 489486
rect 433928 489218 433970 489454
rect 434206 489218 434248 489454
rect 433928 489134 434248 489218
rect 433928 488898 433970 489134
rect 434206 488898 434248 489134
rect 433928 488866 434248 488898
rect 464648 489454 464968 489486
rect 464648 489218 464690 489454
rect 464926 489218 464968 489454
rect 464648 489134 464968 489218
rect 464648 488898 464690 489134
rect 464926 488898 464968 489134
rect 464648 488866 464968 488898
rect 495368 489454 495688 489486
rect 495368 489218 495410 489454
rect 495646 489218 495688 489454
rect 495368 489134 495688 489218
rect 495368 488898 495410 489134
rect 495646 488898 495688 489134
rect 495368 488866 495688 488898
rect 526088 489454 526408 489486
rect 526088 489218 526130 489454
rect 526366 489218 526408 489454
rect 526088 489134 526408 489218
rect 526088 488898 526130 489134
rect 526366 488898 526408 489134
rect 526088 488866 526408 488898
rect 19208 471454 19528 471486
rect 19208 471218 19250 471454
rect 19486 471218 19528 471454
rect 19208 471134 19528 471218
rect 19208 470898 19250 471134
rect 19486 470898 19528 471134
rect 19208 470866 19528 470898
rect 49928 471454 50248 471486
rect 49928 471218 49970 471454
rect 50206 471218 50248 471454
rect 49928 471134 50248 471218
rect 49928 470898 49970 471134
rect 50206 470898 50248 471134
rect 49928 470866 50248 470898
rect 80648 471454 80968 471486
rect 80648 471218 80690 471454
rect 80926 471218 80968 471454
rect 80648 471134 80968 471218
rect 80648 470898 80690 471134
rect 80926 470898 80968 471134
rect 80648 470866 80968 470898
rect 111368 471454 111688 471486
rect 111368 471218 111410 471454
rect 111646 471218 111688 471454
rect 111368 471134 111688 471218
rect 111368 470898 111410 471134
rect 111646 470898 111688 471134
rect 111368 470866 111688 470898
rect 142088 471454 142408 471486
rect 142088 471218 142130 471454
rect 142366 471218 142408 471454
rect 142088 471134 142408 471218
rect 142088 470898 142130 471134
rect 142366 470898 142408 471134
rect 142088 470866 142408 470898
rect 172808 471454 173128 471486
rect 172808 471218 172850 471454
rect 173086 471218 173128 471454
rect 172808 471134 173128 471218
rect 172808 470898 172850 471134
rect 173086 470898 173128 471134
rect 172808 470866 173128 470898
rect 203528 471454 203848 471486
rect 203528 471218 203570 471454
rect 203806 471218 203848 471454
rect 203528 471134 203848 471218
rect 203528 470898 203570 471134
rect 203806 470898 203848 471134
rect 203528 470866 203848 470898
rect 234248 471454 234568 471486
rect 234248 471218 234290 471454
rect 234526 471218 234568 471454
rect 234248 471134 234568 471218
rect 234248 470898 234290 471134
rect 234526 470898 234568 471134
rect 234248 470866 234568 470898
rect 264968 471454 265288 471486
rect 264968 471218 265010 471454
rect 265246 471218 265288 471454
rect 264968 471134 265288 471218
rect 264968 470898 265010 471134
rect 265246 470898 265288 471134
rect 264968 470866 265288 470898
rect 295688 471454 296008 471486
rect 295688 471218 295730 471454
rect 295966 471218 296008 471454
rect 295688 471134 296008 471218
rect 295688 470898 295730 471134
rect 295966 470898 296008 471134
rect 295688 470866 296008 470898
rect 326408 471454 326728 471486
rect 326408 471218 326450 471454
rect 326686 471218 326728 471454
rect 326408 471134 326728 471218
rect 326408 470898 326450 471134
rect 326686 470898 326728 471134
rect 326408 470866 326728 470898
rect 357128 471454 357448 471486
rect 357128 471218 357170 471454
rect 357406 471218 357448 471454
rect 357128 471134 357448 471218
rect 357128 470898 357170 471134
rect 357406 470898 357448 471134
rect 357128 470866 357448 470898
rect 387848 471454 388168 471486
rect 387848 471218 387890 471454
rect 388126 471218 388168 471454
rect 387848 471134 388168 471218
rect 387848 470898 387890 471134
rect 388126 470898 388168 471134
rect 387848 470866 388168 470898
rect 418568 471454 418888 471486
rect 418568 471218 418610 471454
rect 418846 471218 418888 471454
rect 418568 471134 418888 471218
rect 418568 470898 418610 471134
rect 418846 470898 418888 471134
rect 418568 470866 418888 470898
rect 449288 471454 449608 471486
rect 449288 471218 449330 471454
rect 449566 471218 449608 471454
rect 449288 471134 449608 471218
rect 449288 470898 449330 471134
rect 449566 470898 449608 471134
rect 449288 470866 449608 470898
rect 480008 471454 480328 471486
rect 480008 471218 480050 471454
rect 480286 471218 480328 471454
rect 480008 471134 480328 471218
rect 480008 470898 480050 471134
rect 480286 470898 480328 471134
rect 480008 470866 480328 470898
rect 510728 471454 511048 471486
rect 510728 471218 510770 471454
rect 511006 471218 511048 471454
rect 510728 471134 511048 471218
rect 510728 470898 510770 471134
rect 511006 470898 511048 471134
rect 510728 470866 511048 470898
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 34568 453454 34888 453486
rect 34568 453218 34610 453454
rect 34846 453218 34888 453454
rect 34568 453134 34888 453218
rect 34568 452898 34610 453134
rect 34846 452898 34888 453134
rect 34568 452866 34888 452898
rect 65288 453454 65608 453486
rect 65288 453218 65330 453454
rect 65566 453218 65608 453454
rect 65288 453134 65608 453218
rect 65288 452898 65330 453134
rect 65566 452898 65608 453134
rect 65288 452866 65608 452898
rect 96008 453454 96328 453486
rect 96008 453218 96050 453454
rect 96286 453218 96328 453454
rect 96008 453134 96328 453218
rect 96008 452898 96050 453134
rect 96286 452898 96328 453134
rect 96008 452866 96328 452898
rect 126728 453454 127048 453486
rect 126728 453218 126770 453454
rect 127006 453218 127048 453454
rect 126728 453134 127048 453218
rect 126728 452898 126770 453134
rect 127006 452898 127048 453134
rect 126728 452866 127048 452898
rect 157448 453454 157768 453486
rect 157448 453218 157490 453454
rect 157726 453218 157768 453454
rect 157448 453134 157768 453218
rect 157448 452898 157490 453134
rect 157726 452898 157768 453134
rect 157448 452866 157768 452898
rect 188168 453454 188488 453486
rect 188168 453218 188210 453454
rect 188446 453218 188488 453454
rect 188168 453134 188488 453218
rect 188168 452898 188210 453134
rect 188446 452898 188488 453134
rect 188168 452866 188488 452898
rect 218888 453454 219208 453486
rect 218888 453218 218930 453454
rect 219166 453218 219208 453454
rect 218888 453134 219208 453218
rect 218888 452898 218930 453134
rect 219166 452898 219208 453134
rect 218888 452866 219208 452898
rect 249608 453454 249928 453486
rect 249608 453218 249650 453454
rect 249886 453218 249928 453454
rect 249608 453134 249928 453218
rect 249608 452898 249650 453134
rect 249886 452898 249928 453134
rect 249608 452866 249928 452898
rect 280328 453454 280648 453486
rect 280328 453218 280370 453454
rect 280606 453218 280648 453454
rect 280328 453134 280648 453218
rect 280328 452898 280370 453134
rect 280606 452898 280648 453134
rect 280328 452866 280648 452898
rect 311048 453454 311368 453486
rect 311048 453218 311090 453454
rect 311326 453218 311368 453454
rect 311048 453134 311368 453218
rect 311048 452898 311090 453134
rect 311326 452898 311368 453134
rect 311048 452866 311368 452898
rect 341768 453454 342088 453486
rect 341768 453218 341810 453454
rect 342046 453218 342088 453454
rect 341768 453134 342088 453218
rect 341768 452898 341810 453134
rect 342046 452898 342088 453134
rect 341768 452866 342088 452898
rect 372488 453454 372808 453486
rect 372488 453218 372530 453454
rect 372766 453218 372808 453454
rect 372488 453134 372808 453218
rect 372488 452898 372530 453134
rect 372766 452898 372808 453134
rect 372488 452866 372808 452898
rect 403208 453454 403528 453486
rect 403208 453218 403250 453454
rect 403486 453218 403528 453454
rect 403208 453134 403528 453218
rect 403208 452898 403250 453134
rect 403486 452898 403528 453134
rect 403208 452866 403528 452898
rect 433928 453454 434248 453486
rect 433928 453218 433970 453454
rect 434206 453218 434248 453454
rect 433928 453134 434248 453218
rect 433928 452898 433970 453134
rect 434206 452898 434248 453134
rect 433928 452866 434248 452898
rect 464648 453454 464968 453486
rect 464648 453218 464690 453454
rect 464926 453218 464968 453454
rect 464648 453134 464968 453218
rect 464648 452898 464690 453134
rect 464926 452898 464968 453134
rect 464648 452866 464968 452898
rect 495368 453454 495688 453486
rect 495368 453218 495410 453454
rect 495646 453218 495688 453454
rect 495368 453134 495688 453218
rect 495368 452898 495410 453134
rect 495646 452898 495688 453134
rect 495368 452866 495688 452898
rect 526088 453454 526408 453486
rect 526088 453218 526130 453454
rect 526366 453218 526408 453454
rect 526088 453134 526408 453218
rect 526088 452898 526130 453134
rect 526366 452898 526408 453134
rect 526088 452866 526408 452898
rect 19208 435454 19528 435486
rect 19208 435218 19250 435454
rect 19486 435218 19528 435454
rect 19208 435134 19528 435218
rect 19208 434898 19250 435134
rect 19486 434898 19528 435134
rect 19208 434866 19528 434898
rect 49928 435454 50248 435486
rect 49928 435218 49970 435454
rect 50206 435218 50248 435454
rect 49928 435134 50248 435218
rect 49928 434898 49970 435134
rect 50206 434898 50248 435134
rect 49928 434866 50248 434898
rect 80648 435454 80968 435486
rect 80648 435218 80690 435454
rect 80926 435218 80968 435454
rect 80648 435134 80968 435218
rect 80648 434898 80690 435134
rect 80926 434898 80968 435134
rect 80648 434866 80968 434898
rect 111368 435454 111688 435486
rect 111368 435218 111410 435454
rect 111646 435218 111688 435454
rect 111368 435134 111688 435218
rect 111368 434898 111410 435134
rect 111646 434898 111688 435134
rect 111368 434866 111688 434898
rect 142088 435454 142408 435486
rect 142088 435218 142130 435454
rect 142366 435218 142408 435454
rect 142088 435134 142408 435218
rect 142088 434898 142130 435134
rect 142366 434898 142408 435134
rect 142088 434866 142408 434898
rect 172808 435454 173128 435486
rect 172808 435218 172850 435454
rect 173086 435218 173128 435454
rect 172808 435134 173128 435218
rect 172808 434898 172850 435134
rect 173086 434898 173128 435134
rect 172808 434866 173128 434898
rect 203528 435454 203848 435486
rect 203528 435218 203570 435454
rect 203806 435218 203848 435454
rect 203528 435134 203848 435218
rect 203528 434898 203570 435134
rect 203806 434898 203848 435134
rect 203528 434866 203848 434898
rect 234248 435454 234568 435486
rect 234248 435218 234290 435454
rect 234526 435218 234568 435454
rect 234248 435134 234568 435218
rect 234248 434898 234290 435134
rect 234526 434898 234568 435134
rect 234248 434866 234568 434898
rect 264968 435454 265288 435486
rect 264968 435218 265010 435454
rect 265246 435218 265288 435454
rect 264968 435134 265288 435218
rect 264968 434898 265010 435134
rect 265246 434898 265288 435134
rect 264968 434866 265288 434898
rect 295688 435454 296008 435486
rect 295688 435218 295730 435454
rect 295966 435218 296008 435454
rect 295688 435134 296008 435218
rect 295688 434898 295730 435134
rect 295966 434898 296008 435134
rect 295688 434866 296008 434898
rect 326408 435454 326728 435486
rect 326408 435218 326450 435454
rect 326686 435218 326728 435454
rect 326408 435134 326728 435218
rect 326408 434898 326450 435134
rect 326686 434898 326728 435134
rect 326408 434866 326728 434898
rect 357128 435454 357448 435486
rect 357128 435218 357170 435454
rect 357406 435218 357448 435454
rect 357128 435134 357448 435218
rect 357128 434898 357170 435134
rect 357406 434898 357448 435134
rect 357128 434866 357448 434898
rect 387848 435454 388168 435486
rect 387848 435218 387890 435454
rect 388126 435218 388168 435454
rect 387848 435134 388168 435218
rect 387848 434898 387890 435134
rect 388126 434898 388168 435134
rect 387848 434866 388168 434898
rect 418568 435454 418888 435486
rect 418568 435218 418610 435454
rect 418846 435218 418888 435454
rect 418568 435134 418888 435218
rect 418568 434898 418610 435134
rect 418846 434898 418888 435134
rect 418568 434866 418888 434898
rect 449288 435454 449608 435486
rect 449288 435218 449330 435454
rect 449566 435218 449608 435454
rect 449288 435134 449608 435218
rect 449288 434898 449330 435134
rect 449566 434898 449608 435134
rect 449288 434866 449608 434898
rect 480008 435454 480328 435486
rect 480008 435218 480050 435454
rect 480286 435218 480328 435454
rect 480008 435134 480328 435218
rect 480008 434898 480050 435134
rect 480286 434898 480328 435134
rect 480008 434866 480328 434898
rect 510728 435454 511048 435486
rect 510728 435218 510770 435454
rect 511006 435218 511048 435454
rect 510728 435134 511048 435218
rect 510728 434898 510770 435134
rect 511006 434898 511048 435134
rect 510728 434866 511048 434898
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 34568 417454 34888 417486
rect 34568 417218 34610 417454
rect 34846 417218 34888 417454
rect 34568 417134 34888 417218
rect 34568 416898 34610 417134
rect 34846 416898 34888 417134
rect 34568 416866 34888 416898
rect 65288 417454 65608 417486
rect 65288 417218 65330 417454
rect 65566 417218 65608 417454
rect 65288 417134 65608 417218
rect 65288 416898 65330 417134
rect 65566 416898 65608 417134
rect 65288 416866 65608 416898
rect 96008 417454 96328 417486
rect 96008 417218 96050 417454
rect 96286 417218 96328 417454
rect 96008 417134 96328 417218
rect 96008 416898 96050 417134
rect 96286 416898 96328 417134
rect 96008 416866 96328 416898
rect 126728 417454 127048 417486
rect 126728 417218 126770 417454
rect 127006 417218 127048 417454
rect 126728 417134 127048 417218
rect 126728 416898 126770 417134
rect 127006 416898 127048 417134
rect 126728 416866 127048 416898
rect 157448 417454 157768 417486
rect 157448 417218 157490 417454
rect 157726 417218 157768 417454
rect 157448 417134 157768 417218
rect 157448 416898 157490 417134
rect 157726 416898 157768 417134
rect 157448 416866 157768 416898
rect 188168 417454 188488 417486
rect 188168 417218 188210 417454
rect 188446 417218 188488 417454
rect 188168 417134 188488 417218
rect 188168 416898 188210 417134
rect 188446 416898 188488 417134
rect 188168 416866 188488 416898
rect 218888 417454 219208 417486
rect 218888 417218 218930 417454
rect 219166 417218 219208 417454
rect 218888 417134 219208 417218
rect 218888 416898 218930 417134
rect 219166 416898 219208 417134
rect 218888 416866 219208 416898
rect 249608 417454 249928 417486
rect 249608 417218 249650 417454
rect 249886 417218 249928 417454
rect 249608 417134 249928 417218
rect 249608 416898 249650 417134
rect 249886 416898 249928 417134
rect 249608 416866 249928 416898
rect 280328 417454 280648 417486
rect 280328 417218 280370 417454
rect 280606 417218 280648 417454
rect 280328 417134 280648 417218
rect 280328 416898 280370 417134
rect 280606 416898 280648 417134
rect 280328 416866 280648 416898
rect 311048 417454 311368 417486
rect 311048 417218 311090 417454
rect 311326 417218 311368 417454
rect 311048 417134 311368 417218
rect 311048 416898 311090 417134
rect 311326 416898 311368 417134
rect 311048 416866 311368 416898
rect 341768 417454 342088 417486
rect 341768 417218 341810 417454
rect 342046 417218 342088 417454
rect 341768 417134 342088 417218
rect 341768 416898 341810 417134
rect 342046 416898 342088 417134
rect 341768 416866 342088 416898
rect 372488 417454 372808 417486
rect 372488 417218 372530 417454
rect 372766 417218 372808 417454
rect 372488 417134 372808 417218
rect 372488 416898 372530 417134
rect 372766 416898 372808 417134
rect 372488 416866 372808 416898
rect 403208 417454 403528 417486
rect 403208 417218 403250 417454
rect 403486 417218 403528 417454
rect 403208 417134 403528 417218
rect 403208 416898 403250 417134
rect 403486 416898 403528 417134
rect 403208 416866 403528 416898
rect 433928 417454 434248 417486
rect 433928 417218 433970 417454
rect 434206 417218 434248 417454
rect 433928 417134 434248 417218
rect 433928 416898 433970 417134
rect 434206 416898 434248 417134
rect 433928 416866 434248 416898
rect 464648 417454 464968 417486
rect 464648 417218 464690 417454
rect 464926 417218 464968 417454
rect 464648 417134 464968 417218
rect 464648 416898 464690 417134
rect 464926 416898 464968 417134
rect 464648 416866 464968 416898
rect 495368 417454 495688 417486
rect 495368 417218 495410 417454
rect 495646 417218 495688 417454
rect 495368 417134 495688 417218
rect 495368 416898 495410 417134
rect 495646 416898 495688 417134
rect 495368 416866 495688 416898
rect 526088 417454 526408 417486
rect 526088 417218 526130 417454
rect 526366 417218 526408 417454
rect 526088 417134 526408 417218
rect 526088 416898 526130 417134
rect 526366 416898 526408 417134
rect 526088 416866 526408 416898
rect 19208 399454 19528 399486
rect 19208 399218 19250 399454
rect 19486 399218 19528 399454
rect 19208 399134 19528 399218
rect 19208 398898 19250 399134
rect 19486 398898 19528 399134
rect 19208 398866 19528 398898
rect 49928 399454 50248 399486
rect 49928 399218 49970 399454
rect 50206 399218 50248 399454
rect 49928 399134 50248 399218
rect 49928 398898 49970 399134
rect 50206 398898 50248 399134
rect 49928 398866 50248 398898
rect 80648 399454 80968 399486
rect 80648 399218 80690 399454
rect 80926 399218 80968 399454
rect 80648 399134 80968 399218
rect 80648 398898 80690 399134
rect 80926 398898 80968 399134
rect 80648 398866 80968 398898
rect 111368 399454 111688 399486
rect 111368 399218 111410 399454
rect 111646 399218 111688 399454
rect 111368 399134 111688 399218
rect 111368 398898 111410 399134
rect 111646 398898 111688 399134
rect 111368 398866 111688 398898
rect 142088 399454 142408 399486
rect 142088 399218 142130 399454
rect 142366 399218 142408 399454
rect 142088 399134 142408 399218
rect 142088 398898 142130 399134
rect 142366 398898 142408 399134
rect 142088 398866 142408 398898
rect 172808 399454 173128 399486
rect 172808 399218 172850 399454
rect 173086 399218 173128 399454
rect 172808 399134 173128 399218
rect 172808 398898 172850 399134
rect 173086 398898 173128 399134
rect 172808 398866 173128 398898
rect 203528 399454 203848 399486
rect 203528 399218 203570 399454
rect 203806 399218 203848 399454
rect 203528 399134 203848 399218
rect 203528 398898 203570 399134
rect 203806 398898 203848 399134
rect 203528 398866 203848 398898
rect 234248 399454 234568 399486
rect 234248 399218 234290 399454
rect 234526 399218 234568 399454
rect 234248 399134 234568 399218
rect 234248 398898 234290 399134
rect 234526 398898 234568 399134
rect 234248 398866 234568 398898
rect 264968 399454 265288 399486
rect 264968 399218 265010 399454
rect 265246 399218 265288 399454
rect 264968 399134 265288 399218
rect 264968 398898 265010 399134
rect 265246 398898 265288 399134
rect 264968 398866 265288 398898
rect 295688 399454 296008 399486
rect 295688 399218 295730 399454
rect 295966 399218 296008 399454
rect 295688 399134 296008 399218
rect 295688 398898 295730 399134
rect 295966 398898 296008 399134
rect 295688 398866 296008 398898
rect 326408 399454 326728 399486
rect 326408 399218 326450 399454
rect 326686 399218 326728 399454
rect 326408 399134 326728 399218
rect 326408 398898 326450 399134
rect 326686 398898 326728 399134
rect 326408 398866 326728 398898
rect 357128 399454 357448 399486
rect 357128 399218 357170 399454
rect 357406 399218 357448 399454
rect 357128 399134 357448 399218
rect 357128 398898 357170 399134
rect 357406 398898 357448 399134
rect 357128 398866 357448 398898
rect 387848 399454 388168 399486
rect 387848 399218 387890 399454
rect 388126 399218 388168 399454
rect 387848 399134 388168 399218
rect 387848 398898 387890 399134
rect 388126 398898 388168 399134
rect 387848 398866 388168 398898
rect 418568 399454 418888 399486
rect 418568 399218 418610 399454
rect 418846 399218 418888 399454
rect 418568 399134 418888 399218
rect 418568 398898 418610 399134
rect 418846 398898 418888 399134
rect 418568 398866 418888 398898
rect 449288 399454 449608 399486
rect 449288 399218 449330 399454
rect 449566 399218 449608 399454
rect 449288 399134 449608 399218
rect 449288 398898 449330 399134
rect 449566 398898 449608 399134
rect 449288 398866 449608 398898
rect 480008 399454 480328 399486
rect 480008 399218 480050 399454
rect 480286 399218 480328 399454
rect 480008 399134 480328 399218
rect 480008 398898 480050 399134
rect 480286 398898 480328 399134
rect 480008 398866 480328 398898
rect 510728 399454 511048 399486
rect 510728 399218 510770 399454
rect 511006 399218 511048 399454
rect 510728 399134 511048 399218
rect 510728 398898 510770 399134
rect 511006 398898 511048 399134
rect 510728 398866 511048 398898
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 34568 381454 34888 381486
rect 34568 381218 34610 381454
rect 34846 381218 34888 381454
rect 34568 381134 34888 381218
rect 34568 380898 34610 381134
rect 34846 380898 34888 381134
rect 34568 380866 34888 380898
rect 65288 381454 65608 381486
rect 65288 381218 65330 381454
rect 65566 381218 65608 381454
rect 65288 381134 65608 381218
rect 65288 380898 65330 381134
rect 65566 380898 65608 381134
rect 65288 380866 65608 380898
rect 96008 381454 96328 381486
rect 96008 381218 96050 381454
rect 96286 381218 96328 381454
rect 96008 381134 96328 381218
rect 96008 380898 96050 381134
rect 96286 380898 96328 381134
rect 96008 380866 96328 380898
rect 126728 381454 127048 381486
rect 126728 381218 126770 381454
rect 127006 381218 127048 381454
rect 126728 381134 127048 381218
rect 126728 380898 126770 381134
rect 127006 380898 127048 381134
rect 126728 380866 127048 380898
rect 157448 381454 157768 381486
rect 157448 381218 157490 381454
rect 157726 381218 157768 381454
rect 157448 381134 157768 381218
rect 157448 380898 157490 381134
rect 157726 380898 157768 381134
rect 157448 380866 157768 380898
rect 188168 381454 188488 381486
rect 188168 381218 188210 381454
rect 188446 381218 188488 381454
rect 188168 381134 188488 381218
rect 188168 380898 188210 381134
rect 188446 380898 188488 381134
rect 188168 380866 188488 380898
rect 218888 381454 219208 381486
rect 218888 381218 218930 381454
rect 219166 381218 219208 381454
rect 218888 381134 219208 381218
rect 218888 380898 218930 381134
rect 219166 380898 219208 381134
rect 218888 380866 219208 380898
rect 249608 381454 249928 381486
rect 249608 381218 249650 381454
rect 249886 381218 249928 381454
rect 249608 381134 249928 381218
rect 249608 380898 249650 381134
rect 249886 380898 249928 381134
rect 249608 380866 249928 380898
rect 280328 381454 280648 381486
rect 280328 381218 280370 381454
rect 280606 381218 280648 381454
rect 280328 381134 280648 381218
rect 280328 380898 280370 381134
rect 280606 380898 280648 381134
rect 280328 380866 280648 380898
rect 311048 381454 311368 381486
rect 311048 381218 311090 381454
rect 311326 381218 311368 381454
rect 311048 381134 311368 381218
rect 311048 380898 311090 381134
rect 311326 380898 311368 381134
rect 311048 380866 311368 380898
rect 341768 381454 342088 381486
rect 341768 381218 341810 381454
rect 342046 381218 342088 381454
rect 341768 381134 342088 381218
rect 341768 380898 341810 381134
rect 342046 380898 342088 381134
rect 341768 380866 342088 380898
rect 372488 381454 372808 381486
rect 372488 381218 372530 381454
rect 372766 381218 372808 381454
rect 372488 381134 372808 381218
rect 372488 380898 372530 381134
rect 372766 380898 372808 381134
rect 372488 380866 372808 380898
rect 403208 381454 403528 381486
rect 403208 381218 403250 381454
rect 403486 381218 403528 381454
rect 403208 381134 403528 381218
rect 403208 380898 403250 381134
rect 403486 380898 403528 381134
rect 403208 380866 403528 380898
rect 433928 381454 434248 381486
rect 433928 381218 433970 381454
rect 434206 381218 434248 381454
rect 433928 381134 434248 381218
rect 433928 380898 433970 381134
rect 434206 380898 434248 381134
rect 433928 380866 434248 380898
rect 464648 381454 464968 381486
rect 464648 381218 464690 381454
rect 464926 381218 464968 381454
rect 464648 381134 464968 381218
rect 464648 380898 464690 381134
rect 464926 380898 464968 381134
rect 464648 380866 464968 380898
rect 495368 381454 495688 381486
rect 495368 381218 495410 381454
rect 495646 381218 495688 381454
rect 495368 381134 495688 381218
rect 495368 380898 495410 381134
rect 495646 380898 495688 381134
rect 495368 380866 495688 380898
rect 526088 381454 526408 381486
rect 526088 381218 526130 381454
rect 526366 381218 526408 381454
rect 526088 381134 526408 381218
rect 526088 380898 526130 381134
rect 526366 380898 526408 381134
rect 526088 380866 526408 380898
rect 19208 363454 19528 363486
rect 19208 363218 19250 363454
rect 19486 363218 19528 363454
rect 19208 363134 19528 363218
rect 19208 362898 19250 363134
rect 19486 362898 19528 363134
rect 19208 362866 19528 362898
rect 49928 363454 50248 363486
rect 49928 363218 49970 363454
rect 50206 363218 50248 363454
rect 49928 363134 50248 363218
rect 49928 362898 49970 363134
rect 50206 362898 50248 363134
rect 49928 362866 50248 362898
rect 80648 363454 80968 363486
rect 80648 363218 80690 363454
rect 80926 363218 80968 363454
rect 80648 363134 80968 363218
rect 80648 362898 80690 363134
rect 80926 362898 80968 363134
rect 80648 362866 80968 362898
rect 111368 363454 111688 363486
rect 111368 363218 111410 363454
rect 111646 363218 111688 363454
rect 111368 363134 111688 363218
rect 111368 362898 111410 363134
rect 111646 362898 111688 363134
rect 111368 362866 111688 362898
rect 142088 363454 142408 363486
rect 142088 363218 142130 363454
rect 142366 363218 142408 363454
rect 142088 363134 142408 363218
rect 142088 362898 142130 363134
rect 142366 362898 142408 363134
rect 142088 362866 142408 362898
rect 172808 363454 173128 363486
rect 172808 363218 172850 363454
rect 173086 363218 173128 363454
rect 172808 363134 173128 363218
rect 172808 362898 172850 363134
rect 173086 362898 173128 363134
rect 172808 362866 173128 362898
rect 203528 363454 203848 363486
rect 203528 363218 203570 363454
rect 203806 363218 203848 363454
rect 203528 363134 203848 363218
rect 203528 362898 203570 363134
rect 203806 362898 203848 363134
rect 203528 362866 203848 362898
rect 234248 363454 234568 363486
rect 234248 363218 234290 363454
rect 234526 363218 234568 363454
rect 234248 363134 234568 363218
rect 234248 362898 234290 363134
rect 234526 362898 234568 363134
rect 234248 362866 234568 362898
rect 264968 363454 265288 363486
rect 264968 363218 265010 363454
rect 265246 363218 265288 363454
rect 264968 363134 265288 363218
rect 264968 362898 265010 363134
rect 265246 362898 265288 363134
rect 264968 362866 265288 362898
rect 295688 363454 296008 363486
rect 295688 363218 295730 363454
rect 295966 363218 296008 363454
rect 295688 363134 296008 363218
rect 295688 362898 295730 363134
rect 295966 362898 296008 363134
rect 295688 362866 296008 362898
rect 326408 363454 326728 363486
rect 326408 363218 326450 363454
rect 326686 363218 326728 363454
rect 326408 363134 326728 363218
rect 326408 362898 326450 363134
rect 326686 362898 326728 363134
rect 326408 362866 326728 362898
rect 357128 363454 357448 363486
rect 357128 363218 357170 363454
rect 357406 363218 357448 363454
rect 357128 363134 357448 363218
rect 357128 362898 357170 363134
rect 357406 362898 357448 363134
rect 357128 362866 357448 362898
rect 387848 363454 388168 363486
rect 387848 363218 387890 363454
rect 388126 363218 388168 363454
rect 387848 363134 388168 363218
rect 387848 362898 387890 363134
rect 388126 362898 388168 363134
rect 387848 362866 388168 362898
rect 418568 363454 418888 363486
rect 418568 363218 418610 363454
rect 418846 363218 418888 363454
rect 418568 363134 418888 363218
rect 418568 362898 418610 363134
rect 418846 362898 418888 363134
rect 418568 362866 418888 362898
rect 449288 363454 449608 363486
rect 449288 363218 449330 363454
rect 449566 363218 449608 363454
rect 449288 363134 449608 363218
rect 449288 362898 449330 363134
rect 449566 362898 449608 363134
rect 449288 362866 449608 362898
rect 480008 363454 480328 363486
rect 480008 363218 480050 363454
rect 480286 363218 480328 363454
rect 480008 363134 480328 363218
rect 480008 362898 480050 363134
rect 480286 362898 480328 363134
rect 480008 362866 480328 362898
rect 510728 363454 511048 363486
rect 510728 363218 510770 363454
rect 511006 363218 511048 363454
rect 510728 363134 511048 363218
rect 510728 362898 510770 363134
rect 511006 362898 511048 363134
rect 510728 362866 511048 362898
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 34568 345454 34888 345486
rect 34568 345218 34610 345454
rect 34846 345218 34888 345454
rect 34568 345134 34888 345218
rect 34568 344898 34610 345134
rect 34846 344898 34888 345134
rect 34568 344866 34888 344898
rect 65288 345454 65608 345486
rect 65288 345218 65330 345454
rect 65566 345218 65608 345454
rect 65288 345134 65608 345218
rect 65288 344898 65330 345134
rect 65566 344898 65608 345134
rect 65288 344866 65608 344898
rect 96008 345454 96328 345486
rect 96008 345218 96050 345454
rect 96286 345218 96328 345454
rect 96008 345134 96328 345218
rect 96008 344898 96050 345134
rect 96286 344898 96328 345134
rect 96008 344866 96328 344898
rect 126728 345454 127048 345486
rect 126728 345218 126770 345454
rect 127006 345218 127048 345454
rect 126728 345134 127048 345218
rect 126728 344898 126770 345134
rect 127006 344898 127048 345134
rect 126728 344866 127048 344898
rect 157448 345454 157768 345486
rect 157448 345218 157490 345454
rect 157726 345218 157768 345454
rect 157448 345134 157768 345218
rect 157448 344898 157490 345134
rect 157726 344898 157768 345134
rect 157448 344866 157768 344898
rect 188168 345454 188488 345486
rect 188168 345218 188210 345454
rect 188446 345218 188488 345454
rect 188168 345134 188488 345218
rect 188168 344898 188210 345134
rect 188446 344898 188488 345134
rect 188168 344866 188488 344898
rect 218888 345454 219208 345486
rect 218888 345218 218930 345454
rect 219166 345218 219208 345454
rect 218888 345134 219208 345218
rect 218888 344898 218930 345134
rect 219166 344898 219208 345134
rect 218888 344866 219208 344898
rect 249608 345454 249928 345486
rect 249608 345218 249650 345454
rect 249886 345218 249928 345454
rect 249608 345134 249928 345218
rect 249608 344898 249650 345134
rect 249886 344898 249928 345134
rect 249608 344866 249928 344898
rect 280328 345454 280648 345486
rect 280328 345218 280370 345454
rect 280606 345218 280648 345454
rect 280328 345134 280648 345218
rect 280328 344898 280370 345134
rect 280606 344898 280648 345134
rect 280328 344866 280648 344898
rect 311048 345454 311368 345486
rect 311048 345218 311090 345454
rect 311326 345218 311368 345454
rect 311048 345134 311368 345218
rect 311048 344898 311090 345134
rect 311326 344898 311368 345134
rect 311048 344866 311368 344898
rect 341768 345454 342088 345486
rect 341768 345218 341810 345454
rect 342046 345218 342088 345454
rect 341768 345134 342088 345218
rect 341768 344898 341810 345134
rect 342046 344898 342088 345134
rect 341768 344866 342088 344898
rect 372488 345454 372808 345486
rect 372488 345218 372530 345454
rect 372766 345218 372808 345454
rect 372488 345134 372808 345218
rect 372488 344898 372530 345134
rect 372766 344898 372808 345134
rect 372488 344866 372808 344898
rect 403208 345454 403528 345486
rect 403208 345218 403250 345454
rect 403486 345218 403528 345454
rect 403208 345134 403528 345218
rect 403208 344898 403250 345134
rect 403486 344898 403528 345134
rect 403208 344866 403528 344898
rect 433928 345454 434248 345486
rect 433928 345218 433970 345454
rect 434206 345218 434248 345454
rect 433928 345134 434248 345218
rect 433928 344898 433970 345134
rect 434206 344898 434248 345134
rect 433928 344866 434248 344898
rect 464648 345454 464968 345486
rect 464648 345218 464690 345454
rect 464926 345218 464968 345454
rect 464648 345134 464968 345218
rect 464648 344898 464690 345134
rect 464926 344898 464968 345134
rect 464648 344866 464968 344898
rect 495368 345454 495688 345486
rect 495368 345218 495410 345454
rect 495646 345218 495688 345454
rect 495368 345134 495688 345218
rect 495368 344898 495410 345134
rect 495646 344898 495688 345134
rect 495368 344866 495688 344898
rect 526088 345454 526408 345486
rect 526088 345218 526130 345454
rect 526366 345218 526408 345454
rect 526088 345134 526408 345218
rect 526088 344898 526130 345134
rect 526366 344898 526408 345134
rect 526088 344866 526408 344898
rect 19208 327454 19528 327486
rect 19208 327218 19250 327454
rect 19486 327218 19528 327454
rect 19208 327134 19528 327218
rect 19208 326898 19250 327134
rect 19486 326898 19528 327134
rect 19208 326866 19528 326898
rect 49928 327454 50248 327486
rect 49928 327218 49970 327454
rect 50206 327218 50248 327454
rect 49928 327134 50248 327218
rect 49928 326898 49970 327134
rect 50206 326898 50248 327134
rect 49928 326866 50248 326898
rect 80648 327454 80968 327486
rect 80648 327218 80690 327454
rect 80926 327218 80968 327454
rect 80648 327134 80968 327218
rect 80648 326898 80690 327134
rect 80926 326898 80968 327134
rect 80648 326866 80968 326898
rect 111368 327454 111688 327486
rect 111368 327218 111410 327454
rect 111646 327218 111688 327454
rect 111368 327134 111688 327218
rect 111368 326898 111410 327134
rect 111646 326898 111688 327134
rect 111368 326866 111688 326898
rect 142088 327454 142408 327486
rect 142088 327218 142130 327454
rect 142366 327218 142408 327454
rect 142088 327134 142408 327218
rect 142088 326898 142130 327134
rect 142366 326898 142408 327134
rect 142088 326866 142408 326898
rect 172808 327454 173128 327486
rect 172808 327218 172850 327454
rect 173086 327218 173128 327454
rect 172808 327134 173128 327218
rect 172808 326898 172850 327134
rect 173086 326898 173128 327134
rect 172808 326866 173128 326898
rect 203528 327454 203848 327486
rect 203528 327218 203570 327454
rect 203806 327218 203848 327454
rect 203528 327134 203848 327218
rect 203528 326898 203570 327134
rect 203806 326898 203848 327134
rect 203528 326866 203848 326898
rect 234248 327454 234568 327486
rect 234248 327218 234290 327454
rect 234526 327218 234568 327454
rect 234248 327134 234568 327218
rect 234248 326898 234290 327134
rect 234526 326898 234568 327134
rect 234248 326866 234568 326898
rect 264968 327454 265288 327486
rect 264968 327218 265010 327454
rect 265246 327218 265288 327454
rect 264968 327134 265288 327218
rect 264968 326898 265010 327134
rect 265246 326898 265288 327134
rect 264968 326866 265288 326898
rect 295688 327454 296008 327486
rect 295688 327218 295730 327454
rect 295966 327218 296008 327454
rect 295688 327134 296008 327218
rect 295688 326898 295730 327134
rect 295966 326898 296008 327134
rect 295688 326866 296008 326898
rect 326408 327454 326728 327486
rect 326408 327218 326450 327454
rect 326686 327218 326728 327454
rect 326408 327134 326728 327218
rect 326408 326898 326450 327134
rect 326686 326898 326728 327134
rect 326408 326866 326728 326898
rect 357128 327454 357448 327486
rect 357128 327218 357170 327454
rect 357406 327218 357448 327454
rect 357128 327134 357448 327218
rect 357128 326898 357170 327134
rect 357406 326898 357448 327134
rect 357128 326866 357448 326898
rect 387848 327454 388168 327486
rect 387848 327218 387890 327454
rect 388126 327218 388168 327454
rect 387848 327134 388168 327218
rect 387848 326898 387890 327134
rect 388126 326898 388168 327134
rect 387848 326866 388168 326898
rect 418568 327454 418888 327486
rect 418568 327218 418610 327454
rect 418846 327218 418888 327454
rect 418568 327134 418888 327218
rect 418568 326898 418610 327134
rect 418846 326898 418888 327134
rect 418568 326866 418888 326898
rect 449288 327454 449608 327486
rect 449288 327218 449330 327454
rect 449566 327218 449608 327454
rect 449288 327134 449608 327218
rect 449288 326898 449330 327134
rect 449566 326898 449608 327134
rect 449288 326866 449608 326898
rect 480008 327454 480328 327486
rect 480008 327218 480050 327454
rect 480286 327218 480328 327454
rect 480008 327134 480328 327218
rect 480008 326898 480050 327134
rect 480286 326898 480328 327134
rect 480008 326866 480328 326898
rect 510728 327454 511048 327486
rect 510728 327218 510770 327454
rect 511006 327218 511048 327454
rect 510728 327134 511048 327218
rect 510728 326898 510770 327134
rect 511006 326898 511048 327134
rect 510728 326866 511048 326898
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 34568 309454 34888 309486
rect 34568 309218 34610 309454
rect 34846 309218 34888 309454
rect 34568 309134 34888 309218
rect 34568 308898 34610 309134
rect 34846 308898 34888 309134
rect 34568 308866 34888 308898
rect 65288 309454 65608 309486
rect 65288 309218 65330 309454
rect 65566 309218 65608 309454
rect 65288 309134 65608 309218
rect 65288 308898 65330 309134
rect 65566 308898 65608 309134
rect 65288 308866 65608 308898
rect 96008 309454 96328 309486
rect 96008 309218 96050 309454
rect 96286 309218 96328 309454
rect 96008 309134 96328 309218
rect 96008 308898 96050 309134
rect 96286 308898 96328 309134
rect 96008 308866 96328 308898
rect 126728 309454 127048 309486
rect 126728 309218 126770 309454
rect 127006 309218 127048 309454
rect 126728 309134 127048 309218
rect 126728 308898 126770 309134
rect 127006 308898 127048 309134
rect 126728 308866 127048 308898
rect 157448 309454 157768 309486
rect 157448 309218 157490 309454
rect 157726 309218 157768 309454
rect 157448 309134 157768 309218
rect 157448 308898 157490 309134
rect 157726 308898 157768 309134
rect 157448 308866 157768 308898
rect 188168 309454 188488 309486
rect 188168 309218 188210 309454
rect 188446 309218 188488 309454
rect 188168 309134 188488 309218
rect 188168 308898 188210 309134
rect 188446 308898 188488 309134
rect 188168 308866 188488 308898
rect 218888 309454 219208 309486
rect 218888 309218 218930 309454
rect 219166 309218 219208 309454
rect 218888 309134 219208 309218
rect 218888 308898 218930 309134
rect 219166 308898 219208 309134
rect 218888 308866 219208 308898
rect 249608 309454 249928 309486
rect 249608 309218 249650 309454
rect 249886 309218 249928 309454
rect 249608 309134 249928 309218
rect 249608 308898 249650 309134
rect 249886 308898 249928 309134
rect 249608 308866 249928 308898
rect 280328 309454 280648 309486
rect 280328 309218 280370 309454
rect 280606 309218 280648 309454
rect 280328 309134 280648 309218
rect 280328 308898 280370 309134
rect 280606 308898 280648 309134
rect 280328 308866 280648 308898
rect 311048 309454 311368 309486
rect 311048 309218 311090 309454
rect 311326 309218 311368 309454
rect 311048 309134 311368 309218
rect 311048 308898 311090 309134
rect 311326 308898 311368 309134
rect 311048 308866 311368 308898
rect 341768 309454 342088 309486
rect 341768 309218 341810 309454
rect 342046 309218 342088 309454
rect 341768 309134 342088 309218
rect 341768 308898 341810 309134
rect 342046 308898 342088 309134
rect 341768 308866 342088 308898
rect 372488 309454 372808 309486
rect 372488 309218 372530 309454
rect 372766 309218 372808 309454
rect 372488 309134 372808 309218
rect 372488 308898 372530 309134
rect 372766 308898 372808 309134
rect 372488 308866 372808 308898
rect 403208 309454 403528 309486
rect 403208 309218 403250 309454
rect 403486 309218 403528 309454
rect 403208 309134 403528 309218
rect 403208 308898 403250 309134
rect 403486 308898 403528 309134
rect 403208 308866 403528 308898
rect 433928 309454 434248 309486
rect 433928 309218 433970 309454
rect 434206 309218 434248 309454
rect 433928 309134 434248 309218
rect 433928 308898 433970 309134
rect 434206 308898 434248 309134
rect 433928 308866 434248 308898
rect 464648 309454 464968 309486
rect 464648 309218 464690 309454
rect 464926 309218 464968 309454
rect 464648 309134 464968 309218
rect 464648 308898 464690 309134
rect 464926 308898 464968 309134
rect 464648 308866 464968 308898
rect 495368 309454 495688 309486
rect 495368 309218 495410 309454
rect 495646 309218 495688 309454
rect 495368 309134 495688 309218
rect 495368 308898 495410 309134
rect 495646 308898 495688 309134
rect 495368 308866 495688 308898
rect 526088 309454 526408 309486
rect 526088 309218 526130 309454
rect 526366 309218 526408 309454
rect 526088 309134 526408 309218
rect 526088 308898 526130 309134
rect 526366 308898 526408 309134
rect 526088 308866 526408 308898
rect 19208 291454 19528 291486
rect 19208 291218 19250 291454
rect 19486 291218 19528 291454
rect 19208 291134 19528 291218
rect 19208 290898 19250 291134
rect 19486 290898 19528 291134
rect 19208 290866 19528 290898
rect 49928 291454 50248 291486
rect 49928 291218 49970 291454
rect 50206 291218 50248 291454
rect 49928 291134 50248 291218
rect 49928 290898 49970 291134
rect 50206 290898 50248 291134
rect 49928 290866 50248 290898
rect 80648 291454 80968 291486
rect 80648 291218 80690 291454
rect 80926 291218 80968 291454
rect 80648 291134 80968 291218
rect 80648 290898 80690 291134
rect 80926 290898 80968 291134
rect 80648 290866 80968 290898
rect 111368 291454 111688 291486
rect 111368 291218 111410 291454
rect 111646 291218 111688 291454
rect 111368 291134 111688 291218
rect 111368 290898 111410 291134
rect 111646 290898 111688 291134
rect 111368 290866 111688 290898
rect 142088 291454 142408 291486
rect 142088 291218 142130 291454
rect 142366 291218 142408 291454
rect 142088 291134 142408 291218
rect 142088 290898 142130 291134
rect 142366 290898 142408 291134
rect 142088 290866 142408 290898
rect 172808 291454 173128 291486
rect 172808 291218 172850 291454
rect 173086 291218 173128 291454
rect 172808 291134 173128 291218
rect 172808 290898 172850 291134
rect 173086 290898 173128 291134
rect 172808 290866 173128 290898
rect 203528 291454 203848 291486
rect 203528 291218 203570 291454
rect 203806 291218 203848 291454
rect 203528 291134 203848 291218
rect 203528 290898 203570 291134
rect 203806 290898 203848 291134
rect 203528 290866 203848 290898
rect 234248 291454 234568 291486
rect 234248 291218 234290 291454
rect 234526 291218 234568 291454
rect 234248 291134 234568 291218
rect 234248 290898 234290 291134
rect 234526 290898 234568 291134
rect 234248 290866 234568 290898
rect 264968 291454 265288 291486
rect 264968 291218 265010 291454
rect 265246 291218 265288 291454
rect 264968 291134 265288 291218
rect 264968 290898 265010 291134
rect 265246 290898 265288 291134
rect 264968 290866 265288 290898
rect 295688 291454 296008 291486
rect 295688 291218 295730 291454
rect 295966 291218 296008 291454
rect 295688 291134 296008 291218
rect 295688 290898 295730 291134
rect 295966 290898 296008 291134
rect 295688 290866 296008 290898
rect 326408 291454 326728 291486
rect 326408 291218 326450 291454
rect 326686 291218 326728 291454
rect 326408 291134 326728 291218
rect 326408 290898 326450 291134
rect 326686 290898 326728 291134
rect 326408 290866 326728 290898
rect 357128 291454 357448 291486
rect 357128 291218 357170 291454
rect 357406 291218 357448 291454
rect 357128 291134 357448 291218
rect 357128 290898 357170 291134
rect 357406 290898 357448 291134
rect 357128 290866 357448 290898
rect 387848 291454 388168 291486
rect 387848 291218 387890 291454
rect 388126 291218 388168 291454
rect 387848 291134 388168 291218
rect 387848 290898 387890 291134
rect 388126 290898 388168 291134
rect 387848 290866 388168 290898
rect 418568 291454 418888 291486
rect 418568 291218 418610 291454
rect 418846 291218 418888 291454
rect 418568 291134 418888 291218
rect 418568 290898 418610 291134
rect 418846 290898 418888 291134
rect 418568 290866 418888 290898
rect 449288 291454 449608 291486
rect 449288 291218 449330 291454
rect 449566 291218 449608 291454
rect 449288 291134 449608 291218
rect 449288 290898 449330 291134
rect 449566 290898 449608 291134
rect 449288 290866 449608 290898
rect 480008 291454 480328 291486
rect 480008 291218 480050 291454
rect 480286 291218 480328 291454
rect 480008 291134 480328 291218
rect 480008 290898 480050 291134
rect 480286 290898 480328 291134
rect 480008 290866 480328 290898
rect 510728 291454 511048 291486
rect 510728 291218 510770 291454
rect 511006 291218 511048 291454
rect 510728 291134 511048 291218
rect 510728 290898 510770 291134
rect 511006 290898 511048 291134
rect 510728 290866 511048 290898
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 34568 273454 34888 273486
rect 34568 273218 34610 273454
rect 34846 273218 34888 273454
rect 34568 273134 34888 273218
rect 34568 272898 34610 273134
rect 34846 272898 34888 273134
rect 34568 272866 34888 272898
rect 65288 273454 65608 273486
rect 65288 273218 65330 273454
rect 65566 273218 65608 273454
rect 65288 273134 65608 273218
rect 65288 272898 65330 273134
rect 65566 272898 65608 273134
rect 65288 272866 65608 272898
rect 96008 273454 96328 273486
rect 96008 273218 96050 273454
rect 96286 273218 96328 273454
rect 96008 273134 96328 273218
rect 96008 272898 96050 273134
rect 96286 272898 96328 273134
rect 96008 272866 96328 272898
rect 126728 273454 127048 273486
rect 126728 273218 126770 273454
rect 127006 273218 127048 273454
rect 126728 273134 127048 273218
rect 126728 272898 126770 273134
rect 127006 272898 127048 273134
rect 126728 272866 127048 272898
rect 157448 273454 157768 273486
rect 157448 273218 157490 273454
rect 157726 273218 157768 273454
rect 157448 273134 157768 273218
rect 157448 272898 157490 273134
rect 157726 272898 157768 273134
rect 157448 272866 157768 272898
rect 188168 273454 188488 273486
rect 188168 273218 188210 273454
rect 188446 273218 188488 273454
rect 188168 273134 188488 273218
rect 188168 272898 188210 273134
rect 188446 272898 188488 273134
rect 188168 272866 188488 272898
rect 218888 273454 219208 273486
rect 218888 273218 218930 273454
rect 219166 273218 219208 273454
rect 218888 273134 219208 273218
rect 218888 272898 218930 273134
rect 219166 272898 219208 273134
rect 218888 272866 219208 272898
rect 249608 273454 249928 273486
rect 249608 273218 249650 273454
rect 249886 273218 249928 273454
rect 249608 273134 249928 273218
rect 249608 272898 249650 273134
rect 249886 272898 249928 273134
rect 249608 272866 249928 272898
rect 280328 273454 280648 273486
rect 280328 273218 280370 273454
rect 280606 273218 280648 273454
rect 280328 273134 280648 273218
rect 280328 272898 280370 273134
rect 280606 272898 280648 273134
rect 280328 272866 280648 272898
rect 311048 273454 311368 273486
rect 311048 273218 311090 273454
rect 311326 273218 311368 273454
rect 311048 273134 311368 273218
rect 311048 272898 311090 273134
rect 311326 272898 311368 273134
rect 311048 272866 311368 272898
rect 341768 273454 342088 273486
rect 341768 273218 341810 273454
rect 342046 273218 342088 273454
rect 341768 273134 342088 273218
rect 341768 272898 341810 273134
rect 342046 272898 342088 273134
rect 341768 272866 342088 272898
rect 372488 273454 372808 273486
rect 372488 273218 372530 273454
rect 372766 273218 372808 273454
rect 372488 273134 372808 273218
rect 372488 272898 372530 273134
rect 372766 272898 372808 273134
rect 372488 272866 372808 272898
rect 403208 273454 403528 273486
rect 403208 273218 403250 273454
rect 403486 273218 403528 273454
rect 403208 273134 403528 273218
rect 403208 272898 403250 273134
rect 403486 272898 403528 273134
rect 403208 272866 403528 272898
rect 433928 273454 434248 273486
rect 433928 273218 433970 273454
rect 434206 273218 434248 273454
rect 433928 273134 434248 273218
rect 433928 272898 433970 273134
rect 434206 272898 434248 273134
rect 433928 272866 434248 272898
rect 464648 273454 464968 273486
rect 464648 273218 464690 273454
rect 464926 273218 464968 273454
rect 464648 273134 464968 273218
rect 464648 272898 464690 273134
rect 464926 272898 464968 273134
rect 464648 272866 464968 272898
rect 495368 273454 495688 273486
rect 495368 273218 495410 273454
rect 495646 273218 495688 273454
rect 495368 273134 495688 273218
rect 495368 272898 495410 273134
rect 495646 272898 495688 273134
rect 495368 272866 495688 272898
rect 526088 273454 526408 273486
rect 526088 273218 526130 273454
rect 526366 273218 526408 273454
rect 526088 273134 526408 273218
rect 526088 272898 526130 273134
rect 526366 272898 526408 273134
rect 526088 272866 526408 272898
rect 19208 255454 19528 255486
rect 19208 255218 19250 255454
rect 19486 255218 19528 255454
rect 19208 255134 19528 255218
rect 19208 254898 19250 255134
rect 19486 254898 19528 255134
rect 19208 254866 19528 254898
rect 49928 255454 50248 255486
rect 49928 255218 49970 255454
rect 50206 255218 50248 255454
rect 49928 255134 50248 255218
rect 49928 254898 49970 255134
rect 50206 254898 50248 255134
rect 49928 254866 50248 254898
rect 80648 255454 80968 255486
rect 80648 255218 80690 255454
rect 80926 255218 80968 255454
rect 80648 255134 80968 255218
rect 80648 254898 80690 255134
rect 80926 254898 80968 255134
rect 80648 254866 80968 254898
rect 111368 255454 111688 255486
rect 111368 255218 111410 255454
rect 111646 255218 111688 255454
rect 111368 255134 111688 255218
rect 111368 254898 111410 255134
rect 111646 254898 111688 255134
rect 111368 254866 111688 254898
rect 142088 255454 142408 255486
rect 142088 255218 142130 255454
rect 142366 255218 142408 255454
rect 142088 255134 142408 255218
rect 142088 254898 142130 255134
rect 142366 254898 142408 255134
rect 142088 254866 142408 254898
rect 172808 255454 173128 255486
rect 172808 255218 172850 255454
rect 173086 255218 173128 255454
rect 172808 255134 173128 255218
rect 172808 254898 172850 255134
rect 173086 254898 173128 255134
rect 172808 254866 173128 254898
rect 203528 255454 203848 255486
rect 203528 255218 203570 255454
rect 203806 255218 203848 255454
rect 203528 255134 203848 255218
rect 203528 254898 203570 255134
rect 203806 254898 203848 255134
rect 203528 254866 203848 254898
rect 234248 255454 234568 255486
rect 234248 255218 234290 255454
rect 234526 255218 234568 255454
rect 234248 255134 234568 255218
rect 234248 254898 234290 255134
rect 234526 254898 234568 255134
rect 234248 254866 234568 254898
rect 264968 255454 265288 255486
rect 264968 255218 265010 255454
rect 265246 255218 265288 255454
rect 264968 255134 265288 255218
rect 264968 254898 265010 255134
rect 265246 254898 265288 255134
rect 264968 254866 265288 254898
rect 295688 255454 296008 255486
rect 295688 255218 295730 255454
rect 295966 255218 296008 255454
rect 295688 255134 296008 255218
rect 295688 254898 295730 255134
rect 295966 254898 296008 255134
rect 295688 254866 296008 254898
rect 326408 255454 326728 255486
rect 326408 255218 326450 255454
rect 326686 255218 326728 255454
rect 326408 255134 326728 255218
rect 326408 254898 326450 255134
rect 326686 254898 326728 255134
rect 326408 254866 326728 254898
rect 357128 255454 357448 255486
rect 357128 255218 357170 255454
rect 357406 255218 357448 255454
rect 357128 255134 357448 255218
rect 357128 254898 357170 255134
rect 357406 254898 357448 255134
rect 357128 254866 357448 254898
rect 387848 255454 388168 255486
rect 387848 255218 387890 255454
rect 388126 255218 388168 255454
rect 387848 255134 388168 255218
rect 387848 254898 387890 255134
rect 388126 254898 388168 255134
rect 387848 254866 388168 254898
rect 418568 255454 418888 255486
rect 418568 255218 418610 255454
rect 418846 255218 418888 255454
rect 418568 255134 418888 255218
rect 418568 254898 418610 255134
rect 418846 254898 418888 255134
rect 418568 254866 418888 254898
rect 449288 255454 449608 255486
rect 449288 255218 449330 255454
rect 449566 255218 449608 255454
rect 449288 255134 449608 255218
rect 449288 254898 449330 255134
rect 449566 254898 449608 255134
rect 449288 254866 449608 254898
rect 480008 255454 480328 255486
rect 480008 255218 480050 255454
rect 480286 255218 480328 255454
rect 480008 255134 480328 255218
rect 480008 254898 480050 255134
rect 480286 254898 480328 255134
rect 480008 254866 480328 254898
rect 510728 255454 511048 255486
rect 510728 255218 510770 255454
rect 511006 255218 511048 255454
rect 510728 255134 511048 255218
rect 510728 254898 510770 255134
rect 511006 254898 511048 255134
rect 510728 254866 511048 254898
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 34568 237454 34888 237486
rect 34568 237218 34610 237454
rect 34846 237218 34888 237454
rect 34568 237134 34888 237218
rect 34568 236898 34610 237134
rect 34846 236898 34888 237134
rect 34568 236866 34888 236898
rect 65288 237454 65608 237486
rect 65288 237218 65330 237454
rect 65566 237218 65608 237454
rect 65288 237134 65608 237218
rect 65288 236898 65330 237134
rect 65566 236898 65608 237134
rect 65288 236866 65608 236898
rect 96008 237454 96328 237486
rect 96008 237218 96050 237454
rect 96286 237218 96328 237454
rect 96008 237134 96328 237218
rect 96008 236898 96050 237134
rect 96286 236898 96328 237134
rect 96008 236866 96328 236898
rect 126728 237454 127048 237486
rect 126728 237218 126770 237454
rect 127006 237218 127048 237454
rect 126728 237134 127048 237218
rect 126728 236898 126770 237134
rect 127006 236898 127048 237134
rect 126728 236866 127048 236898
rect 157448 237454 157768 237486
rect 157448 237218 157490 237454
rect 157726 237218 157768 237454
rect 157448 237134 157768 237218
rect 157448 236898 157490 237134
rect 157726 236898 157768 237134
rect 157448 236866 157768 236898
rect 188168 237454 188488 237486
rect 188168 237218 188210 237454
rect 188446 237218 188488 237454
rect 188168 237134 188488 237218
rect 188168 236898 188210 237134
rect 188446 236898 188488 237134
rect 188168 236866 188488 236898
rect 218888 237454 219208 237486
rect 218888 237218 218930 237454
rect 219166 237218 219208 237454
rect 218888 237134 219208 237218
rect 218888 236898 218930 237134
rect 219166 236898 219208 237134
rect 218888 236866 219208 236898
rect 249608 237454 249928 237486
rect 249608 237218 249650 237454
rect 249886 237218 249928 237454
rect 249608 237134 249928 237218
rect 249608 236898 249650 237134
rect 249886 236898 249928 237134
rect 249608 236866 249928 236898
rect 280328 237454 280648 237486
rect 280328 237218 280370 237454
rect 280606 237218 280648 237454
rect 280328 237134 280648 237218
rect 280328 236898 280370 237134
rect 280606 236898 280648 237134
rect 280328 236866 280648 236898
rect 311048 237454 311368 237486
rect 311048 237218 311090 237454
rect 311326 237218 311368 237454
rect 311048 237134 311368 237218
rect 311048 236898 311090 237134
rect 311326 236898 311368 237134
rect 311048 236866 311368 236898
rect 341768 237454 342088 237486
rect 341768 237218 341810 237454
rect 342046 237218 342088 237454
rect 341768 237134 342088 237218
rect 341768 236898 341810 237134
rect 342046 236898 342088 237134
rect 341768 236866 342088 236898
rect 372488 237454 372808 237486
rect 372488 237218 372530 237454
rect 372766 237218 372808 237454
rect 372488 237134 372808 237218
rect 372488 236898 372530 237134
rect 372766 236898 372808 237134
rect 372488 236866 372808 236898
rect 403208 237454 403528 237486
rect 403208 237218 403250 237454
rect 403486 237218 403528 237454
rect 403208 237134 403528 237218
rect 403208 236898 403250 237134
rect 403486 236898 403528 237134
rect 403208 236866 403528 236898
rect 433928 237454 434248 237486
rect 433928 237218 433970 237454
rect 434206 237218 434248 237454
rect 433928 237134 434248 237218
rect 433928 236898 433970 237134
rect 434206 236898 434248 237134
rect 433928 236866 434248 236898
rect 464648 237454 464968 237486
rect 464648 237218 464690 237454
rect 464926 237218 464968 237454
rect 464648 237134 464968 237218
rect 464648 236898 464690 237134
rect 464926 236898 464968 237134
rect 464648 236866 464968 236898
rect 495368 237454 495688 237486
rect 495368 237218 495410 237454
rect 495646 237218 495688 237454
rect 495368 237134 495688 237218
rect 495368 236898 495410 237134
rect 495646 236898 495688 237134
rect 495368 236866 495688 236898
rect 526088 237454 526408 237486
rect 526088 237218 526130 237454
rect 526366 237218 526408 237454
rect 526088 237134 526408 237218
rect 526088 236898 526130 237134
rect 526366 236898 526408 237134
rect 526088 236866 526408 236898
rect 19208 219454 19528 219486
rect 19208 219218 19250 219454
rect 19486 219218 19528 219454
rect 19208 219134 19528 219218
rect 19208 218898 19250 219134
rect 19486 218898 19528 219134
rect 19208 218866 19528 218898
rect 49928 219454 50248 219486
rect 49928 219218 49970 219454
rect 50206 219218 50248 219454
rect 49928 219134 50248 219218
rect 49928 218898 49970 219134
rect 50206 218898 50248 219134
rect 49928 218866 50248 218898
rect 80648 219454 80968 219486
rect 80648 219218 80690 219454
rect 80926 219218 80968 219454
rect 80648 219134 80968 219218
rect 80648 218898 80690 219134
rect 80926 218898 80968 219134
rect 80648 218866 80968 218898
rect 111368 219454 111688 219486
rect 111368 219218 111410 219454
rect 111646 219218 111688 219454
rect 111368 219134 111688 219218
rect 111368 218898 111410 219134
rect 111646 218898 111688 219134
rect 111368 218866 111688 218898
rect 142088 219454 142408 219486
rect 142088 219218 142130 219454
rect 142366 219218 142408 219454
rect 142088 219134 142408 219218
rect 142088 218898 142130 219134
rect 142366 218898 142408 219134
rect 142088 218866 142408 218898
rect 172808 219454 173128 219486
rect 172808 219218 172850 219454
rect 173086 219218 173128 219454
rect 172808 219134 173128 219218
rect 172808 218898 172850 219134
rect 173086 218898 173128 219134
rect 172808 218866 173128 218898
rect 203528 219454 203848 219486
rect 203528 219218 203570 219454
rect 203806 219218 203848 219454
rect 203528 219134 203848 219218
rect 203528 218898 203570 219134
rect 203806 218898 203848 219134
rect 203528 218866 203848 218898
rect 234248 219454 234568 219486
rect 234248 219218 234290 219454
rect 234526 219218 234568 219454
rect 234248 219134 234568 219218
rect 234248 218898 234290 219134
rect 234526 218898 234568 219134
rect 234248 218866 234568 218898
rect 264968 219454 265288 219486
rect 264968 219218 265010 219454
rect 265246 219218 265288 219454
rect 264968 219134 265288 219218
rect 264968 218898 265010 219134
rect 265246 218898 265288 219134
rect 264968 218866 265288 218898
rect 295688 219454 296008 219486
rect 295688 219218 295730 219454
rect 295966 219218 296008 219454
rect 295688 219134 296008 219218
rect 295688 218898 295730 219134
rect 295966 218898 296008 219134
rect 295688 218866 296008 218898
rect 326408 219454 326728 219486
rect 326408 219218 326450 219454
rect 326686 219218 326728 219454
rect 326408 219134 326728 219218
rect 326408 218898 326450 219134
rect 326686 218898 326728 219134
rect 326408 218866 326728 218898
rect 357128 219454 357448 219486
rect 357128 219218 357170 219454
rect 357406 219218 357448 219454
rect 357128 219134 357448 219218
rect 357128 218898 357170 219134
rect 357406 218898 357448 219134
rect 357128 218866 357448 218898
rect 387848 219454 388168 219486
rect 387848 219218 387890 219454
rect 388126 219218 388168 219454
rect 387848 219134 388168 219218
rect 387848 218898 387890 219134
rect 388126 218898 388168 219134
rect 387848 218866 388168 218898
rect 418568 219454 418888 219486
rect 418568 219218 418610 219454
rect 418846 219218 418888 219454
rect 418568 219134 418888 219218
rect 418568 218898 418610 219134
rect 418846 218898 418888 219134
rect 418568 218866 418888 218898
rect 449288 219454 449608 219486
rect 449288 219218 449330 219454
rect 449566 219218 449608 219454
rect 449288 219134 449608 219218
rect 449288 218898 449330 219134
rect 449566 218898 449608 219134
rect 449288 218866 449608 218898
rect 480008 219454 480328 219486
rect 480008 219218 480050 219454
rect 480286 219218 480328 219454
rect 480008 219134 480328 219218
rect 480008 218898 480050 219134
rect 480286 218898 480328 219134
rect 480008 218866 480328 218898
rect 510728 219454 511048 219486
rect 510728 219218 510770 219454
rect 511006 219218 511048 219454
rect 510728 219134 511048 219218
rect 510728 218898 510770 219134
rect 511006 218898 511048 219134
rect 510728 218866 511048 218898
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 13675 208180 13741 208181
rect 13675 208116 13676 208180
rect 13740 208116 13741 208180
rect 13675 208115 13741 208116
rect 34568 201454 34888 201486
rect 34568 201218 34610 201454
rect 34846 201218 34888 201454
rect 34568 201134 34888 201218
rect 34568 200898 34610 201134
rect 34846 200898 34888 201134
rect 34568 200866 34888 200898
rect 65288 201454 65608 201486
rect 65288 201218 65330 201454
rect 65566 201218 65608 201454
rect 65288 201134 65608 201218
rect 65288 200898 65330 201134
rect 65566 200898 65608 201134
rect 65288 200866 65608 200898
rect 96008 201454 96328 201486
rect 96008 201218 96050 201454
rect 96286 201218 96328 201454
rect 96008 201134 96328 201218
rect 96008 200898 96050 201134
rect 96286 200898 96328 201134
rect 96008 200866 96328 200898
rect 126728 201454 127048 201486
rect 126728 201218 126770 201454
rect 127006 201218 127048 201454
rect 126728 201134 127048 201218
rect 126728 200898 126770 201134
rect 127006 200898 127048 201134
rect 126728 200866 127048 200898
rect 157448 201454 157768 201486
rect 157448 201218 157490 201454
rect 157726 201218 157768 201454
rect 157448 201134 157768 201218
rect 157448 200898 157490 201134
rect 157726 200898 157768 201134
rect 157448 200866 157768 200898
rect 188168 201454 188488 201486
rect 188168 201218 188210 201454
rect 188446 201218 188488 201454
rect 188168 201134 188488 201218
rect 188168 200898 188210 201134
rect 188446 200898 188488 201134
rect 188168 200866 188488 200898
rect 218888 201454 219208 201486
rect 218888 201218 218930 201454
rect 219166 201218 219208 201454
rect 218888 201134 219208 201218
rect 218888 200898 218930 201134
rect 219166 200898 219208 201134
rect 218888 200866 219208 200898
rect 249608 201454 249928 201486
rect 249608 201218 249650 201454
rect 249886 201218 249928 201454
rect 249608 201134 249928 201218
rect 249608 200898 249650 201134
rect 249886 200898 249928 201134
rect 249608 200866 249928 200898
rect 280328 201454 280648 201486
rect 280328 201218 280370 201454
rect 280606 201218 280648 201454
rect 280328 201134 280648 201218
rect 280328 200898 280370 201134
rect 280606 200898 280648 201134
rect 280328 200866 280648 200898
rect 311048 201454 311368 201486
rect 311048 201218 311090 201454
rect 311326 201218 311368 201454
rect 311048 201134 311368 201218
rect 311048 200898 311090 201134
rect 311326 200898 311368 201134
rect 311048 200866 311368 200898
rect 341768 201454 342088 201486
rect 341768 201218 341810 201454
rect 342046 201218 342088 201454
rect 341768 201134 342088 201218
rect 341768 200898 341810 201134
rect 342046 200898 342088 201134
rect 341768 200866 342088 200898
rect 372488 201454 372808 201486
rect 372488 201218 372530 201454
rect 372766 201218 372808 201454
rect 372488 201134 372808 201218
rect 372488 200898 372530 201134
rect 372766 200898 372808 201134
rect 372488 200866 372808 200898
rect 403208 201454 403528 201486
rect 403208 201218 403250 201454
rect 403486 201218 403528 201454
rect 403208 201134 403528 201218
rect 403208 200898 403250 201134
rect 403486 200898 403528 201134
rect 403208 200866 403528 200898
rect 433928 201454 434248 201486
rect 433928 201218 433970 201454
rect 434206 201218 434248 201454
rect 433928 201134 434248 201218
rect 433928 200898 433970 201134
rect 434206 200898 434248 201134
rect 433928 200866 434248 200898
rect 464648 201454 464968 201486
rect 464648 201218 464690 201454
rect 464926 201218 464968 201454
rect 464648 201134 464968 201218
rect 464648 200898 464690 201134
rect 464926 200898 464968 201134
rect 464648 200866 464968 200898
rect 495368 201454 495688 201486
rect 495368 201218 495410 201454
rect 495646 201218 495688 201454
rect 495368 201134 495688 201218
rect 495368 200898 495410 201134
rect 495646 200898 495688 201134
rect 495368 200866 495688 200898
rect 526088 201454 526408 201486
rect 526088 201218 526130 201454
rect 526366 201218 526408 201454
rect 526088 201134 526408 201218
rect 526088 200898 526130 201134
rect 526366 200898 526408 201134
rect 526088 200866 526408 200898
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 19208 183454 19528 183486
rect 19208 183218 19250 183454
rect 19486 183218 19528 183454
rect 19208 183134 19528 183218
rect 19208 182898 19250 183134
rect 19486 182898 19528 183134
rect 19208 182866 19528 182898
rect 49928 183454 50248 183486
rect 49928 183218 49970 183454
rect 50206 183218 50248 183454
rect 49928 183134 50248 183218
rect 49928 182898 49970 183134
rect 50206 182898 50248 183134
rect 49928 182866 50248 182898
rect 80648 183454 80968 183486
rect 80648 183218 80690 183454
rect 80926 183218 80968 183454
rect 80648 183134 80968 183218
rect 80648 182898 80690 183134
rect 80926 182898 80968 183134
rect 80648 182866 80968 182898
rect 111368 183454 111688 183486
rect 111368 183218 111410 183454
rect 111646 183218 111688 183454
rect 111368 183134 111688 183218
rect 111368 182898 111410 183134
rect 111646 182898 111688 183134
rect 111368 182866 111688 182898
rect 142088 183454 142408 183486
rect 142088 183218 142130 183454
rect 142366 183218 142408 183454
rect 142088 183134 142408 183218
rect 142088 182898 142130 183134
rect 142366 182898 142408 183134
rect 142088 182866 142408 182898
rect 172808 183454 173128 183486
rect 172808 183218 172850 183454
rect 173086 183218 173128 183454
rect 172808 183134 173128 183218
rect 172808 182898 172850 183134
rect 173086 182898 173128 183134
rect 172808 182866 173128 182898
rect 203528 183454 203848 183486
rect 203528 183218 203570 183454
rect 203806 183218 203848 183454
rect 203528 183134 203848 183218
rect 203528 182898 203570 183134
rect 203806 182898 203848 183134
rect 203528 182866 203848 182898
rect 234248 183454 234568 183486
rect 234248 183218 234290 183454
rect 234526 183218 234568 183454
rect 234248 183134 234568 183218
rect 234248 182898 234290 183134
rect 234526 182898 234568 183134
rect 234248 182866 234568 182898
rect 264968 183454 265288 183486
rect 264968 183218 265010 183454
rect 265246 183218 265288 183454
rect 264968 183134 265288 183218
rect 264968 182898 265010 183134
rect 265246 182898 265288 183134
rect 264968 182866 265288 182898
rect 295688 183454 296008 183486
rect 295688 183218 295730 183454
rect 295966 183218 296008 183454
rect 295688 183134 296008 183218
rect 295688 182898 295730 183134
rect 295966 182898 296008 183134
rect 295688 182866 296008 182898
rect 326408 183454 326728 183486
rect 326408 183218 326450 183454
rect 326686 183218 326728 183454
rect 326408 183134 326728 183218
rect 326408 182898 326450 183134
rect 326686 182898 326728 183134
rect 326408 182866 326728 182898
rect 357128 183454 357448 183486
rect 357128 183218 357170 183454
rect 357406 183218 357448 183454
rect 357128 183134 357448 183218
rect 357128 182898 357170 183134
rect 357406 182898 357448 183134
rect 357128 182866 357448 182898
rect 387848 183454 388168 183486
rect 387848 183218 387890 183454
rect 388126 183218 388168 183454
rect 387848 183134 388168 183218
rect 387848 182898 387890 183134
rect 388126 182898 388168 183134
rect 387848 182866 388168 182898
rect 418568 183454 418888 183486
rect 418568 183218 418610 183454
rect 418846 183218 418888 183454
rect 418568 183134 418888 183218
rect 418568 182898 418610 183134
rect 418846 182898 418888 183134
rect 418568 182866 418888 182898
rect 449288 183454 449608 183486
rect 449288 183218 449330 183454
rect 449566 183218 449608 183454
rect 449288 183134 449608 183218
rect 449288 182898 449330 183134
rect 449566 182898 449608 183134
rect 449288 182866 449608 182898
rect 480008 183454 480328 183486
rect 480008 183218 480050 183454
rect 480286 183218 480328 183454
rect 480008 183134 480328 183218
rect 480008 182898 480050 183134
rect 480286 182898 480328 183134
rect 480008 182866 480328 182898
rect 510728 183454 511048 183486
rect 510728 183218 510770 183454
rect 511006 183218 511048 183454
rect 510728 183134 511048 183218
rect 510728 182898 510770 183134
rect 511006 182898 511048 183134
rect 510728 182866 511048 182898
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 34568 165454 34888 165486
rect 34568 165218 34610 165454
rect 34846 165218 34888 165454
rect 34568 165134 34888 165218
rect 34568 164898 34610 165134
rect 34846 164898 34888 165134
rect 34568 164866 34888 164898
rect 65288 165454 65608 165486
rect 65288 165218 65330 165454
rect 65566 165218 65608 165454
rect 65288 165134 65608 165218
rect 65288 164898 65330 165134
rect 65566 164898 65608 165134
rect 65288 164866 65608 164898
rect 96008 165454 96328 165486
rect 96008 165218 96050 165454
rect 96286 165218 96328 165454
rect 96008 165134 96328 165218
rect 96008 164898 96050 165134
rect 96286 164898 96328 165134
rect 96008 164866 96328 164898
rect 126728 165454 127048 165486
rect 126728 165218 126770 165454
rect 127006 165218 127048 165454
rect 126728 165134 127048 165218
rect 126728 164898 126770 165134
rect 127006 164898 127048 165134
rect 126728 164866 127048 164898
rect 157448 165454 157768 165486
rect 157448 165218 157490 165454
rect 157726 165218 157768 165454
rect 157448 165134 157768 165218
rect 157448 164898 157490 165134
rect 157726 164898 157768 165134
rect 157448 164866 157768 164898
rect 188168 165454 188488 165486
rect 188168 165218 188210 165454
rect 188446 165218 188488 165454
rect 188168 165134 188488 165218
rect 188168 164898 188210 165134
rect 188446 164898 188488 165134
rect 188168 164866 188488 164898
rect 218888 165454 219208 165486
rect 218888 165218 218930 165454
rect 219166 165218 219208 165454
rect 218888 165134 219208 165218
rect 218888 164898 218930 165134
rect 219166 164898 219208 165134
rect 218888 164866 219208 164898
rect 249608 165454 249928 165486
rect 249608 165218 249650 165454
rect 249886 165218 249928 165454
rect 249608 165134 249928 165218
rect 249608 164898 249650 165134
rect 249886 164898 249928 165134
rect 249608 164866 249928 164898
rect 280328 165454 280648 165486
rect 280328 165218 280370 165454
rect 280606 165218 280648 165454
rect 280328 165134 280648 165218
rect 280328 164898 280370 165134
rect 280606 164898 280648 165134
rect 280328 164866 280648 164898
rect 311048 165454 311368 165486
rect 311048 165218 311090 165454
rect 311326 165218 311368 165454
rect 311048 165134 311368 165218
rect 311048 164898 311090 165134
rect 311326 164898 311368 165134
rect 311048 164866 311368 164898
rect 341768 165454 342088 165486
rect 341768 165218 341810 165454
rect 342046 165218 342088 165454
rect 341768 165134 342088 165218
rect 341768 164898 341810 165134
rect 342046 164898 342088 165134
rect 341768 164866 342088 164898
rect 372488 165454 372808 165486
rect 372488 165218 372530 165454
rect 372766 165218 372808 165454
rect 372488 165134 372808 165218
rect 372488 164898 372530 165134
rect 372766 164898 372808 165134
rect 372488 164866 372808 164898
rect 403208 165454 403528 165486
rect 403208 165218 403250 165454
rect 403486 165218 403528 165454
rect 403208 165134 403528 165218
rect 403208 164898 403250 165134
rect 403486 164898 403528 165134
rect 403208 164866 403528 164898
rect 433928 165454 434248 165486
rect 433928 165218 433970 165454
rect 434206 165218 434248 165454
rect 433928 165134 434248 165218
rect 433928 164898 433970 165134
rect 434206 164898 434248 165134
rect 433928 164866 434248 164898
rect 464648 165454 464968 165486
rect 464648 165218 464690 165454
rect 464926 165218 464968 165454
rect 464648 165134 464968 165218
rect 464648 164898 464690 165134
rect 464926 164898 464968 165134
rect 464648 164866 464968 164898
rect 495368 165454 495688 165486
rect 495368 165218 495410 165454
rect 495646 165218 495688 165454
rect 495368 165134 495688 165218
rect 495368 164898 495410 165134
rect 495646 164898 495688 165134
rect 495368 164866 495688 164898
rect 526088 165454 526408 165486
rect 526088 165218 526130 165454
rect 526366 165218 526408 165454
rect 526088 165134 526408 165218
rect 526088 164898 526130 165134
rect 526366 164898 526408 165134
rect 526088 164866 526408 164898
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 19208 147454 19528 147486
rect 19208 147218 19250 147454
rect 19486 147218 19528 147454
rect 19208 147134 19528 147218
rect 19208 146898 19250 147134
rect 19486 146898 19528 147134
rect 19208 146866 19528 146898
rect 49928 147454 50248 147486
rect 49928 147218 49970 147454
rect 50206 147218 50248 147454
rect 49928 147134 50248 147218
rect 49928 146898 49970 147134
rect 50206 146898 50248 147134
rect 49928 146866 50248 146898
rect 80648 147454 80968 147486
rect 80648 147218 80690 147454
rect 80926 147218 80968 147454
rect 80648 147134 80968 147218
rect 80648 146898 80690 147134
rect 80926 146898 80968 147134
rect 80648 146866 80968 146898
rect 111368 147454 111688 147486
rect 111368 147218 111410 147454
rect 111646 147218 111688 147454
rect 111368 147134 111688 147218
rect 111368 146898 111410 147134
rect 111646 146898 111688 147134
rect 111368 146866 111688 146898
rect 142088 147454 142408 147486
rect 142088 147218 142130 147454
rect 142366 147218 142408 147454
rect 142088 147134 142408 147218
rect 142088 146898 142130 147134
rect 142366 146898 142408 147134
rect 142088 146866 142408 146898
rect 172808 147454 173128 147486
rect 172808 147218 172850 147454
rect 173086 147218 173128 147454
rect 172808 147134 173128 147218
rect 172808 146898 172850 147134
rect 173086 146898 173128 147134
rect 172808 146866 173128 146898
rect 203528 147454 203848 147486
rect 203528 147218 203570 147454
rect 203806 147218 203848 147454
rect 203528 147134 203848 147218
rect 203528 146898 203570 147134
rect 203806 146898 203848 147134
rect 203528 146866 203848 146898
rect 234248 147454 234568 147486
rect 234248 147218 234290 147454
rect 234526 147218 234568 147454
rect 234248 147134 234568 147218
rect 234248 146898 234290 147134
rect 234526 146898 234568 147134
rect 234248 146866 234568 146898
rect 264968 147454 265288 147486
rect 264968 147218 265010 147454
rect 265246 147218 265288 147454
rect 264968 147134 265288 147218
rect 264968 146898 265010 147134
rect 265246 146898 265288 147134
rect 264968 146866 265288 146898
rect 295688 147454 296008 147486
rect 295688 147218 295730 147454
rect 295966 147218 296008 147454
rect 295688 147134 296008 147218
rect 295688 146898 295730 147134
rect 295966 146898 296008 147134
rect 295688 146866 296008 146898
rect 326408 147454 326728 147486
rect 326408 147218 326450 147454
rect 326686 147218 326728 147454
rect 326408 147134 326728 147218
rect 326408 146898 326450 147134
rect 326686 146898 326728 147134
rect 326408 146866 326728 146898
rect 357128 147454 357448 147486
rect 357128 147218 357170 147454
rect 357406 147218 357448 147454
rect 357128 147134 357448 147218
rect 357128 146898 357170 147134
rect 357406 146898 357448 147134
rect 357128 146866 357448 146898
rect 387848 147454 388168 147486
rect 387848 147218 387890 147454
rect 388126 147218 388168 147454
rect 387848 147134 388168 147218
rect 387848 146898 387890 147134
rect 388126 146898 388168 147134
rect 387848 146866 388168 146898
rect 418568 147454 418888 147486
rect 418568 147218 418610 147454
rect 418846 147218 418888 147454
rect 418568 147134 418888 147218
rect 418568 146898 418610 147134
rect 418846 146898 418888 147134
rect 418568 146866 418888 146898
rect 449288 147454 449608 147486
rect 449288 147218 449330 147454
rect 449566 147218 449608 147454
rect 449288 147134 449608 147218
rect 449288 146898 449330 147134
rect 449566 146898 449608 147134
rect 449288 146866 449608 146898
rect 480008 147454 480328 147486
rect 480008 147218 480050 147454
rect 480286 147218 480328 147454
rect 480008 147134 480328 147218
rect 480008 146898 480050 147134
rect 480286 146898 480328 147134
rect 480008 146866 480328 146898
rect 510728 147454 511048 147486
rect 510728 147218 510770 147454
rect 511006 147218 511048 147454
rect 510728 147134 511048 147218
rect 510728 146898 510770 147134
rect 511006 146898 511048 147134
rect 510728 146866 511048 146898
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 34568 129454 34888 129486
rect 34568 129218 34610 129454
rect 34846 129218 34888 129454
rect 34568 129134 34888 129218
rect 34568 128898 34610 129134
rect 34846 128898 34888 129134
rect 34568 128866 34888 128898
rect 65288 129454 65608 129486
rect 65288 129218 65330 129454
rect 65566 129218 65608 129454
rect 65288 129134 65608 129218
rect 65288 128898 65330 129134
rect 65566 128898 65608 129134
rect 65288 128866 65608 128898
rect 96008 129454 96328 129486
rect 96008 129218 96050 129454
rect 96286 129218 96328 129454
rect 96008 129134 96328 129218
rect 96008 128898 96050 129134
rect 96286 128898 96328 129134
rect 96008 128866 96328 128898
rect 126728 129454 127048 129486
rect 126728 129218 126770 129454
rect 127006 129218 127048 129454
rect 126728 129134 127048 129218
rect 126728 128898 126770 129134
rect 127006 128898 127048 129134
rect 126728 128866 127048 128898
rect 157448 129454 157768 129486
rect 157448 129218 157490 129454
rect 157726 129218 157768 129454
rect 157448 129134 157768 129218
rect 157448 128898 157490 129134
rect 157726 128898 157768 129134
rect 157448 128866 157768 128898
rect 188168 129454 188488 129486
rect 188168 129218 188210 129454
rect 188446 129218 188488 129454
rect 188168 129134 188488 129218
rect 188168 128898 188210 129134
rect 188446 128898 188488 129134
rect 188168 128866 188488 128898
rect 218888 129454 219208 129486
rect 218888 129218 218930 129454
rect 219166 129218 219208 129454
rect 218888 129134 219208 129218
rect 218888 128898 218930 129134
rect 219166 128898 219208 129134
rect 218888 128866 219208 128898
rect 249608 129454 249928 129486
rect 249608 129218 249650 129454
rect 249886 129218 249928 129454
rect 249608 129134 249928 129218
rect 249608 128898 249650 129134
rect 249886 128898 249928 129134
rect 249608 128866 249928 128898
rect 280328 129454 280648 129486
rect 280328 129218 280370 129454
rect 280606 129218 280648 129454
rect 280328 129134 280648 129218
rect 280328 128898 280370 129134
rect 280606 128898 280648 129134
rect 280328 128866 280648 128898
rect 311048 129454 311368 129486
rect 311048 129218 311090 129454
rect 311326 129218 311368 129454
rect 311048 129134 311368 129218
rect 311048 128898 311090 129134
rect 311326 128898 311368 129134
rect 311048 128866 311368 128898
rect 341768 129454 342088 129486
rect 341768 129218 341810 129454
rect 342046 129218 342088 129454
rect 341768 129134 342088 129218
rect 341768 128898 341810 129134
rect 342046 128898 342088 129134
rect 341768 128866 342088 128898
rect 372488 129454 372808 129486
rect 372488 129218 372530 129454
rect 372766 129218 372808 129454
rect 372488 129134 372808 129218
rect 372488 128898 372530 129134
rect 372766 128898 372808 129134
rect 372488 128866 372808 128898
rect 403208 129454 403528 129486
rect 403208 129218 403250 129454
rect 403486 129218 403528 129454
rect 403208 129134 403528 129218
rect 403208 128898 403250 129134
rect 403486 128898 403528 129134
rect 403208 128866 403528 128898
rect 433928 129454 434248 129486
rect 433928 129218 433970 129454
rect 434206 129218 434248 129454
rect 433928 129134 434248 129218
rect 433928 128898 433970 129134
rect 434206 128898 434248 129134
rect 433928 128866 434248 128898
rect 464648 129454 464968 129486
rect 464648 129218 464690 129454
rect 464926 129218 464968 129454
rect 464648 129134 464968 129218
rect 464648 128898 464690 129134
rect 464926 128898 464968 129134
rect 464648 128866 464968 128898
rect 495368 129454 495688 129486
rect 495368 129218 495410 129454
rect 495646 129218 495688 129454
rect 495368 129134 495688 129218
rect 495368 128898 495410 129134
rect 495646 128898 495688 129134
rect 495368 128866 495688 128898
rect 526088 129454 526408 129486
rect 526088 129218 526130 129454
rect 526366 129218 526408 129454
rect 526088 129134 526408 129218
rect 526088 128898 526130 129134
rect 526366 128898 526408 129134
rect 526088 128866 526408 128898
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 19208 111454 19528 111486
rect 19208 111218 19250 111454
rect 19486 111218 19528 111454
rect 19208 111134 19528 111218
rect 19208 110898 19250 111134
rect 19486 110898 19528 111134
rect 19208 110866 19528 110898
rect 49928 111454 50248 111486
rect 49928 111218 49970 111454
rect 50206 111218 50248 111454
rect 49928 111134 50248 111218
rect 49928 110898 49970 111134
rect 50206 110898 50248 111134
rect 49928 110866 50248 110898
rect 80648 111454 80968 111486
rect 80648 111218 80690 111454
rect 80926 111218 80968 111454
rect 80648 111134 80968 111218
rect 80648 110898 80690 111134
rect 80926 110898 80968 111134
rect 80648 110866 80968 110898
rect 111368 111454 111688 111486
rect 111368 111218 111410 111454
rect 111646 111218 111688 111454
rect 111368 111134 111688 111218
rect 111368 110898 111410 111134
rect 111646 110898 111688 111134
rect 111368 110866 111688 110898
rect 142088 111454 142408 111486
rect 142088 111218 142130 111454
rect 142366 111218 142408 111454
rect 142088 111134 142408 111218
rect 142088 110898 142130 111134
rect 142366 110898 142408 111134
rect 142088 110866 142408 110898
rect 172808 111454 173128 111486
rect 172808 111218 172850 111454
rect 173086 111218 173128 111454
rect 172808 111134 173128 111218
rect 172808 110898 172850 111134
rect 173086 110898 173128 111134
rect 172808 110866 173128 110898
rect 203528 111454 203848 111486
rect 203528 111218 203570 111454
rect 203806 111218 203848 111454
rect 203528 111134 203848 111218
rect 203528 110898 203570 111134
rect 203806 110898 203848 111134
rect 203528 110866 203848 110898
rect 234248 111454 234568 111486
rect 234248 111218 234290 111454
rect 234526 111218 234568 111454
rect 234248 111134 234568 111218
rect 234248 110898 234290 111134
rect 234526 110898 234568 111134
rect 234248 110866 234568 110898
rect 264968 111454 265288 111486
rect 264968 111218 265010 111454
rect 265246 111218 265288 111454
rect 264968 111134 265288 111218
rect 264968 110898 265010 111134
rect 265246 110898 265288 111134
rect 264968 110866 265288 110898
rect 295688 111454 296008 111486
rect 295688 111218 295730 111454
rect 295966 111218 296008 111454
rect 295688 111134 296008 111218
rect 295688 110898 295730 111134
rect 295966 110898 296008 111134
rect 295688 110866 296008 110898
rect 326408 111454 326728 111486
rect 326408 111218 326450 111454
rect 326686 111218 326728 111454
rect 326408 111134 326728 111218
rect 326408 110898 326450 111134
rect 326686 110898 326728 111134
rect 326408 110866 326728 110898
rect 357128 111454 357448 111486
rect 357128 111218 357170 111454
rect 357406 111218 357448 111454
rect 357128 111134 357448 111218
rect 357128 110898 357170 111134
rect 357406 110898 357448 111134
rect 357128 110866 357448 110898
rect 387848 111454 388168 111486
rect 387848 111218 387890 111454
rect 388126 111218 388168 111454
rect 387848 111134 388168 111218
rect 387848 110898 387890 111134
rect 388126 110898 388168 111134
rect 387848 110866 388168 110898
rect 418568 111454 418888 111486
rect 418568 111218 418610 111454
rect 418846 111218 418888 111454
rect 418568 111134 418888 111218
rect 418568 110898 418610 111134
rect 418846 110898 418888 111134
rect 418568 110866 418888 110898
rect 449288 111454 449608 111486
rect 449288 111218 449330 111454
rect 449566 111218 449608 111454
rect 449288 111134 449608 111218
rect 449288 110898 449330 111134
rect 449566 110898 449608 111134
rect 449288 110866 449608 110898
rect 480008 111454 480328 111486
rect 480008 111218 480050 111454
rect 480286 111218 480328 111454
rect 480008 111134 480328 111218
rect 480008 110898 480050 111134
rect 480286 110898 480328 111134
rect 480008 110866 480328 110898
rect 510728 111454 511048 111486
rect 510728 111218 510770 111454
rect 511006 111218 511048 111454
rect 510728 111134 511048 111218
rect 510728 110898 510770 111134
rect 511006 110898 511048 111134
rect 510728 110866 511048 110898
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 34568 93454 34888 93486
rect 34568 93218 34610 93454
rect 34846 93218 34888 93454
rect 34568 93134 34888 93218
rect 34568 92898 34610 93134
rect 34846 92898 34888 93134
rect 34568 92866 34888 92898
rect 65288 93454 65608 93486
rect 65288 93218 65330 93454
rect 65566 93218 65608 93454
rect 65288 93134 65608 93218
rect 65288 92898 65330 93134
rect 65566 92898 65608 93134
rect 65288 92866 65608 92898
rect 96008 93454 96328 93486
rect 96008 93218 96050 93454
rect 96286 93218 96328 93454
rect 96008 93134 96328 93218
rect 96008 92898 96050 93134
rect 96286 92898 96328 93134
rect 96008 92866 96328 92898
rect 126728 93454 127048 93486
rect 126728 93218 126770 93454
rect 127006 93218 127048 93454
rect 126728 93134 127048 93218
rect 126728 92898 126770 93134
rect 127006 92898 127048 93134
rect 126728 92866 127048 92898
rect 157448 93454 157768 93486
rect 157448 93218 157490 93454
rect 157726 93218 157768 93454
rect 157448 93134 157768 93218
rect 157448 92898 157490 93134
rect 157726 92898 157768 93134
rect 157448 92866 157768 92898
rect 188168 93454 188488 93486
rect 188168 93218 188210 93454
rect 188446 93218 188488 93454
rect 188168 93134 188488 93218
rect 188168 92898 188210 93134
rect 188446 92898 188488 93134
rect 188168 92866 188488 92898
rect 218888 93454 219208 93486
rect 218888 93218 218930 93454
rect 219166 93218 219208 93454
rect 218888 93134 219208 93218
rect 218888 92898 218930 93134
rect 219166 92898 219208 93134
rect 218888 92866 219208 92898
rect 249608 93454 249928 93486
rect 249608 93218 249650 93454
rect 249886 93218 249928 93454
rect 249608 93134 249928 93218
rect 249608 92898 249650 93134
rect 249886 92898 249928 93134
rect 249608 92866 249928 92898
rect 280328 93454 280648 93486
rect 280328 93218 280370 93454
rect 280606 93218 280648 93454
rect 280328 93134 280648 93218
rect 280328 92898 280370 93134
rect 280606 92898 280648 93134
rect 280328 92866 280648 92898
rect 311048 93454 311368 93486
rect 311048 93218 311090 93454
rect 311326 93218 311368 93454
rect 311048 93134 311368 93218
rect 311048 92898 311090 93134
rect 311326 92898 311368 93134
rect 311048 92866 311368 92898
rect 341768 93454 342088 93486
rect 341768 93218 341810 93454
rect 342046 93218 342088 93454
rect 341768 93134 342088 93218
rect 341768 92898 341810 93134
rect 342046 92898 342088 93134
rect 341768 92866 342088 92898
rect 372488 93454 372808 93486
rect 372488 93218 372530 93454
rect 372766 93218 372808 93454
rect 372488 93134 372808 93218
rect 372488 92898 372530 93134
rect 372766 92898 372808 93134
rect 372488 92866 372808 92898
rect 403208 93454 403528 93486
rect 403208 93218 403250 93454
rect 403486 93218 403528 93454
rect 403208 93134 403528 93218
rect 403208 92898 403250 93134
rect 403486 92898 403528 93134
rect 403208 92866 403528 92898
rect 433928 93454 434248 93486
rect 433928 93218 433970 93454
rect 434206 93218 434248 93454
rect 433928 93134 434248 93218
rect 433928 92898 433970 93134
rect 434206 92898 434248 93134
rect 433928 92866 434248 92898
rect 464648 93454 464968 93486
rect 464648 93218 464690 93454
rect 464926 93218 464968 93454
rect 464648 93134 464968 93218
rect 464648 92898 464690 93134
rect 464926 92898 464968 93134
rect 464648 92866 464968 92898
rect 495368 93454 495688 93486
rect 495368 93218 495410 93454
rect 495646 93218 495688 93454
rect 495368 93134 495688 93218
rect 495368 92898 495410 93134
rect 495646 92898 495688 93134
rect 495368 92866 495688 92898
rect 526088 93454 526408 93486
rect 526088 93218 526130 93454
rect 526366 93218 526408 93454
rect 526088 93134 526408 93218
rect 526088 92898 526130 93134
rect 526366 92898 526408 93134
rect 526088 92866 526408 92898
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 19208 75454 19528 75486
rect 19208 75218 19250 75454
rect 19486 75218 19528 75454
rect 19208 75134 19528 75218
rect 19208 74898 19250 75134
rect 19486 74898 19528 75134
rect 19208 74866 19528 74898
rect 49928 75454 50248 75486
rect 49928 75218 49970 75454
rect 50206 75218 50248 75454
rect 49928 75134 50248 75218
rect 49928 74898 49970 75134
rect 50206 74898 50248 75134
rect 49928 74866 50248 74898
rect 80648 75454 80968 75486
rect 80648 75218 80690 75454
rect 80926 75218 80968 75454
rect 80648 75134 80968 75218
rect 80648 74898 80690 75134
rect 80926 74898 80968 75134
rect 80648 74866 80968 74898
rect 111368 75454 111688 75486
rect 111368 75218 111410 75454
rect 111646 75218 111688 75454
rect 111368 75134 111688 75218
rect 111368 74898 111410 75134
rect 111646 74898 111688 75134
rect 111368 74866 111688 74898
rect 142088 75454 142408 75486
rect 142088 75218 142130 75454
rect 142366 75218 142408 75454
rect 142088 75134 142408 75218
rect 142088 74898 142130 75134
rect 142366 74898 142408 75134
rect 142088 74866 142408 74898
rect 172808 75454 173128 75486
rect 172808 75218 172850 75454
rect 173086 75218 173128 75454
rect 172808 75134 173128 75218
rect 172808 74898 172850 75134
rect 173086 74898 173128 75134
rect 172808 74866 173128 74898
rect 203528 75454 203848 75486
rect 203528 75218 203570 75454
rect 203806 75218 203848 75454
rect 203528 75134 203848 75218
rect 203528 74898 203570 75134
rect 203806 74898 203848 75134
rect 203528 74866 203848 74898
rect 234248 75454 234568 75486
rect 234248 75218 234290 75454
rect 234526 75218 234568 75454
rect 234248 75134 234568 75218
rect 234248 74898 234290 75134
rect 234526 74898 234568 75134
rect 234248 74866 234568 74898
rect 264968 75454 265288 75486
rect 264968 75218 265010 75454
rect 265246 75218 265288 75454
rect 264968 75134 265288 75218
rect 264968 74898 265010 75134
rect 265246 74898 265288 75134
rect 264968 74866 265288 74898
rect 295688 75454 296008 75486
rect 295688 75218 295730 75454
rect 295966 75218 296008 75454
rect 295688 75134 296008 75218
rect 295688 74898 295730 75134
rect 295966 74898 296008 75134
rect 295688 74866 296008 74898
rect 326408 75454 326728 75486
rect 326408 75218 326450 75454
rect 326686 75218 326728 75454
rect 326408 75134 326728 75218
rect 326408 74898 326450 75134
rect 326686 74898 326728 75134
rect 326408 74866 326728 74898
rect 357128 75454 357448 75486
rect 357128 75218 357170 75454
rect 357406 75218 357448 75454
rect 357128 75134 357448 75218
rect 357128 74898 357170 75134
rect 357406 74898 357448 75134
rect 357128 74866 357448 74898
rect 387848 75454 388168 75486
rect 387848 75218 387890 75454
rect 388126 75218 388168 75454
rect 387848 75134 388168 75218
rect 387848 74898 387890 75134
rect 388126 74898 388168 75134
rect 387848 74866 388168 74898
rect 418568 75454 418888 75486
rect 418568 75218 418610 75454
rect 418846 75218 418888 75454
rect 418568 75134 418888 75218
rect 418568 74898 418610 75134
rect 418846 74898 418888 75134
rect 418568 74866 418888 74898
rect 449288 75454 449608 75486
rect 449288 75218 449330 75454
rect 449566 75218 449608 75454
rect 449288 75134 449608 75218
rect 449288 74898 449330 75134
rect 449566 74898 449608 75134
rect 449288 74866 449608 74898
rect 480008 75454 480328 75486
rect 480008 75218 480050 75454
rect 480286 75218 480328 75454
rect 480008 75134 480328 75218
rect 480008 74898 480050 75134
rect 480286 74898 480328 75134
rect 480008 74866 480328 74898
rect 510728 75454 511048 75486
rect 510728 75218 510770 75454
rect 511006 75218 511048 75454
rect 510728 75134 511048 75218
rect 510728 74898 510770 75134
rect 511006 74898 511048 75134
rect 510728 74866 511048 74898
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 34568 57454 34888 57486
rect 34568 57218 34610 57454
rect 34846 57218 34888 57454
rect 34568 57134 34888 57218
rect 34568 56898 34610 57134
rect 34846 56898 34888 57134
rect 34568 56866 34888 56898
rect 65288 57454 65608 57486
rect 65288 57218 65330 57454
rect 65566 57218 65608 57454
rect 65288 57134 65608 57218
rect 65288 56898 65330 57134
rect 65566 56898 65608 57134
rect 65288 56866 65608 56898
rect 96008 57454 96328 57486
rect 96008 57218 96050 57454
rect 96286 57218 96328 57454
rect 96008 57134 96328 57218
rect 96008 56898 96050 57134
rect 96286 56898 96328 57134
rect 96008 56866 96328 56898
rect 126728 57454 127048 57486
rect 126728 57218 126770 57454
rect 127006 57218 127048 57454
rect 126728 57134 127048 57218
rect 126728 56898 126770 57134
rect 127006 56898 127048 57134
rect 126728 56866 127048 56898
rect 157448 57454 157768 57486
rect 157448 57218 157490 57454
rect 157726 57218 157768 57454
rect 157448 57134 157768 57218
rect 157448 56898 157490 57134
rect 157726 56898 157768 57134
rect 157448 56866 157768 56898
rect 188168 57454 188488 57486
rect 188168 57218 188210 57454
rect 188446 57218 188488 57454
rect 188168 57134 188488 57218
rect 188168 56898 188210 57134
rect 188446 56898 188488 57134
rect 188168 56866 188488 56898
rect 218888 57454 219208 57486
rect 218888 57218 218930 57454
rect 219166 57218 219208 57454
rect 218888 57134 219208 57218
rect 218888 56898 218930 57134
rect 219166 56898 219208 57134
rect 218888 56866 219208 56898
rect 249608 57454 249928 57486
rect 249608 57218 249650 57454
rect 249886 57218 249928 57454
rect 249608 57134 249928 57218
rect 249608 56898 249650 57134
rect 249886 56898 249928 57134
rect 249608 56866 249928 56898
rect 280328 57454 280648 57486
rect 280328 57218 280370 57454
rect 280606 57218 280648 57454
rect 280328 57134 280648 57218
rect 280328 56898 280370 57134
rect 280606 56898 280648 57134
rect 280328 56866 280648 56898
rect 311048 57454 311368 57486
rect 311048 57218 311090 57454
rect 311326 57218 311368 57454
rect 311048 57134 311368 57218
rect 311048 56898 311090 57134
rect 311326 56898 311368 57134
rect 311048 56866 311368 56898
rect 341768 57454 342088 57486
rect 341768 57218 341810 57454
rect 342046 57218 342088 57454
rect 341768 57134 342088 57218
rect 341768 56898 341810 57134
rect 342046 56898 342088 57134
rect 341768 56866 342088 56898
rect 372488 57454 372808 57486
rect 372488 57218 372530 57454
rect 372766 57218 372808 57454
rect 372488 57134 372808 57218
rect 372488 56898 372530 57134
rect 372766 56898 372808 57134
rect 372488 56866 372808 56898
rect 403208 57454 403528 57486
rect 403208 57218 403250 57454
rect 403486 57218 403528 57454
rect 403208 57134 403528 57218
rect 403208 56898 403250 57134
rect 403486 56898 403528 57134
rect 403208 56866 403528 56898
rect 433928 57454 434248 57486
rect 433928 57218 433970 57454
rect 434206 57218 434248 57454
rect 433928 57134 434248 57218
rect 433928 56898 433970 57134
rect 434206 56898 434248 57134
rect 433928 56866 434248 56898
rect 464648 57454 464968 57486
rect 464648 57218 464690 57454
rect 464926 57218 464968 57454
rect 464648 57134 464968 57218
rect 464648 56898 464690 57134
rect 464926 56898 464968 57134
rect 464648 56866 464968 56898
rect 495368 57454 495688 57486
rect 495368 57218 495410 57454
rect 495646 57218 495688 57454
rect 495368 57134 495688 57218
rect 495368 56898 495410 57134
rect 495646 56898 495688 57134
rect 495368 56866 495688 56898
rect 526088 57454 526408 57486
rect 526088 57218 526130 57454
rect 526366 57218 526408 57454
rect 526088 57134 526408 57218
rect 526088 56898 526130 57134
rect 526366 56898 526408 57134
rect 526088 56866 526408 56898
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 19208 39454 19528 39486
rect 19208 39218 19250 39454
rect 19486 39218 19528 39454
rect 19208 39134 19528 39218
rect 19208 38898 19250 39134
rect 19486 38898 19528 39134
rect 19208 38866 19528 38898
rect 49928 39454 50248 39486
rect 49928 39218 49970 39454
rect 50206 39218 50248 39454
rect 49928 39134 50248 39218
rect 49928 38898 49970 39134
rect 50206 38898 50248 39134
rect 49928 38866 50248 38898
rect 80648 39454 80968 39486
rect 80648 39218 80690 39454
rect 80926 39218 80968 39454
rect 80648 39134 80968 39218
rect 80648 38898 80690 39134
rect 80926 38898 80968 39134
rect 80648 38866 80968 38898
rect 111368 39454 111688 39486
rect 111368 39218 111410 39454
rect 111646 39218 111688 39454
rect 111368 39134 111688 39218
rect 111368 38898 111410 39134
rect 111646 38898 111688 39134
rect 111368 38866 111688 38898
rect 142088 39454 142408 39486
rect 142088 39218 142130 39454
rect 142366 39218 142408 39454
rect 142088 39134 142408 39218
rect 142088 38898 142130 39134
rect 142366 38898 142408 39134
rect 142088 38866 142408 38898
rect 172808 39454 173128 39486
rect 172808 39218 172850 39454
rect 173086 39218 173128 39454
rect 172808 39134 173128 39218
rect 172808 38898 172850 39134
rect 173086 38898 173128 39134
rect 172808 38866 173128 38898
rect 203528 39454 203848 39486
rect 203528 39218 203570 39454
rect 203806 39218 203848 39454
rect 203528 39134 203848 39218
rect 203528 38898 203570 39134
rect 203806 38898 203848 39134
rect 203528 38866 203848 38898
rect 234248 39454 234568 39486
rect 234248 39218 234290 39454
rect 234526 39218 234568 39454
rect 234248 39134 234568 39218
rect 234248 38898 234290 39134
rect 234526 38898 234568 39134
rect 234248 38866 234568 38898
rect 264968 39454 265288 39486
rect 264968 39218 265010 39454
rect 265246 39218 265288 39454
rect 264968 39134 265288 39218
rect 264968 38898 265010 39134
rect 265246 38898 265288 39134
rect 264968 38866 265288 38898
rect 295688 39454 296008 39486
rect 295688 39218 295730 39454
rect 295966 39218 296008 39454
rect 295688 39134 296008 39218
rect 295688 38898 295730 39134
rect 295966 38898 296008 39134
rect 295688 38866 296008 38898
rect 326408 39454 326728 39486
rect 326408 39218 326450 39454
rect 326686 39218 326728 39454
rect 326408 39134 326728 39218
rect 326408 38898 326450 39134
rect 326686 38898 326728 39134
rect 326408 38866 326728 38898
rect 357128 39454 357448 39486
rect 357128 39218 357170 39454
rect 357406 39218 357448 39454
rect 357128 39134 357448 39218
rect 357128 38898 357170 39134
rect 357406 38898 357448 39134
rect 357128 38866 357448 38898
rect 387848 39454 388168 39486
rect 387848 39218 387890 39454
rect 388126 39218 388168 39454
rect 387848 39134 388168 39218
rect 387848 38898 387890 39134
rect 388126 38898 388168 39134
rect 387848 38866 388168 38898
rect 418568 39454 418888 39486
rect 418568 39218 418610 39454
rect 418846 39218 418888 39454
rect 418568 39134 418888 39218
rect 418568 38898 418610 39134
rect 418846 38898 418888 39134
rect 418568 38866 418888 38898
rect 449288 39454 449608 39486
rect 449288 39218 449330 39454
rect 449566 39218 449608 39454
rect 449288 39134 449608 39218
rect 449288 38898 449330 39134
rect 449566 38898 449608 39134
rect 449288 38866 449608 38898
rect 480008 39454 480328 39486
rect 480008 39218 480050 39454
rect 480286 39218 480328 39454
rect 480008 39134 480328 39218
rect 480008 38898 480050 39134
rect 480286 38898 480328 39134
rect 480008 38866 480328 38898
rect 510728 39454 511048 39486
rect 510728 39218 510770 39454
rect 511006 39218 511048 39454
rect 510728 39134 511048 39218
rect 510728 38898 510770 39134
rect 511006 38898 511048 39134
rect 510728 38866 511048 38898
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 34568 21454 34888 21486
rect 34568 21218 34610 21454
rect 34846 21218 34888 21454
rect 34568 21134 34888 21218
rect 34568 20898 34610 21134
rect 34846 20898 34888 21134
rect 34568 20866 34888 20898
rect 65288 21454 65608 21486
rect 65288 21218 65330 21454
rect 65566 21218 65608 21454
rect 65288 21134 65608 21218
rect 65288 20898 65330 21134
rect 65566 20898 65608 21134
rect 65288 20866 65608 20898
rect 96008 21454 96328 21486
rect 96008 21218 96050 21454
rect 96286 21218 96328 21454
rect 96008 21134 96328 21218
rect 96008 20898 96050 21134
rect 96286 20898 96328 21134
rect 96008 20866 96328 20898
rect 126728 21454 127048 21486
rect 126728 21218 126770 21454
rect 127006 21218 127048 21454
rect 126728 21134 127048 21218
rect 126728 20898 126770 21134
rect 127006 20898 127048 21134
rect 126728 20866 127048 20898
rect 157448 21454 157768 21486
rect 157448 21218 157490 21454
rect 157726 21218 157768 21454
rect 157448 21134 157768 21218
rect 157448 20898 157490 21134
rect 157726 20898 157768 21134
rect 157448 20866 157768 20898
rect 188168 21454 188488 21486
rect 188168 21218 188210 21454
rect 188446 21218 188488 21454
rect 188168 21134 188488 21218
rect 188168 20898 188210 21134
rect 188446 20898 188488 21134
rect 188168 20866 188488 20898
rect 218888 21454 219208 21486
rect 218888 21218 218930 21454
rect 219166 21218 219208 21454
rect 218888 21134 219208 21218
rect 218888 20898 218930 21134
rect 219166 20898 219208 21134
rect 218888 20866 219208 20898
rect 249608 21454 249928 21486
rect 249608 21218 249650 21454
rect 249886 21218 249928 21454
rect 249608 21134 249928 21218
rect 249608 20898 249650 21134
rect 249886 20898 249928 21134
rect 249608 20866 249928 20898
rect 280328 21454 280648 21486
rect 280328 21218 280370 21454
rect 280606 21218 280648 21454
rect 280328 21134 280648 21218
rect 280328 20898 280370 21134
rect 280606 20898 280648 21134
rect 280328 20866 280648 20898
rect 311048 21454 311368 21486
rect 311048 21218 311090 21454
rect 311326 21218 311368 21454
rect 311048 21134 311368 21218
rect 311048 20898 311090 21134
rect 311326 20898 311368 21134
rect 311048 20866 311368 20898
rect 341768 21454 342088 21486
rect 341768 21218 341810 21454
rect 342046 21218 342088 21454
rect 341768 21134 342088 21218
rect 341768 20898 341810 21134
rect 342046 20898 342088 21134
rect 341768 20866 342088 20898
rect 372488 21454 372808 21486
rect 372488 21218 372530 21454
rect 372766 21218 372808 21454
rect 372488 21134 372808 21218
rect 372488 20898 372530 21134
rect 372766 20898 372808 21134
rect 372488 20866 372808 20898
rect 403208 21454 403528 21486
rect 403208 21218 403250 21454
rect 403486 21218 403528 21454
rect 403208 21134 403528 21218
rect 403208 20898 403250 21134
rect 403486 20898 403528 21134
rect 403208 20866 403528 20898
rect 433928 21454 434248 21486
rect 433928 21218 433970 21454
rect 434206 21218 434248 21454
rect 433928 21134 434248 21218
rect 433928 20898 433970 21134
rect 434206 20898 434248 21134
rect 433928 20866 434248 20898
rect 464648 21454 464968 21486
rect 464648 21218 464690 21454
rect 464926 21218 464968 21454
rect 464648 21134 464968 21218
rect 464648 20898 464690 21134
rect 464926 20898 464968 21134
rect 464648 20866 464968 20898
rect 495368 21454 495688 21486
rect 495368 21218 495410 21454
rect 495646 21218 495688 21454
rect 495368 21134 495688 21218
rect 495368 20898 495410 21134
rect 495646 20898 495688 21134
rect 495368 20866 495688 20898
rect 526088 21454 526408 21486
rect 526088 21218 526130 21454
rect 526366 21218 526408 21454
rect 526088 21134 526408 21218
rect 526088 20898 526130 21134
rect 526366 20898 526408 21134
rect 526088 20866 526408 20898
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 13000
rect 19794 -1306 20414 13000
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 -3226 24134 13000
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 -5146 27854 13000
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 13000
rect 37794 3454 38414 13000
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 7174 42134 13000
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 10894 45854 13000
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 13000
rect 55794 -1306 56414 13000
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 -3226 60134 13000
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 -5146 63854 13000
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 13000
rect 73794 3454 74414 13000
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 7174 78134 13000
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 10894 81854 13000
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 13000
rect 91794 -1306 92414 13000
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 -3226 96134 13000
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 -5146 99854 13000
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 13000
rect 109794 3454 110414 13000
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 7174 114134 13000
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 10894 117854 13000
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 13000
rect 127794 -1306 128414 13000
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 -3226 132134 13000
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 -5146 135854 13000
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 13000
rect 145794 3454 146414 13000
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 7174 150134 13000
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 10894 153854 13000
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 13000
rect 163794 -1306 164414 13000
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 -3226 168134 13000
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 -5146 171854 13000
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 13000
rect 181794 3454 182414 13000
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 7174 186134 13000
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 10894 189854 13000
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 13000
rect 199794 -1306 200414 13000
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 -3226 204134 13000
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 -5146 207854 13000
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 13000
rect 217794 3454 218414 13000
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 7174 222134 13000
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 10894 225854 13000
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 13000
rect 235794 -1306 236414 13000
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 -3226 240134 13000
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 -5146 243854 13000
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 13000
rect 253794 3454 254414 13000
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 7174 258134 13000
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 10894 261854 13000
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 13000
rect 271794 -1306 272414 13000
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 -3226 276134 13000
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 -5146 279854 13000
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 13000
rect 289794 3454 290414 13000
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 7174 294134 13000
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 10894 297854 13000
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 13000
rect 307794 -1306 308414 13000
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 -3226 312134 13000
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 -5146 315854 13000
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 13000
rect 325794 3454 326414 13000
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 7174 330134 13000
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 10894 333854 13000
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 13000
rect 343794 -1306 344414 13000
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 -3226 348134 13000
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 -5146 351854 13000
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 13000
rect 361794 3454 362414 13000
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 7174 366134 13000
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 10894 369854 13000
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 13000
rect 379794 -1306 380414 13000
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 -3226 384134 13000
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 -5146 387854 13000
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 13000
rect 397794 3454 398414 13000
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 7174 402134 13000
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 10894 405854 13000
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 13000
rect 415794 -1306 416414 13000
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 -3226 420134 13000
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 -5146 423854 13000
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 13000
rect 433794 3454 434414 13000
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 7174 438134 13000
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 10894 441854 13000
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 13000
rect 451794 -1306 452414 13000
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 -3226 456134 13000
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 -5146 459854 13000
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 13000
rect 469794 3454 470414 13000
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 7174 474134 13000
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 10894 477854 13000
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 13000
rect 487794 -1306 488414 13000
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 -3226 492134 13000
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 -5146 495854 13000
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 13000
rect 505794 3454 506414 13000
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 7174 510134 13000
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 10894 513854 13000
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 13000
rect 523794 -1306 524414 13000
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 -3226 528134 13000
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 -5146 531854 13000
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 13000
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 19250 651218 19486 651454
rect 19250 650898 19486 651134
rect 49970 651218 50206 651454
rect 49970 650898 50206 651134
rect 80690 651218 80926 651454
rect 80690 650898 80926 651134
rect 111410 651218 111646 651454
rect 111410 650898 111646 651134
rect 142130 651218 142366 651454
rect 142130 650898 142366 651134
rect 172850 651218 173086 651454
rect 172850 650898 173086 651134
rect 203570 651218 203806 651454
rect 203570 650898 203806 651134
rect 234290 651218 234526 651454
rect 234290 650898 234526 651134
rect 265010 651218 265246 651454
rect 265010 650898 265246 651134
rect 295730 651218 295966 651454
rect 295730 650898 295966 651134
rect 326450 651218 326686 651454
rect 326450 650898 326686 651134
rect 357170 651218 357406 651454
rect 357170 650898 357406 651134
rect 387890 651218 388126 651454
rect 387890 650898 388126 651134
rect 418610 651218 418846 651454
rect 418610 650898 418846 651134
rect 449330 651218 449566 651454
rect 449330 650898 449566 651134
rect 480050 651218 480286 651454
rect 480050 650898 480286 651134
rect 510770 651218 511006 651454
rect 510770 650898 511006 651134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 34610 633218 34846 633454
rect 34610 632898 34846 633134
rect 65330 633218 65566 633454
rect 65330 632898 65566 633134
rect 96050 633218 96286 633454
rect 96050 632898 96286 633134
rect 126770 633218 127006 633454
rect 126770 632898 127006 633134
rect 157490 633218 157726 633454
rect 157490 632898 157726 633134
rect 188210 633218 188446 633454
rect 188210 632898 188446 633134
rect 218930 633218 219166 633454
rect 218930 632898 219166 633134
rect 249650 633218 249886 633454
rect 249650 632898 249886 633134
rect 280370 633218 280606 633454
rect 280370 632898 280606 633134
rect 311090 633218 311326 633454
rect 311090 632898 311326 633134
rect 341810 633218 342046 633454
rect 341810 632898 342046 633134
rect 372530 633218 372766 633454
rect 372530 632898 372766 633134
rect 403250 633218 403486 633454
rect 403250 632898 403486 633134
rect 433970 633218 434206 633454
rect 433970 632898 434206 633134
rect 464690 633218 464926 633454
rect 464690 632898 464926 633134
rect 495410 633218 495646 633454
rect 495410 632898 495646 633134
rect 526130 633218 526366 633454
rect 526130 632898 526366 633134
rect 19250 615218 19486 615454
rect 19250 614898 19486 615134
rect 49970 615218 50206 615454
rect 49970 614898 50206 615134
rect 80690 615218 80926 615454
rect 80690 614898 80926 615134
rect 111410 615218 111646 615454
rect 111410 614898 111646 615134
rect 142130 615218 142366 615454
rect 142130 614898 142366 615134
rect 172850 615218 173086 615454
rect 172850 614898 173086 615134
rect 203570 615218 203806 615454
rect 203570 614898 203806 615134
rect 234290 615218 234526 615454
rect 234290 614898 234526 615134
rect 265010 615218 265246 615454
rect 265010 614898 265246 615134
rect 295730 615218 295966 615454
rect 295730 614898 295966 615134
rect 326450 615218 326686 615454
rect 326450 614898 326686 615134
rect 357170 615218 357406 615454
rect 357170 614898 357406 615134
rect 387890 615218 388126 615454
rect 387890 614898 388126 615134
rect 418610 615218 418846 615454
rect 418610 614898 418846 615134
rect 449330 615218 449566 615454
rect 449330 614898 449566 615134
rect 480050 615218 480286 615454
rect 480050 614898 480286 615134
rect 510770 615218 511006 615454
rect 510770 614898 511006 615134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 34610 597218 34846 597454
rect 34610 596898 34846 597134
rect 65330 597218 65566 597454
rect 65330 596898 65566 597134
rect 96050 597218 96286 597454
rect 96050 596898 96286 597134
rect 126770 597218 127006 597454
rect 126770 596898 127006 597134
rect 157490 597218 157726 597454
rect 157490 596898 157726 597134
rect 188210 597218 188446 597454
rect 188210 596898 188446 597134
rect 218930 597218 219166 597454
rect 218930 596898 219166 597134
rect 249650 597218 249886 597454
rect 249650 596898 249886 597134
rect 280370 597218 280606 597454
rect 280370 596898 280606 597134
rect 311090 597218 311326 597454
rect 311090 596898 311326 597134
rect 341810 597218 342046 597454
rect 341810 596898 342046 597134
rect 372530 597218 372766 597454
rect 372530 596898 372766 597134
rect 403250 597218 403486 597454
rect 403250 596898 403486 597134
rect 433970 597218 434206 597454
rect 433970 596898 434206 597134
rect 464690 597218 464926 597454
rect 464690 596898 464926 597134
rect 495410 597218 495646 597454
rect 495410 596898 495646 597134
rect 526130 597218 526366 597454
rect 526130 596898 526366 597134
rect 19250 579218 19486 579454
rect 19250 578898 19486 579134
rect 49970 579218 50206 579454
rect 49970 578898 50206 579134
rect 80690 579218 80926 579454
rect 80690 578898 80926 579134
rect 111410 579218 111646 579454
rect 111410 578898 111646 579134
rect 142130 579218 142366 579454
rect 142130 578898 142366 579134
rect 172850 579218 173086 579454
rect 172850 578898 173086 579134
rect 203570 579218 203806 579454
rect 203570 578898 203806 579134
rect 234290 579218 234526 579454
rect 234290 578898 234526 579134
rect 265010 579218 265246 579454
rect 265010 578898 265246 579134
rect 295730 579218 295966 579454
rect 295730 578898 295966 579134
rect 326450 579218 326686 579454
rect 326450 578898 326686 579134
rect 357170 579218 357406 579454
rect 357170 578898 357406 579134
rect 387890 579218 388126 579454
rect 387890 578898 388126 579134
rect 418610 579218 418846 579454
rect 418610 578898 418846 579134
rect 449330 579218 449566 579454
rect 449330 578898 449566 579134
rect 480050 579218 480286 579454
rect 480050 578898 480286 579134
rect 510770 579218 511006 579454
rect 510770 578898 511006 579134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 34610 561218 34846 561454
rect 34610 560898 34846 561134
rect 65330 561218 65566 561454
rect 65330 560898 65566 561134
rect 96050 561218 96286 561454
rect 96050 560898 96286 561134
rect 126770 561218 127006 561454
rect 126770 560898 127006 561134
rect 157490 561218 157726 561454
rect 157490 560898 157726 561134
rect 188210 561218 188446 561454
rect 188210 560898 188446 561134
rect 218930 561218 219166 561454
rect 218930 560898 219166 561134
rect 249650 561218 249886 561454
rect 249650 560898 249886 561134
rect 280370 561218 280606 561454
rect 280370 560898 280606 561134
rect 311090 561218 311326 561454
rect 311090 560898 311326 561134
rect 341810 561218 342046 561454
rect 341810 560898 342046 561134
rect 372530 561218 372766 561454
rect 372530 560898 372766 561134
rect 403250 561218 403486 561454
rect 403250 560898 403486 561134
rect 433970 561218 434206 561454
rect 433970 560898 434206 561134
rect 464690 561218 464926 561454
rect 464690 560898 464926 561134
rect 495410 561218 495646 561454
rect 495410 560898 495646 561134
rect 526130 561218 526366 561454
rect 526130 560898 526366 561134
rect 19250 543218 19486 543454
rect 19250 542898 19486 543134
rect 49970 543218 50206 543454
rect 49970 542898 50206 543134
rect 80690 543218 80926 543454
rect 80690 542898 80926 543134
rect 111410 543218 111646 543454
rect 111410 542898 111646 543134
rect 142130 543218 142366 543454
rect 142130 542898 142366 543134
rect 172850 543218 173086 543454
rect 172850 542898 173086 543134
rect 203570 543218 203806 543454
rect 203570 542898 203806 543134
rect 234290 543218 234526 543454
rect 234290 542898 234526 543134
rect 265010 543218 265246 543454
rect 265010 542898 265246 543134
rect 295730 543218 295966 543454
rect 295730 542898 295966 543134
rect 326450 543218 326686 543454
rect 326450 542898 326686 543134
rect 357170 543218 357406 543454
rect 357170 542898 357406 543134
rect 387890 543218 388126 543454
rect 387890 542898 388126 543134
rect 418610 543218 418846 543454
rect 418610 542898 418846 543134
rect 449330 543218 449566 543454
rect 449330 542898 449566 543134
rect 480050 543218 480286 543454
rect 480050 542898 480286 543134
rect 510770 543218 511006 543454
rect 510770 542898 511006 543134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 34610 525218 34846 525454
rect 34610 524898 34846 525134
rect 65330 525218 65566 525454
rect 65330 524898 65566 525134
rect 96050 525218 96286 525454
rect 96050 524898 96286 525134
rect 126770 525218 127006 525454
rect 126770 524898 127006 525134
rect 157490 525218 157726 525454
rect 157490 524898 157726 525134
rect 188210 525218 188446 525454
rect 188210 524898 188446 525134
rect 218930 525218 219166 525454
rect 218930 524898 219166 525134
rect 249650 525218 249886 525454
rect 249650 524898 249886 525134
rect 280370 525218 280606 525454
rect 280370 524898 280606 525134
rect 311090 525218 311326 525454
rect 311090 524898 311326 525134
rect 341810 525218 342046 525454
rect 341810 524898 342046 525134
rect 372530 525218 372766 525454
rect 372530 524898 372766 525134
rect 403250 525218 403486 525454
rect 403250 524898 403486 525134
rect 433970 525218 434206 525454
rect 433970 524898 434206 525134
rect 464690 525218 464926 525454
rect 464690 524898 464926 525134
rect 495410 525218 495646 525454
rect 495410 524898 495646 525134
rect 526130 525218 526366 525454
rect 526130 524898 526366 525134
rect 19250 507218 19486 507454
rect 19250 506898 19486 507134
rect 49970 507218 50206 507454
rect 49970 506898 50206 507134
rect 80690 507218 80926 507454
rect 80690 506898 80926 507134
rect 111410 507218 111646 507454
rect 111410 506898 111646 507134
rect 142130 507218 142366 507454
rect 142130 506898 142366 507134
rect 172850 507218 173086 507454
rect 172850 506898 173086 507134
rect 203570 507218 203806 507454
rect 203570 506898 203806 507134
rect 234290 507218 234526 507454
rect 234290 506898 234526 507134
rect 265010 507218 265246 507454
rect 265010 506898 265246 507134
rect 295730 507218 295966 507454
rect 295730 506898 295966 507134
rect 326450 507218 326686 507454
rect 326450 506898 326686 507134
rect 357170 507218 357406 507454
rect 357170 506898 357406 507134
rect 387890 507218 388126 507454
rect 387890 506898 388126 507134
rect 418610 507218 418846 507454
rect 418610 506898 418846 507134
rect 449330 507218 449566 507454
rect 449330 506898 449566 507134
rect 480050 507218 480286 507454
rect 480050 506898 480286 507134
rect 510770 507218 511006 507454
rect 510770 506898 511006 507134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 34610 489218 34846 489454
rect 34610 488898 34846 489134
rect 65330 489218 65566 489454
rect 65330 488898 65566 489134
rect 96050 489218 96286 489454
rect 96050 488898 96286 489134
rect 126770 489218 127006 489454
rect 126770 488898 127006 489134
rect 157490 489218 157726 489454
rect 157490 488898 157726 489134
rect 188210 489218 188446 489454
rect 188210 488898 188446 489134
rect 218930 489218 219166 489454
rect 218930 488898 219166 489134
rect 249650 489218 249886 489454
rect 249650 488898 249886 489134
rect 280370 489218 280606 489454
rect 280370 488898 280606 489134
rect 311090 489218 311326 489454
rect 311090 488898 311326 489134
rect 341810 489218 342046 489454
rect 341810 488898 342046 489134
rect 372530 489218 372766 489454
rect 372530 488898 372766 489134
rect 403250 489218 403486 489454
rect 403250 488898 403486 489134
rect 433970 489218 434206 489454
rect 433970 488898 434206 489134
rect 464690 489218 464926 489454
rect 464690 488898 464926 489134
rect 495410 489218 495646 489454
rect 495410 488898 495646 489134
rect 526130 489218 526366 489454
rect 526130 488898 526366 489134
rect 19250 471218 19486 471454
rect 19250 470898 19486 471134
rect 49970 471218 50206 471454
rect 49970 470898 50206 471134
rect 80690 471218 80926 471454
rect 80690 470898 80926 471134
rect 111410 471218 111646 471454
rect 111410 470898 111646 471134
rect 142130 471218 142366 471454
rect 142130 470898 142366 471134
rect 172850 471218 173086 471454
rect 172850 470898 173086 471134
rect 203570 471218 203806 471454
rect 203570 470898 203806 471134
rect 234290 471218 234526 471454
rect 234290 470898 234526 471134
rect 265010 471218 265246 471454
rect 265010 470898 265246 471134
rect 295730 471218 295966 471454
rect 295730 470898 295966 471134
rect 326450 471218 326686 471454
rect 326450 470898 326686 471134
rect 357170 471218 357406 471454
rect 357170 470898 357406 471134
rect 387890 471218 388126 471454
rect 387890 470898 388126 471134
rect 418610 471218 418846 471454
rect 418610 470898 418846 471134
rect 449330 471218 449566 471454
rect 449330 470898 449566 471134
rect 480050 471218 480286 471454
rect 480050 470898 480286 471134
rect 510770 471218 511006 471454
rect 510770 470898 511006 471134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 34610 453218 34846 453454
rect 34610 452898 34846 453134
rect 65330 453218 65566 453454
rect 65330 452898 65566 453134
rect 96050 453218 96286 453454
rect 96050 452898 96286 453134
rect 126770 453218 127006 453454
rect 126770 452898 127006 453134
rect 157490 453218 157726 453454
rect 157490 452898 157726 453134
rect 188210 453218 188446 453454
rect 188210 452898 188446 453134
rect 218930 453218 219166 453454
rect 218930 452898 219166 453134
rect 249650 453218 249886 453454
rect 249650 452898 249886 453134
rect 280370 453218 280606 453454
rect 280370 452898 280606 453134
rect 311090 453218 311326 453454
rect 311090 452898 311326 453134
rect 341810 453218 342046 453454
rect 341810 452898 342046 453134
rect 372530 453218 372766 453454
rect 372530 452898 372766 453134
rect 403250 453218 403486 453454
rect 403250 452898 403486 453134
rect 433970 453218 434206 453454
rect 433970 452898 434206 453134
rect 464690 453218 464926 453454
rect 464690 452898 464926 453134
rect 495410 453218 495646 453454
rect 495410 452898 495646 453134
rect 526130 453218 526366 453454
rect 526130 452898 526366 453134
rect 19250 435218 19486 435454
rect 19250 434898 19486 435134
rect 49970 435218 50206 435454
rect 49970 434898 50206 435134
rect 80690 435218 80926 435454
rect 80690 434898 80926 435134
rect 111410 435218 111646 435454
rect 111410 434898 111646 435134
rect 142130 435218 142366 435454
rect 142130 434898 142366 435134
rect 172850 435218 173086 435454
rect 172850 434898 173086 435134
rect 203570 435218 203806 435454
rect 203570 434898 203806 435134
rect 234290 435218 234526 435454
rect 234290 434898 234526 435134
rect 265010 435218 265246 435454
rect 265010 434898 265246 435134
rect 295730 435218 295966 435454
rect 295730 434898 295966 435134
rect 326450 435218 326686 435454
rect 326450 434898 326686 435134
rect 357170 435218 357406 435454
rect 357170 434898 357406 435134
rect 387890 435218 388126 435454
rect 387890 434898 388126 435134
rect 418610 435218 418846 435454
rect 418610 434898 418846 435134
rect 449330 435218 449566 435454
rect 449330 434898 449566 435134
rect 480050 435218 480286 435454
rect 480050 434898 480286 435134
rect 510770 435218 511006 435454
rect 510770 434898 511006 435134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 34610 417218 34846 417454
rect 34610 416898 34846 417134
rect 65330 417218 65566 417454
rect 65330 416898 65566 417134
rect 96050 417218 96286 417454
rect 96050 416898 96286 417134
rect 126770 417218 127006 417454
rect 126770 416898 127006 417134
rect 157490 417218 157726 417454
rect 157490 416898 157726 417134
rect 188210 417218 188446 417454
rect 188210 416898 188446 417134
rect 218930 417218 219166 417454
rect 218930 416898 219166 417134
rect 249650 417218 249886 417454
rect 249650 416898 249886 417134
rect 280370 417218 280606 417454
rect 280370 416898 280606 417134
rect 311090 417218 311326 417454
rect 311090 416898 311326 417134
rect 341810 417218 342046 417454
rect 341810 416898 342046 417134
rect 372530 417218 372766 417454
rect 372530 416898 372766 417134
rect 403250 417218 403486 417454
rect 403250 416898 403486 417134
rect 433970 417218 434206 417454
rect 433970 416898 434206 417134
rect 464690 417218 464926 417454
rect 464690 416898 464926 417134
rect 495410 417218 495646 417454
rect 495410 416898 495646 417134
rect 526130 417218 526366 417454
rect 526130 416898 526366 417134
rect 19250 399218 19486 399454
rect 19250 398898 19486 399134
rect 49970 399218 50206 399454
rect 49970 398898 50206 399134
rect 80690 399218 80926 399454
rect 80690 398898 80926 399134
rect 111410 399218 111646 399454
rect 111410 398898 111646 399134
rect 142130 399218 142366 399454
rect 142130 398898 142366 399134
rect 172850 399218 173086 399454
rect 172850 398898 173086 399134
rect 203570 399218 203806 399454
rect 203570 398898 203806 399134
rect 234290 399218 234526 399454
rect 234290 398898 234526 399134
rect 265010 399218 265246 399454
rect 265010 398898 265246 399134
rect 295730 399218 295966 399454
rect 295730 398898 295966 399134
rect 326450 399218 326686 399454
rect 326450 398898 326686 399134
rect 357170 399218 357406 399454
rect 357170 398898 357406 399134
rect 387890 399218 388126 399454
rect 387890 398898 388126 399134
rect 418610 399218 418846 399454
rect 418610 398898 418846 399134
rect 449330 399218 449566 399454
rect 449330 398898 449566 399134
rect 480050 399218 480286 399454
rect 480050 398898 480286 399134
rect 510770 399218 511006 399454
rect 510770 398898 511006 399134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 34610 381218 34846 381454
rect 34610 380898 34846 381134
rect 65330 381218 65566 381454
rect 65330 380898 65566 381134
rect 96050 381218 96286 381454
rect 96050 380898 96286 381134
rect 126770 381218 127006 381454
rect 126770 380898 127006 381134
rect 157490 381218 157726 381454
rect 157490 380898 157726 381134
rect 188210 381218 188446 381454
rect 188210 380898 188446 381134
rect 218930 381218 219166 381454
rect 218930 380898 219166 381134
rect 249650 381218 249886 381454
rect 249650 380898 249886 381134
rect 280370 381218 280606 381454
rect 280370 380898 280606 381134
rect 311090 381218 311326 381454
rect 311090 380898 311326 381134
rect 341810 381218 342046 381454
rect 341810 380898 342046 381134
rect 372530 381218 372766 381454
rect 372530 380898 372766 381134
rect 403250 381218 403486 381454
rect 403250 380898 403486 381134
rect 433970 381218 434206 381454
rect 433970 380898 434206 381134
rect 464690 381218 464926 381454
rect 464690 380898 464926 381134
rect 495410 381218 495646 381454
rect 495410 380898 495646 381134
rect 526130 381218 526366 381454
rect 526130 380898 526366 381134
rect 19250 363218 19486 363454
rect 19250 362898 19486 363134
rect 49970 363218 50206 363454
rect 49970 362898 50206 363134
rect 80690 363218 80926 363454
rect 80690 362898 80926 363134
rect 111410 363218 111646 363454
rect 111410 362898 111646 363134
rect 142130 363218 142366 363454
rect 142130 362898 142366 363134
rect 172850 363218 173086 363454
rect 172850 362898 173086 363134
rect 203570 363218 203806 363454
rect 203570 362898 203806 363134
rect 234290 363218 234526 363454
rect 234290 362898 234526 363134
rect 265010 363218 265246 363454
rect 265010 362898 265246 363134
rect 295730 363218 295966 363454
rect 295730 362898 295966 363134
rect 326450 363218 326686 363454
rect 326450 362898 326686 363134
rect 357170 363218 357406 363454
rect 357170 362898 357406 363134
rect 387890 363218 388126 363454
rect 387890 362898 388126 363134
rect 418610 363218 418846 363454
rect 418610 362898 418846 363134
rect 449330 363218 449566 363454
rect 449330 362898 449566 363134
rect 480050 363218 480286 363454
rect 480050 362898 480286 363134
rect 510770 363218 511006 363454
rect 510770 362898 511006 363134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 34610 345218 34846 345454
rect 34610 344898 34846 345134
rect 65330 345218 65566 345454
rect 65330 344898 65566 345134
rect 96050 345218 96286 345454
rect 96050 344898 96286 345134
rect 126770 345218 127006 345454
rect 126770 344898 127006 345134
rect 157490 345218 157726 345454
rect 157490 344898 157726 345134
rect 188210 345218 188446 345454
rect 188210 344898 188446 345134
rect 218930 345218 219166 345454
rect 218930 344898 219166 345134
rect 249650 345218 249886 345454
rect 249650 344898 249886 345134
rect 280370 345218 280606 345454
rect 280370 344898 280606 345134
rect 311090 345218 311326 345454
rect 311090 344898 311326 345134
rect 341810 345218 342046 345454
rect 341810 344898 342046 345134
rect 372530 345218 372766 345454
rect 372530 344898 372766 345134
rect 403250 345218 403486 345454
rect 403250 344898 403486 345134
rect 433970 345218 434206 345454
rect 433970 344898 434206 345134
rect 464690 345218 464926 345454
rect 464690 344898 464926 345134
rect 495410 345218 495646 345454
rect 495410 344898 495646 345134
rect 526130 345218 526366 345454
rect 526130 344898 526366 345134
rect 19250 327218 19486 327454
rect 19250 326898 19486 327134
rect 49970 327218 50206 327454
rect 49970 326898 50206 327134
rect 80690 327218 80926 327454
rect 80690 326898 80926 327134
rect 111410 327218 111646 327454
rect 111410 326898 111646 327134
rect 142130 327218 142366 327454
rect 142130 326898 142366 327134
rect 172850 327218 173086 327454
rect 172850 326898 173086 327134
rect 203570 327218 203806 327454
rect 203570 326898 203806 327134
rect 234290 327218 234526 327454
rect 234290 326898 234526 327134
rect 265010 327218 265246 327454
rect 265010 326898 265246 327134
rect 295730 327218 295966 327454
rect 295730 326898 295966 327134
rect 326450 327218 326686 327454
rect 326450 326898 326686 327134
rect 357170 327218 357406 327454
rect 357170 326898 357406 327134
rect 387890 327218 388126 327454
rect 387890 326898 388126 327134
rect 418610 327218 418846 327454
rect 418610 326898 418846 327134
rect 449330 327218 449566 327454
rect 449330 326898 449566 327134
rect 480050 327218 480286 327454
rect 480050 326898 480286 327134
rect 510770 327218 511006 327454
rect 510770 326898 511006 327134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 34610 309218 34846 309454
rect 34610 308898 34846 309134
rect 65330 309218 65566 309454
rect 65330 308898 65566 309134
rect 96050 309218 96286 309454
rect 96050 308898 96286 309134
rect 126770 309218 127006 309454
rect 126770 308898 127006 309134
rect 157490 309218 157726 309454
rect 157490 308898 157726 309134
rect 188210 309218 188446 309454
rect 188210 308898 188446 309134
rect 218930 309218 219166 309454
rect 218930 308898 219166 309134
rect 249650 309218 249886 309454
rect 249650 308898 249886 309134
rect 280370 309218 280606 309454
rect 280370 308898 280606 309134
rect 311090 309218 311326 309454
rect 311090 308898 311326 309134
rect 341810 309218 342046 309454
rect 341810 308898 342046 309134
rect 372530 309218 372766 309454
rect 372530 308898 372766 309134
rect 403250 309218 403486 309454
rect 403250 308898 403486 309134
rect 433970 309218 434206 309454
rect 433970 308898 434206 309134
rect 464690 309218 464926 309454
rect 464690 308898 464926 309134
rect 495410 309218 495646 309454
rect 495410 308898 495646 309134
rect 526130 309218 526366 309454
rect 526130 308898 526366 309134
rect 19250 291218 19486 291454
rect 19250 290898 19486 291134
rect 49970 291218 50206 291454
rect 49970 290898 50206 291134
rect 80690 291218 80926 291454
rect 80690 290898 80926 291134
rect 111410 291218 111646 291454
rect 111410 290898 111646 291134
rect 142130 291218 142366 291454
rect 142130 290898 142366 291134
rect 172850 291218 173086 291454
rect 172850 290898 173086 291134
rect 203570 291218 203806 291454
rect 203570 290898 203806 291134
rect 234290 291218 234526 291454
rect 234290 290898 234526 291134
rect 265010 291218 265246 291454
rect 265010 290898 265246 291134
rect 295730 291218 295966 291454
rect 295730 290898 295966 291134
rect 326450 291218 326686 291454
rect 326450 290898 326686 291134
rect 357170 291218 357406 291454
rect 357170 290898 357406 291134
rect 387890 291218 388126 291454
rect 387890 290898 388126 291134
rect 418610 291218 418846 291454
rect 418610 290898 418846 291134
rect 449330 291218 449566 291454
rect 449330 290898 449566 291134
rect 480050 291218 480286 291454
rect 480050 290898 480286 291134
rect 510770 291218 511006 291454
rect 510770 290898 511006 291134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 34610 273218 34846 273454
rect 34610 272898 34846 273134
rect 65330 273218 65566 273454
rect 65330 272898 65566 273134
rect 96050 273218 96286 273454
rect 96050 272898 96286 273134
rect 126770 273218 127006 273454
rect 126770 272898 127006 273134
rect 157490 273218 157726 273454
rect 157490 272898 157726 273134
rect 188210 273218 188446 273454
rect 188210 272898 188446 273134
rect 218930 273218 219166 273454
rect 218930 272898 219166 273134
rect 249650 273218 249886 273454
rect 249650 272898 249886 273134
rect 280370 273218 280606 273454
rect 280370 272898 280606 273134
rect 311090 273218 311326 273454
rect 311090 272898 311326 273134
rect 341810 273218 342046 273454
rect 341810 272898 342046 273134
rect 372530 273218 372766 273454
rect 372530 272898 372766 273134
rect 403250 273218 403486 273454
rect 403250 272898 403486 273134
rect 433970 273218 434206 273454
rect 433970 272898 434206 273134
rect 464690 273218 464926 273454
rect 464690 272898 464926 273134
rect 495410 273218 495646 273454
rect 495410 272898 495646 273134
rect 526130 273218 526366 273454
rect 526130 272898 526366 273134
rect 19250 255218 19486 255454
rect 19250 254898 19486 255134
rect 49970 255218 50206 255454
rect 49970 254898 50206 255134
rect 80690 255218 80926 255454
rect 80690 254898 80926 255134
rect 111410 255218 111646 255454
rect 111410 254898 111646 255134
rect 142130 255218 142366 255454
rect 142130 254898 142366 255134
rect 172850 255218 173086 255454
rect 172850 254898 173086 255134
rect 203570 255218 203806 255454
rect 203570 254898 203806 255134
rect 234290 255218 234526 255454
rect 234290 254898 234526 255134
rect 265010 255218 265246 255454
rect 265010 254898 265246 255134
rect 295730 255218 295966 255454
rect 295730 254898 295966 255134
rect 326450 255218 326686 255454
rect 326450 254898 326686 255134
rect 357170 255218 357406 255454
rect 357170 254898 357406 255134
rect 387890 255218 388126 255454
rect 387890 254898 388126 255134
rect 418610 255218 418846 255454
rect 418610 254898 418846 255134
rect 449330 255218 449566 255454
rect 449330 254898 449566 255134
rect 480050 255218 480286 255454
rect 480050 254898 480286 255134
rect 510770 255218 511006 255454
rect 510770 254898 511006 255134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 34610 237218 34846 237454
rect 34610 236898 34846 237134
rect 65330 237218 65566 237454
rect 65330 236898 65566 237134
rect 96050 237218 96286 237454
rect 96050 236898 96286 237134
rect 126770 237218 127006 237454
rect 126770 236898 127006 237134
rect 157490 237218 157726 237454
rect 157490 236898 157726 237134
rect 188210 237218 188446 237454
rect 188210 236898 188446 237134
rect 218930 237218 219166 237454
rect 218930 236898 219166 237134
rect 249650 237218 249886 237454
rect 249650 236898 249886 237134
rect 280370 237218 280606 237454
rect 280370 236898 280606 237134
rect 311090 237218 311326 237454
rect 311090 236898 311326 237134
rect 341810 237218 342046 237454
rect 341810 236898 342046 237134
rect 372530 237218 372766 237454
rect 372530 236898 372766 237134
rect 403250 237218 403486 237454
rect 403250 236898 403486 237134
rect 433970 237218 434206 237454
rect 433970 236898 434206 237134
rect 464690 237218 464926 237454
rect 464690 236898 464926 237134
rect 495410 237218 495646 237454
rect 495410 236898 495646 237134
rect 526130 237218 526366 237454
rect 526130 236898 526366 237134
rect 19250 219218 19486 219454
rect 19250 218898 19486 219134
rect 49970 219218 50206 219454
rect 49970 218898 50206 219134
rect 80690 219218 80926 219454
rect 80690 218898 80926 219134
rect 111410 219218 111646 219454
rect 111410 218898 111646 219134
rect 142130 219218 142366 219454
rect 142130 218898 142366 219134
rect 172850 219218 173086 219454
rect 172850 218898 173086 219134
rect 203570 219218 203806 219454
rect 203570 218898 203806 219134
rect 234290 219218 234526 219454
rect 234290 218898 234526 219134
rect 265010 219218 265246 219454
rect 265010 218898 265246 219134
rect 295730 219218 295966 219454
rect 295730 218898 295966 219134
rect 326450 219218 326686 219454
rect 326450 218898 326686 219134
rect 357170 219218 357406 219454
rect 357170 218898 357406 219134
rect 387890 219218 388126 219454
rect 387890 218898 388126 219134
rect 418610 219218 418846 219454
rect 418610 218898 418846 219134
rect 449330 219218 449566 219454
rect 449330 218898 449566 219134
rect 480050 219218 480286 219454
rect 480050 218898 480286 219134
rect 510770 219218 511006 219454
rect 510770 218898 511006 219134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 34610 201218 34846 201454
rect 34610 200898 34846 201134
rect 65330 201218 65566 201454
rect 65330 200898 65566 201134
rect 96050 201218 96286 201454
rect 96050 200898 96286 201134
rect 126770 201218 127006 201454
rect 126770 200898 127006 201134
rect 157490 201218 157726 201454
rect 157490 200898 157726 201134
rect 188210 201218 188446 201454
rect 188210 200898 188446 201134
rect 218930 201218 219166 201454
rect 218930 200898 219166 201134
rect 249650 201218 249886 201454
rect 249650 200898 249886 201134
rect 280370 201218 280606 201454
rect 280370 200898 280606 201134
rect 311090 201218 311326 201454
rect 311090 200898 311326 201134
rect 341810 201218 342046 201454
rect 341810 200898 342046 201134
rect 372530 201218 372766 201454
rect 372530 200898 372766 201134
rect 403250 201218 403486 201454
rect 403250 200898 403486 201134
rect 433970 201218 434206 201454
rect 433970 200898 434206 201134
rect 464690 201218 464926 201454
rect 464690 200898 464926 201134
rect 495410 201218 495646 201454
rect 495410 200898 495646 201134
rect 526130 201218 526366 201454
rect 526130 200898 526366 201134
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 19250 183218 19486 183454
rect 19250 182898 19486 183134
rect 49970 183218 50206 183454
rect 49970 182898 50206 183134
rect 80690 183218 80926 183454
rect 80690 182898 80926 183134
rect 111410 183218 111646 183454
rect 111410 182898 111646 183134
rect 142130 183218 142366 183454
rect 142130 182898 142366 183134
rect 172850 183218 173086 183454
rect 172850 182898 173086 183134
rect 203570 183218 203806 183454
rect 203570 182898 203806 183134
rect 234290 183218 234526 183454
rect 234290 182898 234526 183134
rect 265010 183218 265246 183454
rect 265010 182898 265246 183134
rect 295730 183218 295966 183454
rect 295730 182898 295966 183134
rect 326450 183218 326686 183454
rect 326450 182898 326686 183134
rect 357170 183218 357406 183454
rect 357170 182898 357406 183134
rect 387890 183218 388126 183454
rect 387890 182898 388126 183134
rect 418610 183218 418846 183454
rect 418610 182898 418846 183134
rect 449330 183218 449566 183454
rect 449330 182898 449566 183134
rect 480050 183218 480286 183454
rect 480050 182898 480286 183134
rect 510770 183218 511006 183454
rect 510770 182898 511006 183134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 34610 165218 34846 165454
rect 34610 164898 34846 165134
rect 65330 165218 65566 165454
rect 65330 164898 65566 165134
rect 96050 165218 96286 165454
rect 96050 164898 96286 165134
rect 126770 165218 127006 165454
rect 126770 164898 127006 165134
rect 157490 165218 157726 165454
rect 157490 164898 157726 165134
rect 188210 165218 188446 165454
rect 188210 164898 188446 165134
rect 218930 165218 219166 165454
rect 218930 164898 219166 165134
rect 249650 165218 249886 165454
rect 249650 164898 249886 165134
rect 280370 165218 280606 165454
rect 280370 164898 280606 165134
rect 311090 165218 311326 165454
rect 311090 164898 311326 165134
rect 341810 165218 342046 165454
rect 341810 164898 342046 165134
rect 372530 165218 372766 165454
rect 372530 164898 372766 165134
rect 403250 165218 403486 165454
rect 403250 164898 403486 165134
rect 433970 165218 434206 165454
rect 433970 164898 434206 165134
rect 464690 165218 464926 165454
rect 464690 164898 464926 165134
rect 495410 165218 495646 165454
rect 495410 164898 495646 165134
rect 526130 165218 526366 165454
rect 526130 164898 526366 165134
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 19250 147218 19486 147454
rect 19250 146898 19486 147134
rect 49970 147218 50206 147454
rect 49970 146898 50206 147134
rect 80690 147218 80926 147454
rect 80690 146898 80926 147134
rect 111410 147218 111646 147454
rect 111410 146898 111646 147134
rect 142130 147218 142366 147454
rect 142130 146898 142366 147134
rect 172850 147218 173086 147454
rect 172850 146898 173086 147134
rect 203570 147218 203806 147454
rect 203570 146898 203806 147134
rect 234290 147218 234526 147454
rect 234290 146898 234526 147134
rect 265010 147218 265246 147454
rect 265010 146898 265246 147134
rect 295730 147218 295966 147454
rect 295730 146898 295966 147134
rect 326450 147218 326686 147454
rect 326450 146898 326686 147134
rect 357170 147218 357406 147454
rect 357170 146898 357406 147134
rect 387890 147218 388126 147454
rect 387890 146898 388126 147134
rect 418610 147218 418846 147454
rect 418610 146898 418846 147134
rect 449330 147218 449566 147454
rect 449330 146898 449566 147134
rect 480050 147218 480286 147454
rect 480050 146898 480286 147134
rect 510770 147218 511006 147454
rect 510770 146898 511006 147134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 34610 129218 34846 129454
rect 34610 128898 34846 129134
rect 65330 129218 65566 129454
rect 65330 128898 65566 129134
rect 96050 129218 96286 129454
rect 96050 128898 96286 129134
rect 126770 129218 127006 129454
rect 126770 128898 127006 129134
rect 157490 129218 157726 129454
rect 157490 128898 157726 129134
rect 188210 129218 188446 129454
rect 188210 128898 188446 129134
rect 218930 129218 219166 129454
rect 218930 128898 219166 129134
rect 249650 129218 249886 129454
rect 249650 128898 249886 129134
rect 280370 129218 280606 129454
rect 280370 128898 280606 129134
rect 311090 129218 311326 129454
rect 311090 128898 311326 129134
rect 341810 129218 342046 129454
rect 341810 128898 342046 129134
rect 372530 129218 372766 129454
rect 372530 128898 372766 129134
rect 403250 129218 403486 129454
rect 403250 128898 403486 129134
rect 433970 129218 434206 129454
rect 433970 128898 434206 129134
rect 464690 129218 464926 129454
rect 464690 128898 464926 129134
rect 495410 129218 495646 129454
rect 495410 128898 495646 129134
rect 526130 129218 526366 129454
rect 526130 128898 526366 129134
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 19250 111218 19486 111454
rect 19250 110898 19486 111134
rect 49970 111218 50206 111454
rect 49970 110898 50206 111134
rect 80690 111218 80926 111454
rect 80690 110898 80926 111134
rect 111410 111218 111646 111454
rect 111410 110898 111646 111134
rect 142130 111218 142366 111454
rect 142130 110898 142366 111134
rect 172850 111218 173086 111454
rect 172850 110898 173086 111134
rect 203570 111218 203806 111454
rect 203570 110898 203806 111134
rect 234290 111218 234526 111454
rect 234290 110898 234526 111134
rect 265010 111218 265246 111454
rect 265010 110898 265246 111134
rect 295730 111218 295966 111454
rect 295730 110898 295966 111134
rect 326450 111218 326686 111454
rect 326450 110898 326686 111134
rect 357170 111218 357406 111454
rect 357170 110898 357406 111134
rect 387890 111218 388126 111454
rect 387890 110898 388126 111134
rect 418610 111218 418846 111454
rect 418610 110898 418846 111134
rect 449330 111218 449566 111454
rect 449330 110898 449566 111134
rect 480050 111218 480286 111454
rect 480050 110898 480286 111134
rect 510770 111218 511006 111454
rect 510770 110898 511006 111134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 34610 93218 34846 93454
rect 34610 92898 34846 93134
rect 65330 93218 65566 93454
rect 65330 92898 65566 93134
rect 96050 93218 96286 93454
rect 96050 92898 96286 93134
rect 126770 93218 127006 93454
rect 126770 92898 127006 93134
rect 157490 93218 157726 93454
rect 157490 92898 157726 93134
rect 188210 93218 188446 93454
rect 188210 92898 188446 93134
rect 218930 93218 219166 93454
rect 218930 92898 219166 93134
rect 249650 93218 249886 93454
rect 249650 92898 249886 93134
rect 280370 93218 280606 93454
rect 280370 92898 280606 93134
rect 311090 93218 311326 93454
rect 311090 92898 311326 93134
rect 341810 93218 342046 93454
rect 341810 92898 342046 93134
rect 372530 93218 372766 93454
rect 372530 92898 372766 93134
rect 403250 93218 403486 93454
rect 403250 92898 403486 93134
rect 433970 93218 434206 93454
rect 433970 92898 434206 93134
rect 464690 93218 464926 93454
rect 464690 92898 464926 93134
rect 495410 93218 495646 93454
rect 495410 92898 495646 93134
rect 526130 93218 526366 93454
rect 526130 92898 526366 93134
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 19250 75218 19486 75454
rect 19250 74898 19486 75134
rect 49970 75218 50206 75454
rect 49970 74898 50206 75134
rect 80690 75218 80926 75454
rect 80690 74898 80926 75134
rect 111410 75218 111646 75454
rect 111410 74898 111646 75134
rect 142130 75218 142366 75454
rect 142130 74898 142366 75134
rect 172850 75218 173086 75454
rect 172850 74898 173086 75134
rect 203570 75218 203806 75454
rect 203570 74898 203806 75134
rect 234290 75218 234526 75454
rect 234290 74898 234526 75134
rect 265010 75218 265246 75454
rect 265010 74898 265246 75134
rect 295730 75218 295966 75454
rect 295730 74898 295966 75134
rect 326450 75218 326686 75454
rect 326450 74898 326686 75134
rect 357170 75218 357406 75454
rect 357170 74898 357406 75134
rect 387890 75218 388126 75454
rect 387890 74898 388126 75134
rect 418610 75218 418846 75454
rect 418610 74898 418846 75134
rect 449330 75218 449566 75454
rect 449330 74898 449566 75134
rect 480050 75218 480286 75454
rect 480050 74898 480286 75134
rect 510770 75218 511006 75454
rect 510770 74898 511006 75134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 34610 57218 34846 57454
rect 34610 56898 34846 57134
rect 65330 57218 65566 57454
rect 65330 56898 65566 57134
rect 96050 57218 96286 57454
rect 96050 56898 96286 57134
rect 126770 57218 127006 57454
rect 126770 56898 127006 57134
rect 157490 57218 157726 57454
rect 157490 56898 157726 57134
rect 188210 57218 188446 57454
rect 188210 56898 188446 57134
rect 218930 57218 219166 57454
rect 218930 56898 219166 57134
rect 249650 57218 249886 57454
rect 249650 56898 249886 57134
rect 280370 57218 280606 57454
rect 280370 56898 280606 57134
rect 311090 57218 311326 57454
rect 311090 56898 311326 57134
rect 341810 57218 342046 57454
rect 341810 56898 342046 57134
rect 372530 57218 372766 57454
rect 372530 56898 372766 57134
rect 403250 57218 403486 57454
rect 403250 56898 403486 57134
rect 433970 57218 434206 57454
rect 433970 56898 434206 57134
rect 464690 57218 464926 57454
rect 464690 56898 464926 57134
rect 495410 57218 495646 57454
rect 495410 56898 495646 57134
rect 526130 57218 526366 57454
rect 526130 56898 526366 57134
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 19250 39218 19486 39454
rect 19250 38898 19486 39134
rect 49970 39218 50206 39454
rect 49970 38898 50206 39134
rect 80690 39218 80926 39454
rect 80690 38898 80926 39134
rect 111410 39218 111646 39454
rect 111410 38898 111646 39134
rect 142130 39218 142366 39454
rect 142130 38898 142366 39134
rect 172850 39218 173086 39454
rect 172850 38898 173086 39134
rect 203570 39218 203806 39454
rect 203570 38898 203806 39134
rect 234290 39218 234526 39454
rect 234290 38898 234526 39134
rect 265010 39218 265246 39454
rect 265010 38898 265246 39134
rect 295730 39218 295966 39454
rect 295730 38898 295966 39134
rect 326450 39218 326686 39454
rect 326450 38898 326686 39134
rect 357170 39218 357406 39454
rect 357170 38898 357406 39134
rect 387890 39218 388126 39454
rect 387890 38898 388126 39134
rect 418610 39218 418846 39454
rect 418610 38898 418846 39134
rect 449330 39218 449566 39454
rect 449330 38898 449566 39134
rect 480050 39218 480286 39454
rect 480050 38898 480286 39134
rect 510770 39218 511006 39454
rect 510770 38898 511006 39134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 34610 21218 34846 21454
rect 34610 20898 34846 21134
rect 65330 21218 65566 21454
rect 65330 20898 65566 21134
rect 96050 21218 96286 21454
rect 96050 20898 96286 21134
rect 126770 21218 127006 21454
rect 126770 20898 127006 21134
rect 157490 21218 157726 21454
rect 157490 20898 157726 21134
rect 188210 21218 188446 21454
rect 188210 20898 188446 21134
rect 218930 21218 219166 21454
rect 218930 20898 219166 21134
rect 249650 21218 249886 21454
rect 249650 20898 249886 21134
rect 280370 21218 280606 21454
rect 280370 20898 280606 21134
rect 311090 21218 311326 21454
rect 311090 20898 311326 21134
rect 341810 21218 342046 21454
rect 341810 20898 342046 21134
rect 372530 21218 372766 21454
rect 372530 20898 372766 21134
rect 403250 21218 403486 21454
rect 403250 20898 403486 21134
rect 433970 21218 434206 21454
rect 433970 20898 434206 21134
rect 464690 21218 464926 21454
rect 464690 20898 464926 21134
rect 495410 21218 495646 21454
rect 495410 20898 495646 21134
rect 526130 21218 526366 21454
rect 526130 20898 526366 21134
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 19250 651454
rect 19486 651218 49970 651454
rect 50206 651218 80690 651454
rect 80926 651218 111410 651454
rect 111646 651218 142130 651454
rect 142366 651218 172850 651454
rect 173086 651218 203570 651454
rect 203806 651218 234290 651454
rect 234526 651218 265010 651454
rect 265246 651218 295730 651454
rect 295966 651218 326450 651454
rect 326686 651218 357170 651454
rect 357406 651218 387890 651454
rect 388126 651218 418610 651454
rect 418846 651218 449330 651454
rect 449566 651218 480050 651454
rect 480286 651218 510770 651454
rect 511006 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 19250 651134
rect 19486 650898 49970 651134
rect 50206 650898 80690 651134
rect 80926 650898 111410 651134
rect 111646 650898 142130 651134
rect 142366 650898 172850 651134
rect 173086 650898 203570 651134
rect 203806 650898 234290 651134
rect 234526 650898 265010 651134
rect 265246 650898 295730 651134
rect 295966 650898 326450 651134
rect 326686 650898 357170 651134
rect 357406 650898 387890 651134
rect 388126 650898 418610 651134
rect 418846 650898 449330 651134
rect 449566 650898 480050 651134
rect 480286 650898 510770 651134
rect 511006 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 34610 633454
rect 34846 633218 65330 633454
rect 65566 633218 96050 633454
rect 96286 633218 126770 633454
rect 127006 633218 157490 633454
rect 157726 633218 188210 633454
rect 188446 633218 218930 633454
rect 219166 633218 249650 633454
rect 249886 633218 280370 633454
rect 280606 633218 311090 633454
rect 311326 633218 341810 633454
rect 342046 633218 372530 633454
rect 372766 633218 403250 633454
rect 403486 633218 433970 633454
rect 434206 633218 464690 633454
rect 464926 633218 495410 633454
rect 495646 633218 526130 633454
rect 526366 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 34610 633134
rect 34846 632898 65330 633134
rect 65566 632898 96050 633134
rect 96286 632898 126770 633134
rect 127006 632898 157490 633134
rect 157726 632898 188210 633134
rect 188446 632898 218930 633134
rect 219166 632898 249650 633134
rect 249886 632898 280370 633134
rect 280606 632898 311090 633134
rect 311326 632898 341810 633134
rect 342046 632898 372530 633134
rect 372766 632898 403250 633134
rect 403486 632898 433970 633134
rect 434206 632898 464690 633134
rect 464926 632898 495410 633134
rect 495646 632898 526130 633134
rect 526366 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 19250 615454
rect 19486 615218 49970 615454
rect 50206 615218 80690 615454
rect 80926 615218 111410 615454
rect 111646 615218 142130 615454
rect 142366 615218 172850 615454
rect 173086 615218 203570 615454
rect 203806 615218 234290 615454
rect 234526 615218 265010 615454
rect 265246 615218 295730 615454
rect 295966 615218 326450 615454
rect 326686 615218 357170 615454
rect 357406 615218 387890 615454
rect 388126 615218 418610 615454
rect 418846 615218 449330 615454
rect 449566 615218 480050 615454
rect 480286 615218 510770 615454
rect 511006 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 19250 615134
rect 19486 614898 49970 615134
rect 50206 614898 80690 615134
rect 80926 614898 111410 615134
rect 111646 614898 142130 615134
rect 142366 614898 172850 615134
rect 173086 614898 203570 615134
rect 203806 614898 234290 615134
rect 234526 614898 265010 615134
rect 265246 614898 295730 615134
rect 295966 614898 326450 615134
rect 326686 614898 357170 615134
rect 357406 614898 387890 615134
rect 388126 614898 418610 615134
rect 418846 614898 449330 615134
rect 449566 614898 480050 615134
rect 480286 614898 510770 615134
rect 511006 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 34610 597454
rect 34846 597218 65330 597454
rect 65566 597218 96050 597454
rect 96286 597218 126770 597454
rect 127006 597218 157490 597454
rect 157726 597218 188210 597454
rect 188446 597218 218930 597454
rect 219166 597218 249650 597454
rect 249886 597218 280370 597454
rect 280606 597218 311090 597454
rect 311326 597218 341810 597454
rect 342046 597218 372530 597454
rect 372766 597218 403250 597454
rect 403486 597218 433970 597454
rect 434206 597218 464690 597454
rect 464926 597218 495410 597454
rect 495646 597218 526130 597454
rect 526366 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 34610 597134
rect 34846 596898 65330 597134
rect 65566 596898 96050 597134
rect 96286 596898 126770 597134
rect 127006 596898 157490 597134
rect 157726 596898 188210 597134
rect 188446 596898 218930 597134
rect 219166 596898 249650 597134
rect 249886 596898 280370 597134
rect 280606 596898 311090 597134
rect 311326 596898 341810 597134
rect 342046 596898 372530 597134
rect 372766 596898 403250 597134
rect 403486 596898 433970 597134
rect 434206 596898 464690 597134
rect 464926 596898 495410 597134
rect 495646 596898 526130 597134
rect 526366 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 19250 579454
rect 19486 579218 49970 579454
rect 50206 579218 80690 579454
rect 80926 579218 111410 579454
rect 111646 579218 142130 579454
rect 142366 579218 172850 579454
rect 173086 579218 203570 579454
rect 203806 579218 234290 579454
rect 234526 579218 265010 579454
rect 265246 579218 295730 579454
rect 295966 579218 326450 579454
rect 326686 579218 357170 579454
rect 357406 579218 387890 579454
rect 388126 579218 418610 579454
rect 418846 579218 449330 579454
rect 449566 579218 480050 579454
rect 480286 579218 510770 579454
rect 511006 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 19250 579134
rect 19486 578898 49970 579134
rect 50206 578898 80690 579134
rect 80926 578898 111410 579134
rect 111646 578898 142130 579134
rect 142366 578898 172850 579134
rect 173086 578898 203570 579134
rect 203806 578898 234290 579134
rect 234526 578898 265010 579134
rect 265246 578898 295730 579134
rect 295966 578898 326450 579134
rect 326686 578898 357170 579134
rect 357406 578898 387890 579134
rect 388126 578898 418610 579134
rect 418846 578898 449330 579134
rect 449566 578898 480050 579134
rect 480286 578898 510770 579134
rect 511006 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 34610 561454
rect 34846 561218 65330 561454
rect 65566 561218 96050 561454
rect 96286 561218 126770 561454
rect 127006 561218 157490 561454
rect 157726 561218 188210 561454
rect 188446 561218 218930 561454
rect 219166 561218 249650 561454
rect 249886 561218 280370 561454
rect 280606 561218 311090 561454
rect 311326 561218 341810 561454
rect 342046 561218 372530 561454
rect 372766 561218 403250 561454
rect 403486 561218 433970 561454
rect 434206 561218 464690 561454
rect 464926 561218 495410 561454
rect 495646 561218 526130 561454
rect 526366 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 34610 561134
rect 34846 560898 65330 561134
rect 65566 560898 96050 561134
rect 96286 560898 126770 561134
rect 127006 560898 157490 561134
rect 157726 560898 188210 561134
rect 188446 560898 218930 561134
rect 219166 560898 249650 561134
rect 249886 560898 280370 561134
rect 280606 560898 311090 561134
rect 311326 560898 341810 561134
rect 342046 560898 372530 561134
rect 372766 560898 403250 561134
rect 403486 560898 433970 561134
rect 434206 560898 464690 561134
rect 464926 560898 495410 561134
rect 495646 560898 526130 561134
rect 526366 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 19250 543454
rect 19486 543218 49970 543454
rect 50206 543218 80690 543454
rect 80926 543218 111410 543454
rect 111646 543218 142130 543454
rect 142366 543218 172850 543454
rect 173086 543218 203570 543454
rect 203806 543218 234290 543454
rect 234526 543218 265010 543454
rect 265246 543218 295730 543454
rect 295966 543218 326450 543454
rect 326686 543218 357170 543454
rect 357406 543218 387890 543454
rect 388126 543218 418610 543454
rect 418846 543218 449330 543454
rect 449566 543218 480050 543454
rect 480286 543218 510770 543454
rect 511006 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 19250 543134
rect 19486 542898 49970 543134
rect 50206 542898 80690 543134
rect 80926 542898 111410 543134
rect 111646 542898 142130 543134
rect 142366 542898 172850 543134
rect 173086 542898 203570 543134
rect 203806 542898 234290 543134
rect 234526 542898 265010 543134
rect 265246 542898 295730 543134
rect 295966 542898 326450 543134
rect 326686 542898 357170 543134
rect 357406 542898 387890 543134
rect 388126 542898 418610 543134
rect 418846 542898 449330 543134
rect 449566 542898 480050 543134
rect 480286 542898 510770 543134
rect 511006 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 34610 525454
rect 34846 525218 65330 525454
rect 65566 525218 96050 525454
rect 96286 525218 126770 525454
rect 127006 525218 157490 525454
rect 157726 525218 188210 525454
rect 188446 525218 218930 525454
rect 219166 525218 249650 525454
rect 249886 525218 280370 525454
rect 280606 525218 311090 525454
rect 311326 525218 341810 525454
rect 342046 525218 372530 525454
rect 372766 525218 403250 525454
rect 403486 525218 433970 525454
rect 434206 525218 464690 525454
rect 464926 525218 495410 525454
rect 495646 525218 526130 525454
rect 526366 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 34610 525134
rect 34846 524898 65330 525134
rect 65566 524898 96050 525134
rect 96286 524898 126770 525134
rect 127006 524898 157490 525134
rect 157726 524898 188210 525134
rect 188446 524898 218930 525134
rect 219166 524898 249650 525134
rect 249886 524898 280370 525134
rect 280606 524898 311090 525134
rect 311326 524898 341810 525134
rect 342046 524898 372530 525134
rect 372766 524898 403250 525134
rect 403486 524898 433970 525134
rect 434206 524898 464690 525134
rect 464926 524898 495410 525134
rect 495646 524898 526130 525134
rect 526366 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 19250 507454
rect 19486 507218 49970 507454
rect 50206 507218 80690 507454
rect 80926 507218 111410 507454
rect 111646 507218 142130 507454
rect 142366 507218 172850 507454
rect 173086 507218 203570 507454
rect 203806 507218 234290 507454
rect 234526 507218 265010 507454
rect 265246 507218 295730 507454
rect 295966 507218 326450 507454
rect 326686 507218 357170 507454
rect 357406 507218 387890 507454
rect 388126 507218 418610 507454
rect 418846 507218 449330 507454
rect 449566 507218 480050 507454
rect 480286 507218 510770 507454
rect 511006 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 19250 507134
rect 19486 506898 49970 507134
rect 50206 506898 80690 507134
rect 80926 506898 111410 507134
rect 111646 506898 142130 507134
rect 142366 506898 172850 507134
rect 173086 506898 203570 507134
rect 203806 506898 234290 507134
rect 234526 506898 265010 507134
rect 265246 506898 295730 507134
rect 295966 506898 326450 507134
rect 326686 506898 357170 507134
rect 357406 506898 387890 507134
rect 388126 506898 418610 507134
rect 418846 506898 449330 507134
rect 449566 506898 480050 507134
rect 480286 506898 510770 507134
rect 511006 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 34610 489454
rect 34846 489218 65330 489454
rect 65566 489218 96050 489454
rect 96286 489218 126770 489454
rect 127006 489218 157490 489454
rect 157726 489218 188210 489454
rect 188446 489218 218930 489454
rect 219166 489218 249650 489454
rect 249886 489218 280370 489454
rect 280606 489218 311090 489454
rect 311326 489218 341810 489454
rect 342046 489218 372530 489454
rect 372766 489218 403250 489454
rect 403486 489218 433970 489454
rect 434206 489218 464690 489454
rect 464926 489218 495410 489454
rect 495646 489218 526130 489454
rect 526366 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 34610 489134
rect 34846 488898 65330 489134
rect 65566 488898 96050 489134
rect 96286 488898 126770 489134
rect 127006 488898 157490 489134
rect 157726 488898 188210 489134
rect 188446 488898 218930 489134
rect 219166 488898 249650 489134
rect 249886 488898 280370 489134
rect 280606 488898 311090 489134
rect 311326 488898 341810 489134
rect 342046 488898 372530 489134
rect 372766 488898 403250 489134
rect 403486 488898 433970 489134
rect 434206 488898 464690 489134
rect 464926 488898 495410 489134
rect 495646 488898 526130 489134
rect 526366 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 19250 471454
rect 19486 471218 49970 471454
rect 50206 471218 80690 471454
rect 80926 471218 111410 471454
rect 111646 471218 142130 471454
rect 142366 471218 172850 471454
rect 173086 471218 203570 471454
rect 203806 471218 234290 471454
rect 234526 471218 265010 471454
rect 265246 471218 295730 471454
rect 295966 471218 326450 471454
rect 326686 471218 357170 471454
rect 357406 471218 387890 471454
rect 388126 471218 418610 471454
rect 418846 471218 449330 471454
rect 449566 471218 480050 471454
rect 480286 471218 510770 471454
rect 511006 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 19250 471134
rect 19486 470898 49970 471134
rect 50206 470898 80690 471134
rect 80926 470898 111410 471134
rect 111646 470898 142130 471134
rect 142366 470898 172850 471134
rect 173086 470898 203570 471134
rect 203806 470898 234290 471134
rect 234526 470898 265010 471134
rect 265246 470898 295730 471134
rect 295966 470898 326450 471134
rect 326686 470898 357170 471134
rect 357406 470898 387890 471134
rect 388126 470898 418610 471134
rect 418846 470898 449330 471134
rect 449566 470898 480050 471134
rect 480286 470898 510770 471134
rect 511006 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 34610 453454
rect 34846 453218 65330 453454
rect 65566 453218 96050 453454
rect 96286 453218 126770 453454
rect 127006 453218 157490 453454
rect 157726 453218 188210 453454
rect 188446 453218 218930 453454
rect 219166 453218 249650 453454
rect 249886 453218 280370 453454
rect 280606 453218 311090 453454
rect 311326 453218 341810 453454
rect 342046 453218 372530 453454
rect 372766 453218 403250 453454
rect 403486 453218 433970 453454
rect 434206 453218 464690 453454
rect 464926 453218 495410 453454
rect 495646 453218 526130 453454
rect 526366 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 34610 453134
rect 34846 452898 65330 453134
rect 65566 452898 96050 453134
rect 96286 452898 126770 453134
rect 127006 452898 157490 453134
rect 157726 452898 188210 453134
rect 188446 452898 218930 453134
rect 219166 452898 249650 453134
rect 249886 452898 280370 453134
rect 280606 452898 311090 453134
rect 311326 452898 341810 453134
rect 342046 452898 372530 453134
rect 372766 452898 403250 453134
rect 403486 452898 433970 453134
rect 434206 452898 464690 453134
rect 464926 452898 495410 453134
rect 495646 452898 526130 453134
rect 526366 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 19250 435454
rect 19486 435218 49970 435454
rect 50206 435218 80690 435454
rect 80926 435218 111410 435454
rect 111646 435218 142130 435454
rect 142366 435218 172850 435454
rect 173086 435218 203570 435454
rect 203806 435218 234290 435454
rect 234526 435218 265010 435454
rect 265246 435218 295730 435454
rect 295966 435218 326450 435454
rect 326686 435218 357170 435454
rect 357406 435218 387890 435454
rect 388126 435218 418610 435454
rect 418846 435218 449330 435454
rect 449566 435218 480050 435454
rect 480286 435218 510770 435454
rect 511006 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 19250 435134
rect 19486 434898 49970 435134
rect 50206 434898 80690 435134
rect 80926 434898 111410 435134
rect 111646 434898 142130 435134
rect 142366 434898 172850 435134
rect 173086 434898 203570 435134
rect 203806 434898 234290 435134
rect 234526 434898 265010 435134
rect 265246 434898 295730 435134
rect 295966 434898 326450 435134
rect 326686 434898 357170 435134
rect 357406 434898 387890 435134
rect 388126 434898 418610 435134
rect 418846 434898 449330 435134
rect 449566 434898 480050 435134
rect 480286 434898 510770 435134
rect 511006 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 34610 417454
rect 34846 417218 65330 417454
rect 65566 417218 96050 417454
rect 96286 417218 126770 417454
rect 127006 417218 157490 417454
rect 157726 417218 188210 417454
rect 188446 417218 218930 417454
rect 219166 417218 249650 417454
rect 249886 417218 280370 417454
rect 280606 417218 311090 417454
rect 311326 417218 341810 417454
rect 342046 417218 372530 417454
rect 372766 417218 403250 417454
rect 403486 417218 433970 417454
rect 434206 417218 464690 417454
rect 464926 417218 495410 417454
rect 495646 417218 526130 417454
rect 526366 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 34610 417134
rect 34846 416898 65330 417134
rect 65566 416898 96050 417134
rect 96286 416898 126770 417134
rect 127006 416898 157490 417134
rect 157726 416898 188210 417134
rect 188446 416898 218930 417134
rect 219166 416898 249650 417134
rect 249886 416898 280370 417134
rect 280606 416898 311090 417134
rect 311326 416898 341810 417134
rect 342046 416898 372530 417134
rect 372766 416898 403250 417134
rect 403486 416898 433970 417134
rect 434206 416898 464690 417134
rect 464926 416898 495410 417134
rect 495646 416898 526130 417134
rect 526366 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 19250 399454
rect 19486 399218 49970 399454
rect 50206 399218 80690 399454
rect 80926 399218 111410 399454
rect 111646 399218 142130 399454
rect 142366 399218 172850 399454
rect 173086 399218 203570 399454
rect 203806 399218 234290 399454
rect 234526 399218 265010 399454
rect 265246 399218 295730 399454
rect 295966 399218 326450 399454
rect 326686 399218 357170 399454
rect 357406 399218 387890 399454
rect 388126 399218 418610 399454
rect 418846 399218 449330 399454
rect 449566 399218 480050 399454
rect 480286 399218 510770 399454
rect 511006 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 19250 399134
rect 19486 398898 49970 399134
rect 50206 398898 80690 399134
rect 80926 398898 111410 399134
rect 111646 398898 142130 399134
rect 142366 398898 172850 399134
rect 173086 398898 203570 399134
rect 203806 398898 234290 399134
rect 234526 398898 265010 399134
rect 265246 398898 295730 399134
rect 295966 398898 326450 399134
rect 326686 398898 357170 399134
rect 357406 398898 387890 399134
rect 388126 398898 418610 399134
rect 418846 398898 449330 399134
rect 449566 398898 480050 399134
rect 480286 398898 510770 399134
rect 511006 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 34610 381454
rect 34846 381218 65330 381454
rect 65566 381218 96050 381454
rect 96286 381218 126770 381454
rect 127006 381218 157490 381454
rect 157726 381218 188210 381454
rect 188446 381218 218930 381454
rect 219166 381218 249650 381454
rect 249886 381218 280370 381454
rect 280606 381218 311090 381454
rect 311326 381218 341810 381454
rect 342046 381218 372530 381454
rect 372766 381218 403250 381454
rect 403486 381218 433970 381454
rect 434206 381218 464690 381454
rect 464926 381218 495410 381454
rect 495646 381218 526130 381454
rect 526366 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 34610 381134
rect 34846 380898 65330 381134
rect 65566 380898 96050 381134
rect 96286 380898 126770 381134
rect 127006 380898 157490 381134
rect 157726 380898 188210 381134
rect 188446 380898 218930 381134
rect 219166 380898 249650 381134
rect 249886 380898 280370 381134
rect 280606 380898 311090 381134
rect 311326 380898 341810 381134
rect 342046 380898 372530 381134
rect 372766 380898 403250 381134
rect 403486 380898 433970 381134
rect 434206 380898 464690 381134
rect 464926 380898 495410 381134
rect 495646 380898 526130 381134
rect 526366 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 19250 363454
rect 19486 363218 49970 363454
rect 50206 363218 80690 363454
rect 80926 363218 111410 363454
rect 111646 363218 142130 363454
rect 142366 363218 172850 363454
rect 173086 363218 203570 363454
rect 203806 363218 234290 363454
rect 234526 363218 265010 363454
rect 265246 363218 295730 363454
rect 295966 363218 326450 363454
rect 326686 363218 357170 363454
rect 357406 363218 387890 363454
rect 388126 363218 418610 363454
rect 418846 363218 449330 363454
rect 449566 363218 480050 363454
rect 480286 363218 510770 363454
rect 511006 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 19250 363134
rect 19486 362898 49970 363134
rect 50206 362898 80690 363134
rect 80926 362898 111410 363134
rect 111646 362898 142130 363134
rect 142366 362898 172850 363134
rect 173086 362898 203570 363134
rect 203806 362898 234290 363134
rect 234526 362898 265010 363134
rect 265246 362898 295730 363134
rect 295966 362898 326450 363134
rect 326686 362898 357170 363134
rect 357406 362898 387890 363134
rect 388126 362898 418610 363134
rect 418846 362898 449330 363134
rect 449566 362898 480050 363134
rect 480286 362898 510770 363134
rect 511006 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 34610 345454
rect 34846 345218 65330 345454
rect 65566 345218 96050 345454
rect 96286 345218 126770 345454
rect 127006 345218 157490 345454
rect 157726 345218 188210 345454
rect 188446 345218 218930 345454
rect 219166 345218 249650 345454
rect 249886 345218 280370 345454
rect 280606 345218 311090 345454
rect 311326 345218 341810 345454
rect 342046 345218 372530 345454
rect 372766 345218 403250 345454
rect 403486 345218 433970 345454
rect 434206 345218 464690 345454
rect 464926 345218 495410 345454
rect 495646 345218 526130 345454
rect 526366 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 34610 345134
rect 34846 344898 65330 345134
rect 65566 344898 96050 345134
rect 96286 344898 126770 345134
rect 127006 344898 157490 345134
rect 157726 344898 188210 345134
rect 188446 344898 218930 345134
rect 219166 344898 249650 345134
rect 249886 344898 280370 345134
rect 280606 344898 311090 345134
rect 311326 344898 341810 345134
rect 342046 344898 372530 345134
rect 372766 344898 403250 345134
rect 403486 344898 433970 345134
rect 434206 344898 464690 345134
rect 464926 344898 495410 345134
rect 495646 344898 526130 345134
rect 526366 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 19250 327454
rect 19486 327218 49970 327454
rect 50206 327218 80690 327454
rect 80926 327218 111410 327454
rect 111646 327218 142130 327454
rect 142366 327218 172850 327454
rect 173086 327218 203570 327454
rect 203806 327218 234290 327454
rect 234526 327218 265010 327454
rect 265246 327218 295730 327454
rect 295966 327218 326450 327454
rect 326686 327218 357170 327454
rect 357406 327218 387890 327454
rect 388126 327218 418610 327454
rect 418846 327218 449330 327454
rect 449566 327218 480050 327454
rect 480286 327218 510770 327454
rect 511006 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 19250 327134
rect 19486 326898 49970 327134
rect 50206 326898 80690 327134
rect 80926 326898 111410 327134
rect 111646 326898 142130 327134
rect 142366 326898 172850 327134
rect 173086 326898 203570 327134
rect 203806 326898 234290 327134
rect 234526 326898 265010 327134
rect 265246 326898 295730 327134
rect 295966 326898 326450 327134
rect 326686 326898 357170 327134
rect 357406 326898 387890 327134
rect 388126 326898 418610 327134
rect 418846 326898 449330 327134
rect 449566 326898 480050 327134
rect 480286 326898 510770 327134
rect 511006 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 34610 309454
rect 34846 309218 65330 309454
rect 65566 309218 96050 309454
rect 96286 309218 126770 309454
rect 127006 309218 157490 309454
rect 157726 309218 188210 309454
rect 188446 309218 218930 309454
rect 219166 309218 249650 309454
rect 249886 309218 280370 309454
rect 280606 309218 311090 309454
rect 311326 309218 341810 309454
rect 342046 309218 372530 309454
rect 372766 309218 403250 309454
rect 403486 309218 433970 309454
rect 434206 309218 464690 309454
rect 464926 309218 495410 309454
rect 495646 309218 526130 309454
rect 526366 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 34610 309134
rect 34846 308898 65330 309134
rect 65566 308898 96050 309134
rect 96286 308898 126770 309134
rect 127006 308898 157490 309134
rect 157726 308898 188210 309134
rect 188446 308898 218930 309134
rect 219166 308898 249650 309134
rect 249886 308898 280370 309134
rect 280606 308898 311090 309134
rect 311326 308898 341810 309134
rect 342046 308898 372530 309134
rect 372766 308898 403250 309134
rect 403486 308898 433970 309134
rect 434206 308898 464690 309134
rect 464926 308898 495410 309134
rect 495646 308898 526130 309134
rect 526366 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 19250 291454
rect 19486 291218 49970 291454
rect 50206 291218 80690 291454
rect 80926 291218 111410 291454
rect 111646 291218 142130 291454
rect 142366 291218 172850 291454
rect 173086 291218 203570 291454
rect 203806 291218 234290 291454
rect 234526 291218 265010 291454
rect 265246 291218 295730 291454
rect 295966 291218 326450 291454
rect 326686 291218 357170 291454
rect 357406 291218 387890 291454
rect 388126 291218 418610 291454
rect 418846 291218 449330 291454
rect 449566 291218 480050 291454
rect 480286 291218 510770 291454
rect 511006 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 19250 291134
rect 19486 290898 49970 291134
rect 50206 290898 80690 291134
rect 80926 290898 111410 291134
rect 111646 290898 142130 291134
rect 142366 290898 172850 291134
rect 173086 290898 203570 291134
rect 203806 290898 234290 291134
rect 234526 290898 265010 291134
rect 265246 290898 295730 291134
rect 295966 290898 326450 291134
rect 326686 290898 357170 291134
rect 357406 290898 387890 291134
rect 388126 290898 418610 291134
rect 418846 290898 449330 291134
rect 449566 290898 480050 291134
rect 480286 290898 510770 291134
rect 511006 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 34610 273454
rect 34846 273218 65330 273454
rect 65566 273218 96050 273454
rect 96286 273218 126770 273454
rect 127006 273218 157490 273454
rect 157726 273218 188210 273454
rect 188446 273218 218930 273454
rect 219166 273218 249650 273454
rect 249886 273218 280370 273454
rect 280606 273218 311090 273454
rect 311326 273218 341810 273454
rect 342046 273218 372530 273454
rect 372766 273218 403250 273454
rect 403486 273218 433970 273454
rect 434206 273218 464690 273454
rect 464926 273218 495410 273454
rect 495646 273218 526130 273454
rect 526366 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 34610 273134
rect 34846 272898 65330 273134
rect 65566 272898 96050 273134
rect 96286 272898 126770 273134
rect 127006 272898 157490 273134
rect 157726 272898 188210 273134
rect 188446 272898 218930 273134
rect 219166 272898 249650 273134
rect 249886 272898 280370 273134
rect 280606 272898 311090 273134
rect 311326 272898 341810 273134
rect 342046 272898 372530 273134
rect 372766 272898 403250 273134
rect 403486 272898 433970 273134
rect 434206 272898 464690 273134
rect 464926 272898 495410 273134
rect 495646 272898 526130 273134
rect 526366 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 19250 255454
rect 19486 255218 49970 255454
rect 50206 255218 80690 255454
rect 80926 255218 111410 255454
rect 111646 255218 142130 255454
rect 142366 255218 172850 255454
rect 173086 255218 203570 255454
rect 203806 255218 234290 255454
rect 234526 255218 265010 255454
rect 265246 255218 295730 255454
rect 295966 255218 326450 255454
rect 326686 255218 357170 255454
rect 357406 255218 387890 255454
rect 388126 255218 418610 255454
rect 418846 255218 449330 255454
rect 449566 255218 480050 255454
rect 480286 255218 510770 255454
rect 511006 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 19250 255134
rect 19486 254898 49970 255134
rect 50206 254898 80690 255134
rect 80926 254898 111410 255134
rect 111646 254898 142130 255134
rect 142366 254898 172850 255134
rect 173086 254898 203570 255134
rect 203806 254898 234290 255134
rect 234526 254898 265010 255134
rect 265246 254898 295730 255134
rect 295966 254898 326450 255134
rect 326686 254898 357170 255134
rect 357406 254898 387890 255134
rect 388126 254898 418610 255134
rect 418846 254898 449330 255134
rect 449566 254898 480050 255134
rect 480286 254898 510770 255134
rect 511006 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 34610 237454
rect 34846 237218 65330 237454
rect 65566 237218 96050 237454
rect 96286 237218 126770 237454
rect 127006 237218 157490 237454
rect 157726 237218 188210 237454
rect 188446 237218 218930 237454
rect 219166 237218 249650 237454
rect 249886 237218 280370 237454
rect 280606 237218 311090 237454
rect 311326 237218 341810 237454
rect 342046 237218 372530 237454
rect 372766 237218 403250 237454
rect 403486 237218 433970 237454
rect 434206 237218 464690 237454
rect 464926 237218 495410 237454
rect 495646 237218 526130 237454
rect 526366 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 34610 237134
rect 34846 236898 65330 237134
rect 65566 236898 96050 237134
rect 96286 236898 126770 237134
rect 127006 236898 157490 237134
rect 157726 236898 188210 237134
rect 188446 236898 218930 237134
rect 219166 236898 249650 237134
rect 249886 236898 280370 237134
rect 280606 236898 311090 237134
rect 311326 236898 341810 237134
rect 342046 236898 372530 237134
rect 372766 236898 403250 237134
rect 403486 236898 433970 237134
rect 434206 236898 464690 237134
rect 464926 236898 495410 237134
rect 495646 236898 526130 237134
rect 526366 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 19250 219454
rect 19486 219218 49970 219454
rect 50206 219218 80690 219454
rect 80926 219218 111410 219454
rect 111646 219218 142130 219454
rect 142366 219218 172850 219454
rect 173086 219218 203570 219454
rect 203806 219218 234290 219454
rect 234526 219218 265010 219454
rect 265246 219218 295730 219454
rect 295966 219218 326450 219454
rect 326686 219218 357170 219454
rect 357406 219218 387890 219454
rect 388126 219218 418610 219454
rect 418846 219218 449330 219454
rect 449566 219218 480050 219454
rect 480286 219218 510770 219454
rect 511006 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 19250 219134
rect 19486 218898 49970 219134
rect 50206 218898 80690 219134
rect 80926 218898 111410 219134
rect 111646 218898 142130 219134
rect 142366 218898 172850 219134
rect 173086 218898 203570 219134
rect 203806 218898 234290 219134
rect 234526 218898 265010 219134
rect 265246 218898 295730 219134
rect 295966 218898 326450 219134
rect 326686 218898 357170 219134
rect 357406 218898 387890 219134
rect 388126 218898 418610 219134
rect 418846 218898 449330 219134
rect 449566 218898 480050 219134
rect 480286 218898 510770 219134
rect 511006 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 34610 201454
rect 34846 201218 65330 201454
rect 65566 201218 96050 201454
rect 96286 201218 126770 201454
rect 127006 201218 157490 201454
rect 157726 201218 188210 201454
rect 188446 201218 218930 201454
rect 219166 201218 249650 201454
rect 249886 201218 280370 201454
rect 280606 201218 311090 201454
rect 311326 201218 341810 201454
rect 342046 201218 372530 201454
rect 372766 201218 403250 201454
rect 403486 201218 433970 201454
rect 434206 201218 464690 201454
rect 464926 201218 495410 201454
rect 495646 201218 526130 201454
rect 526366 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 34610 201134
rect 34846 200898 65330 201134
rect 65566 200898 96050 201134
rect 96286 200898 126770 201134
rect 127006 200898 157490 201134
rect 157726 200898 188210 201134
rect 188446 200898 218930 201134
rect 219166 200898 249650 201134
rect 249886 200898 280370 201134
rect 280606 200898 311090 201134
rect 311326 200898 341810 201134
rect 342046 200898 372530 201134
rect 372766 200898 403250 201134
rect 403486 200898 433970 201134
rect 434206 200898 464690 201134
rect 464926 200898 495410 201134
rect 495646 200898 526130 201134
rect 526366 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 19250 183454
rect 19486 183218 49970 183454
rect 50206 183218 80690 183454
rect 80926 183218 111410 183454
rect 111646 183218 142130 183454
rect 142366 183218 172850 183454
rect 173086 183218 203570 183454
rect 203806 183218 234290 183454
rect 234526 183218 265010 183454
rect 265246 183218 295730 183454
rect 295966 183218 326450 183454
rect 326686 183218 357170 183454
rect 357406 183218 387890 183454
rect 388126 183218 418610 183454
rect 418846 183218 449330 183454
rect 449566 183218 480050 183454
rect 480286 183218 510770 183454
rect 511006 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 19250 183134
rect 19486 182898 49970 183134
rect 50206 182898 80690 183134
rect 80926 182898 111410 183134
rect 111646 182898 142130 183134
rect 142366 182898 172850 183134
rect 173086 182898 203570 183134
rect 203806 182898 234290 183134
rect 234526 182898 265010 183134
rect 265246 182898 295730 183134
rect 295966 182898 326450 183134
rect 326686 182898 357170 183134
rect 357406 182898 387890 183134
rect 388126 182898 418610 183134
rect 418846 182898 449330 183134
rect 449566 182898 480050 183134
rect 480286 182898 510770 183134
rect 511006 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 34610 165454
rect 34846 165218 65330 165454
rect 65566 165218 96050 165454
rect 96286 165218 126770 165454
rect 127006 165218 157490 165454
rect 157726 165218 188210 165454
rect 188446 165218 218930 165454
rect 219166 165218 249650 165454
rect 249886 165218 280370 165454
rect 280606 165218 311090 165454
rect 311326 165218 341810 165454
rect 342046 165218 372530 165454
rect 372766 165218 403250 165454
rect 403486 165218 433970 165454
rect 434206 165218 464690 165454
rect 464926 165218 495410 165454
rect 495646 165218 526130 165454
rect 526366 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 34610 165134
rect 34846 164898 65330 165134
rect 65566 164898 96050 165134
rect 96286 164898 126770 165134
rect 127006 164898 157490 165134
rect 157726 164898 188210 165134
rect 188446 164898 218930 165134
rect 219166 164898 249650 165134
rect 249886 164898 280370 165134
rect 280606 164898 311090 165134
rect 311326 164898 341810 165134
rect 342046 164898 372530 165134
rect 372766 164898 403250 165134
rect 403486 164898 433970 165134
rect 434206 164898 464690 165134
rect 464926 164898 495410 165134
rect 495646 164898 526130 165134
rect 526366 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 19250 147454
rect 19486 147218 49970 147454
rect 50206 147218 80690 147454
rect 80926 147218 111410 147454
rect 111646 147218 142130 147454
rect 142366 147218 172850 147454
rect 173086 147218 203570 147454
rect 203806 147218 234290 147454
rect 234526 147218 265010 147454
rect 265246 147218 295730 147454
rect 295966 147218 326450 147454
rect 326686 147218 357170 147454
rect 357406 147218 387890 147454
rect 388126 147218 418610 147454
rect 418846 147218 449330 147454
rect 449566 147218 480050 147454
rect 480286 147218 510770 147454
rect 511006 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 19250 147134
rect 19486 146898 49970 147134
rect 50206 146898 80690 147134
rect 80926 146898 111410 147134
rect 111646 146898 142130 147134
rect 142366 146898 172850 147134
rect 173086 146898 203570 147134
rect 203806 146898 234290 147134
rect 234526 146898 265010 147134
rect 265246 146898 295730 147134
rect 295966 146898 326450 147134
rect 326686 146898 357170 147134
rect 357406 146898 387890 147134
rect 388126 146898 418610 147134
rect 418846 146898 449330 147134
rect 449566 146898 480050 147134
rect 480286 146898 510770 147134
rect 511006 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 34610 129454
rect 34846 129218 65330 129454
rect 65566 129218 96050 129454
rect 96286 129218 126770 129454
rect 127006 129218 157490 129454
rect 157726 129218 188210 129454
rect 188446 129218 218930 129454
rect 219166 129218 249650 129454
rect 249886 129218 280370 129454
rect 280606 129218 311090 129454
rect 311326 129218 341810 129454
rect 342046 129218 372530 129454
rect 372766 129218 403250 129454
rect 403486 129218 433970 129454
rect 434206 129218 464690 129454
rect 464926 129218 495410 129454
rect 495646 129218 526130 129454
rect 526366 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 34610 129134
rect 34846 128898 65330 129134
rect 65566 128898 96050 129134
rect 96286 128898 126770 129134
rect 127006 128898 157490 129134
rect 157726 128898 188210 129134
rect 188446 128898 218930 129134
rect 219166 128898 249650 129134
rect 249886 128898 280370 129134
rect 280606 128898 311090 129134
rect 311326 128898 341810 129134
rect 342046 128898 372530 129134
rect 372766 128898 403250 129134
rect 403486 128898 433970 129134
rect 434206 128898 464690 129134
rect 464926 128898 495410 129134
rect 495646 128898 526130 129134
rect 526366 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 19250 111454
rect 19486 111218 49970 111454
rect 50206 111218 80690 111454
rect 80926 111218 111410 111454
rect 111646 111218 142130 111454
rect 142366 111218 172850 111454
rect 173086 111218 203570 111454
rect 203806 111218 234290 111454
rect 234526 111218 265010 111454
rect 265246 111218 295730 111454
rect 295966 111218 326450 111454
rect 326686 111218 357170 111454
rect 357406 111218 387890 111454
rect 388126 111218 418610 111454
rect 418846 111218 449330 111454
rect 449566 111218 480050 111454
rect 480286 111218 510770 111454
rect 511006 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 19250 111134
rect 19486 110898 49970 111134
rect 50206 110898 80690 111134
rect 80926 110898 111410 111134
rect 111646 110898 142130 111134
rect 142366 110898 172850 111134
rect 173086 110898 203570 111134
rect 203806 110898 234290 111134
rect 234526 110898 265010 111134
rect 265246 110898 295730 111134
rect 295966 110898 326450 111134
rect 326686 110898 357170 111134
rect 357406 110898 387890 111134
rect 388126 110898 418610 111134
rect 418846 110898 449330 111134
rect 449566 110898 480050 111134
rect 480286 110898 510770 111134
rect 511006 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 34610 93454
rect 34846 93218 65330 93454
rect 65566 93218 96050 93454
rect 96286 93218 126770 93454
rect 127006 93218 157490 93454
rect 157726 93218 188210 93454
rect 188446 93218 218930 93454
rect 219166 93218 249650 93454
rect 249886 93218 280370 93454
rect 280606 93218 311090 93454
rect 311326 93218 341810 93454
rect 342046 93218 372530 93454
rect 372766 93218 403250 93454
rect 403486 93218 433970 93454
rect 434206 93218 464690 93454
rect 464926 93218 495410 93454
rect 495646 93218 526130 93454
rect 526366 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 34610 93134
rect 34846 92898 65330 93134
rect 65566 92898 96050 93134
rect 96286 92898 126770 93134
rect 127006 92898 157490 93134
rect 157726 92898 188210 93134
rect 188446 92898 218930 93134
rect 219166 92898 249650 93134
rect 249886 92898 280370 93134
rect 280606 92898 311090 93134
rect 311326 92898 341810 93134
rect 342046 92898 372530 93134
rect 372766 92898 403250 93134
rect 403486 92898 433970 93134
rect 434206 92898 464690 93134
rect 464926 92898 495410 93134
rect 495646 92898 526130 93134
rect 526366 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 19250 75454
rect 19486 75218 49970 75454
rect 50206 75218 80690 75454
rect 80926 75218 111410 75454
rect 111646 75218 142130 75454
rect 142366 75218 172850 75454
rect 173086 75218 203570 75454
rect 203806 75218 234290 75454
rect 234526 75218 265010 75454
rect 265246 75218 295730 75454
rect 295966 75218 326450 75454
rect 326686 75218 357170 75454
rect 357406 75218 387890 75454
rect 388126 75218 418610 75454
rect 418846 75218 449330 75454
rect 449566 75218 480050 75454
rect 480286 75218 510770 75454
rect 511006 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 19250 75134
rect 19486 74898 49970 75134
rect 50206 74898 80690 75134
rect 80926 74898 111410 75134
rect 111646 74898 142130 75134
rect 142366 74898 172850 75134
rect 173086 74898 203570 75134
rect 203806 74898 234290 75134
rect 234526 74898 265010 75134
rect 265246 74898 295730 75134
rect 295966 74898 326450 75134
rect 326686 74898 357170 75134
rect 357406 74898 387890 75134
rect 388126 74898 418610 75134
rect 418846 74898 449330 75134
rect 449566 74898 480050 75134
rect 480286 74898 510770 75134
rect 511006 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 34610 57454
rect 34846 57218 65330 57454
rect 65566 57218 96050 57454
rect 96286 57218 126770 57454
rect 127006 57218 157490 57454
rect 157726 57218 188210 57454
rect 188446 57218 218930 57454
rect 219166 57218 249650 57454
rect 249886 57218 280370 57454
rect 280606 57218 311090 57454
rect 311326 57218 341810 57454
rect 342046 57218 372530 57454
rect 372766 57218 403250 57454
rect 403486 57218 433970 57454
rect 434206 57218 464690 57454
rect 464926 57218 495410 57454
rect 495646 57218 526130 57454
rect 526366 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 34610 57134
rect 34846 56898 65330 57134
rect 65566 56898 96050 57134
rect 96286 56898 126770 57134
rect 127006 56898 157490 57134
rect 157726 56898 188210 57134
rect 188446 56898 218930 57134
rect 219166 56898 249650 57134
rect 249886 56898 280370 57134
rect 280606 56898 311090 57134
rect 311326 56898 341810 57134
rect 342046 56898 372530 57134
rect 372766 56898 403250 57134
rect 403486 56898 433970 57134
rect 434206 56898 464690 57134
rect 464926 56898 495410 57134
rect 495646 56898 526130 57134
rect 526366 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 19250 39454
rect 19486 39218 49970 39454
rect 50206 39218 80690 39454
rect 80926 39218 111410 39454
rect 111646 39218 142130 39454
rect 142366 39218 172850 39454
rect 173086 39218 203570 39454
rect 203806 39218 234290 39454
rect 234526 39218 265010 39454
rect 265246 39218 295730 39454
rect 295966 39218 326450 39454
rect 326686 39218 357170 39454
rect 357406 39218 387890 39454
rect 388126 39218 418610 39454
rect 418846 39218 449330 39454
rect 449566 39218 480050 39454
rect 480286 39218 510770 39454
rect 511006 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 19250 39134
rect 19486 38898 49970 39134
rect 50206 38898 80690 39134
rect 80926 38898 111410 39134
rect 111646 38898 142130 39134
rect 142366 38898 172850 39134
rect 173086 38898 203570 39134
rect 203806 38898 234290 39134
rect 234526 38898 265010 39134
rect 265246 38898 295730 39134
rect 295966 38898 326450 39134
rect 326686 38898 357170 39134
rect 357406 38898 387890 39134
rect 388126 38898 418610 39134
rect 418846 38898 449330 39134
rect 449566 38898 480050 39134
rect 480286 38898 510770 39134
rect 511006 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 34610 21454
rect 34846 21218 65330 21454
rect 65566 21218 96050 21454
rect 96286 21218 126770 21454
rect 127006 21218 157490 21454
rect 157726 21218 188210 21454
rect 188446 21218 218930 21454
rect 219166 21218 249650 21454
rect 249886 21218 280370 21454
rect 280606 21218 311090 21454
rect 311326 21218 341810 21454
rect 342046 21218 372530 21454
rect 372766 21218 403250 21454
rect 403486 21218 433970 21454
rect 434206 21218 464690 21454
rect 464926 21218 495410 21454
rect 495646 21218 526130 21454
rect 526366 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 34610 21134
rect 34846 20898 65330 21134
rect 65566 20898 96050 21134
rect 96286 20898 126770 21134
rect 127006 20898 157490 21134
rect 157726 20898 188210 21134
rect 188446 20898 218930 21134
rect 219166 20898 249650 21134
rect 249886 20898 280370 21134
rect 280606 20898 311090 21134
rect 311326 20898 341810 21134
rect 342046 20898 372530 21134
rect 372766 20898 403250 21134
rect 403486 20898 433970 21134
rect 434206 20898 464690 21134
rect 464926 20898 495410 21134
rect 495646 20898 526130 21134
rect 526366 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use top  dut
timestamp 0
transform 1 0 15000 0 1 15000
box 0 0 520000 640000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 13000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 657000 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 657000 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 657000 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 657000 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 657000 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 657000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 657000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 657000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 657000 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 657000 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 657000 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 657000 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 657000 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 657000 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 13000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 657000 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 657000 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 657000 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 657000 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 657000 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 657000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 657000 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 657000 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 657000 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 657000 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 657000 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 657000 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 657000 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 657000 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 13000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 657000 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 657000 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 657000 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 657000 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 657000 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 657000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 657000 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 657000 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 657000 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 657000 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 657000 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 657000 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 657000 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 657000 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 13000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 657000 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 657000 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 657000 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 657000 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 657000 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 657000 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 657000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 657000 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 657000 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 657000 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 657000 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 657000 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 657000 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 657000 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 657000 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 13000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 657000 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 657000 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 657000 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 657000 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 657000 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 657000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 657000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 657000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 657000 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 657000 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 657000 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 657000 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 657000 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 657000 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 657000 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 13000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 657000 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 657000 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 657000 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 657000 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 657000 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 657000 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 657000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 657000 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 657000 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 657000 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 657000 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 657000 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 657000 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 657000 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 657000 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 13000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 657000 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 657000 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 657000 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 657000 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 657000 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 657000 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 657000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 657000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 657000 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 657000 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 657000 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 657000 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 657000 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 657000 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 657000 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 13000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 657000 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 657000 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 657000 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 657000 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 657000 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 657000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 657000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 657000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 657000 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 657000 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 657000 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 657000 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 657000 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 657000 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 657000 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
