magic
tech sky130A
magscale 1 2
timestamp 1647133557
<< obsli1 >>
rect 1104 2159 548872 677841
<< obsm1 >>
rect 1104 2128 548872 677872
<< metal2 >>
rect 5722 679200 5778 680000
rect 17130 679200 17186 680000
rect 28630 679200 28686 680000
rect 40038 679200 40094 680000
rect 51538 679200 51594 680000
rect 62946 679200 63002 680000
rect 74446 679200 74502 680000
rect 85854 679200 85910 680000
rect 97354 679200 97410 680000
rect 108762 679200 108818 680000
rect 120262 679200 120318 680000
rect 131670 679200 131726 680000
rect 143170 679200 143226 680000
rect 154670 679200 154726 680000
rect 166078 679200 166134 680000
rect 177578 679200 177634 680000
rect 188986 679200 189042 680000
rect 200486 679200 200542 680000
rect 211894 679200 211950 680000
rect 223394 679200 223450 680000
rect 234802 679200 234858 680000
rect 246302 679200 246358 680000
rect 257710 679200 257766 680000
rect 269210 679200 269266 680000
rect 280710 679200 280766 680000
rect 292118 679200 292174 680000
rect 303618 679200 303674 680000
rect 315026 679200 315082 680000
rect 326526 679200 326582 680000
rect 337934 679200 337990 680000
rect 349434 679200 349490 680000
rect 360842 679200 360898 680000
rect 372342 679200 372398 680000
rect 383750 679200 383806 680000
rect 395250 679200 395306 680000
rect 406658 679200 406714 680000
rect 418158 679200 418214 680000
rect 429658 679200 429714 680000
rect 441066 679200 441122 680000
rect 452566 679200 452622 680000
rect 463974 679200 464030 680000
rect 475474 679200 475530 680000
rect 486882 679200 486938 680000
rect 498382 679200 498438 680000
rect 509790 679200 509846 680000
rect 521290 679200 521346 680000
rect 532698 679200 532754 680000
rect 544198 679200 544254 680000
rect 39302 0 39358 800
rect 117870 0 117926 800
rect 196438 0 196494 800
rect 275006 0 275062 800
rect 353574 0 353630 800
rect 432142 0 432198 800
rect 510710 0 510766 800
<< obsm2 >>
rect 1398 679144 5666 679266
rect 5834 679144 17074 679266
rect 17242 679144 28574 679266
rect 28742 679144 39982 679266
rect 40150 679144 51482 679266
rect 51650 679144 62890 679266
rect 63058 679144 74390 679266
rect 74558 679144 85798 679266
rect 85966 679144 97298 679266
rect 97466 679144 108706 679266
rect 108874 679144 120206 679266
rect 120374 679144 131614 679266
rect 131782 679144 143114 679266
rect 143282 679144 154614 679266
rect 154782 679144 166022 679266
rect 166190 679144 177522 679266
rect 177690 679144 188930 679266
rect 189098 679144 200430 679266
rect 200598 679144 211838 679266
rect 212006 679144 223338 679266
rect 223506 679144 234746 679266
rect 234914 679144 246246 679266
rect 246414 679144 257654 679266
rect 257822 679144 269154 679266
rect 269322 679144 280654 679266
rect 280822 679144 292062 679266
rect 292230 679144 303562 679266
rect 303730 679144 314970 679266
rect 315138 679144 326470 679266
rect 326638 679144 337878 679266
rect 338046 679144 349378 679266
rect 349546 679144 360786 679266
rect 360954 679144 372286 679266
rect 372454 679144 383694 679266
rect 383862 679144 395194 679266
rect 395362 679144 406602 679266
rect 406770 679144 418102 679266
rect 418270 679144 429602 679266
rect 429770 679144 441010 679266
rect 441178 679144 452510 679266
rect 452678 679144 463918 679266
rect 464086 679144 475418 679266
rect 475586 679144 486826 679266
rect 486994 679144 498326 679266
rect 498494 679144 509734 679266
rect 509902 679144 521234 679266
rect 521402 679144 532642 679266
rect 532810 679144 544142 679266
rect 544310 679144 548210 679266
rect 1398 856 548210 679144
rect 1398 800 39246 856
rect 39414 800 117814 856
rect 117982 800 196382 856
rect 196550 800 274950 856
rect 275118 800 353518 856
rect 353686 800 432086 856
rect 432254 800 510654 856
rect 510822 800 548210 856
<< metal3 >>
rect 0 672800 800 672920
rect 549200 672800 550000 672920
rect 0 658656 800 658776
rect 549200 658656 550000 658776
rect 0 644512 800 644632
rect 549200 644512 550000 644632
rect 0 630368 800 630488
rect 549200 630368 550000 630488
rect 0 616224 800 616344
rect 549200 616224 550000 616344
rect 0 602080 800 602200
rect 549200 602080 550000 602200
rect 0 587800 800 587920
rect 549200 587800 550000 587920
rect 0 573656 800 573776
rect 549200 573656 550000 573776
rect 0 559512 800 559632
rect 549200 559512 550000 559632
rect 0 545368 800 545488
rect 549200 545368 550000 545488
rect 0 531224 800 531344
rect 549200 531224 550000 531344
rect 0 517080 800 517200
rect 549200 517080 550000 517200
rect 0 502800 800 502920
rect 549200 502800 550000 502920
rect 0 488656 800 488776
rect 549200 488656 550000 488776
rect 0 474512 800 474632
rect 549200 474512 550000 474632
rect 0 460368 800 460488
rect 549200 460368 550000 460488
rect 0 446224 800 446344
rect 549200 446224 550000 446344
rect 0 432080 800 432200
rect 549200 432080 550000 432200
rect 0 417800 800 417920
rect 549200 417800 550000 417920
rect 0 403656 800 403776
rect 549200 403656 550000 403776
rect 0 389512 800 389632
rect 549200 389512 550000 389632
rect 0 375368 800 375488
rect 549200 375368 550000 375488
rect 0 361224 800 361344
rect 549200 361224 550000 361344
rect 0 347080 800 347200
rect 549200 347080 550000 347200
rect 0 332800 800 332920
rect 549200 332800 550000 332920
rect 0 318656 800 318776
rect 549200 318656 550000 318776
rect 0 304512 800 304632
rect 549200 304512 550000 304632
rect 0 290368 800 290488
rect 549200 290368 550000 290488
rect 0 276224 800 276344
rect 549200 276224 550000 276344
rect 0 262080 800 262200
rect 549200 262080 550000 262200
rect 0 247800 800 247920
rect 549200 247800 550000 247920
rect 0 233656 800 233776
rect 549200 233656 550000 233776
rect 0 219512 800 219632
rect 549200 219512 550000 219632
rect 0 205368 800 205488
rect 549200 205368 550000 205488
rect 0 191224 800 191344
rect 549200 191224 550000 191344
rect 0 177080 800 177200
rect 549200 177080 550000 177200
rect 0 162800 800 162920
rect 549200 162800 550000 162920
rect 0 148656 800 148776
rect 549200 148656 550000 148776
rect 0 134512 800 134632
rect 549200 134512 550000 134632
rect 0 120368 800 120488
rect 549200 120368 550000 120488
rect 0 106224 800 106344
rect 549200 106224 550000 106344
rect 0 92080 800 92200
rect 549200 92080 550000 92200
rect 0 77800 800 77920
rect 549200 77800 550000 77920
rect 0 63656 800 63776
rect 549200 63656 550000 63776
rect 0 49512 800 49632
rect 549200 49512 550000 49632
rect 0 35368 800 35488
rect 549200 35368 550000 35488
rect 0 21224 800 21344
rect 549200 21224 550000 21344
rect 0 7080 800 7200
rect 549200 7080 550000 7200
<< obsm3 >>
rect 800 673000 549200 677857
rect 880 672720 549120 673000
rect 800 658856 549200 672720
rect 880 658576 549120 658856
rect 800 644712 549200 658576
rect 880 644432 549120 644712
rect 800 630568 549200 644432
rect 880 630288 549120 630568
rect 800 616424 549200 630288
rect 880 616144 549120 616424
rect 800 602280 549200 616144
rect 880 602000 549120 602280
rect 800 588000 549200 602000
rect 880 587720 549120 588000
rect 800 573856 549200 587720
rect 880 573576 549120 573856
rect 800 559712 549200 573576
rect 880 559432 549120 559712
rect 800 545568 549200 559432
rect 880 545288 549120 545568
rect 800 531424 549200 545288
rect 880 531144 549120 531424
rect 800 517280 549200 531144
rect 880 517000 549120 517280
rect 800 503000 549200 517000
rect 880 502720 549120 503000
rect 800 488856 549200 502720
rect 880 488576 549120 488856
rect 800 474712 549200 488576
rect 880 474432 549120 474712
rect 800 460568 549200 474432
rect 880 460288 549120 460568
rect 800 446424 549200 460288
rect 880 446144 549120 446424
rect 800 432280 549200 446144
rect 880 432000 549120 432280
rect 800 418000 549200 432000
rect 880 417720 549120 418000
rect 800 403856 549200 417720
rect 880 403576 549120 403856
rect 800 389712 549200 403576
rect 880 389432 549120 389712
rect 800 375568 549200 389432
rect 880 375288 549120 375568
rect 800 361424 549200 375288
rect 880 361144 549120 361424
rect 800 347280 549200 361144
rect 880 347000 549120 347280
rect 800 333000 549200 347000
rect 880 332720 549120 333000
rect 800 318856 549200 332720
rect 880 318576 549120 318856
rect 800 304712 549200 318576
rect 880 304432 549120 304712
rect 800 290568 549200 304432
rect 880 290288 549120 290568
rect 800 276424 549200 290288
rect 880 276144 549120 276424
rect 800 262280 549200 276144
rect 880 262000 549120 262280
rect 800 248000 549200 262000
rect 880 247720 549120 248000
rect 800 233856 549200 247720
rect 880 233576 549120 233856
rect 800 219712 549200 233576
rect 880 219432 549120 219712
rect 800 205568 549200 219432
rect 880 205288 549120 205568
rect 800 191424 549200 205288
rect 880 191144 549120 191424
rect 800 177280 549200 191144
rect 880 177000 549120 177280
rect 800 163000 549200 177000
rect 880 162720 549120 163000
rect 800 148856 549200 162720
rect 880 148576 549120 148856
rect 800 134712 549200 148576
rect 880 134432 549120 134712
rect 800 120568 549200 134432
rect 880 120288 549120 120568
rect 800 106424 549200 120288
rect 880 106144 549120 106424
rect 800 92280 549200 106144
rect 880 92000 549120 92280
rect 800 78000 549200 92000
rect 880 77720 549120 78000
rect 800 63856 549200 77720
rect 880 63576 549120 63856
rect 800 49712 549200 63576
rect 880 49432 549120 49712
rect 800 35568 549200 49432
rect 880 35288 549120 35568
rect 800 21424 549200 35288
rect 880 21144 549120 21424
rect 800 7280 549200 21144
rect 880 7000 549120 7280
rect 800 2143 549200 7000
<< metal4 >>
rect 4208 2128 4528 677872
rect 19568 2128 19888 677872
rect 34928 2128 35248 677872
rect 50288 2128 50608 677872
rect 65648 2128 65968 677872
rect 81008 2128 81328 677872
rect 96368 2128 96688 677872
rect 111728 2128 112048 677872
rect 127088 2128 127408 677872
rect 142448 2128 142768 677872
rect 157808 2128 158128 677872
rect 173168 2128 173488 677872
rect 188528 2128 188848 677872
rect 203888 2128 204208 677872
rect 219248 2128 219568 677872
rect 234608 2128 234928 677872
rect 249968 2128 250288 677872
rect 265328 2128 265648 677872
rect 280688 2128 281008 677872
rect 296048 2128 296368 677872
rect 311408 2128 311728 677872
rect 326768 2128 327088 677872
rect 342128 2128 342448 677872
rect 357488 2128 357808 677872
rect 372848 2128 373168 677872
rect 388208 2128 388528 677872
rect 403568 2128 403888 677872
rect 418928 2128 419248 677872
rect 434288 2128 434608 677872
rect 449648 2128 449968 677872
rect 465008 2128 465328 677872
rect 480368 2128 480688 677872
rect 495728 2128 496048 677872
rect 511088 2128 511408 677872
rect 526448 2128 526768 677872
rect 541808 2128 542128 677872
<< obsm4 >>
rect 27107 2347 34848 677653
rect 35328 2347 50208 677653
rect 50688 2347 65568 677653
rect 66048 2347 80928 677653
rect 81408 2347 96288 677653
rect 96768 2347 111648 677653
rect 112128 2347 127008 677653
rect 127488 2347 142368 677653
rect 142848 2347 157728 677653
rect 158208 2347 173088 677653
rect 173568 2347 188448 677653
rect 188928 2347 203808 677653
rect 204288 2347 219168 677653
rect 219648 2347 234528 677653
rect 235008 2347 249888 677653
rect 250368 2347 265248 677653
rect 265728 2347 280608 677653
rect 281088 2347 295968 677653
rect 296448 2347 311328 677653
rect 311808 2347 326688 677653
rect 327168 2347 342048 677653
rect 342528 2347 357408 677653
rect 357888 2347 372768 677653
rect 373248 2347 388128 677653
rect 388608 2347 403488 677653
rect 403968 2347 418848 677653
rect 419328 2347 434208 677653
rect 434688 2347 449568 677653
rect 450048 2347 464928 677653
rect 465408 2347 480288 677653
rect 480768 2347 495648 677653
rect 496128 2347 496373 677653
<< labels >>
rlabel metal3 s 0 7080 800 7200 6 ipin_x0y1_0
port 1 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 ipin_x0y1_1
port 2 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 ipin_x0y2_0
port 3 nsew signal input
rlabel metal3 s 0 49512 800 49632 6 ipin_x0y2_1
port 4 nsew signal input
rlabel metal3 s 0 63656 800 63776 6 ipin_x0y3_0
port 5 nsew signal input
rlabel metal3 s 0 77800 800 77920 6 ipin_x0y3_1
port 6 nsew signal input
rlabel metal3 s 0 92080 800 92200 6 ipin_x0y4_0
port 7 nsew signal input
rlabel metal3 s 0 106224 800 106344 6 ipin_x0y4_1
port 8 nsew signal input
rlabel metal3 s 0 120368 800 120488 6 ipin_x0y5_0
port 9 nsew signal input
rlabel metal3 s 0 134512 800 134632 6 ipin_x0y5_1
port 10 nsew signal input
rlabel metal3 s 0 148656 800 148776 6 ipin_x0y6_0
port 11 nsew signal input
rlabel metal3 s 0 162800 800 162920 6 ipin_x0y6_1
port 12 nsew signal input
rlabel metal3 s 0 177080 800 177200 6 ipin_x0y7_0
port 13 nsew signal input
rlabel metal3 s 0 191224 800 191344 6 ipin_x0y7_1
port 14 nsew signal input
rlabel metal3 s 0 205368 800 205488 6 ipin_x0y8_0
port 15 nsew signal input
rlabel metal3 s 0 219512 800 219632 6 ipin_x0y8_1
port 16 nsew signal input
rlabel metal2 s 5722 679200 5778 680000 6 ipin_x1y9_0
port 17 nsew signal input
rlabel metal2 s 17130 679200 17186 680000 6 ipin_x1y9_1
port 18 nsew signal input
rlabel metal2 s 28630 679200 28686 680000 6 ipin_x2y9_0
port 19 nsew signal input
rlabel metal2 s 40038 679200 40094 680000 6 ipin_x2y9_1
port 20 nsew signal input
rlabel metal2 s 51538 679200 51594 680000 6 ipin_x3y9_0
port 21 nsew signal input
rlabel metal2 s 62946 679200 63002 680000 6 ipin_x3y9_1
port 22 nsew signal input
rlabel metal2 s 74446 679200 74502 680000 6 ipin_x4y9_0
port 23 nsew signal input
rlabel metal2 s 85854 679200 85910 680000 6 ipin_x4y9_1
port 24 nsew signal input
rlabel metal2 s 97354 679200 97410 680000 6 ipin_x5y9_0
port 25 nsew signal input
rlabel metal2 s 108762 679200 108818 680000 6 ipin_x5y9_1
port 26 nsew signal input
rlabel metal2 s 120262 679200 120318 680000 6 ipin_x6y9_0
port 27 nsew signal input
rlabel metal2 s 131670 679200 131726 680000 6 ipin_x6y9_1
port 28 nsew signal input
rlabel metal2 s 143170 679200 143226 680000 6 ipin_x7y9_0
port 29 nsew signal input
rlabel metal2 s 154670 679200 154726 680000 6 ipin_x7y9_1
port 30 nsew signal input
rlabel metal2 s 166078 679200 166134 680000 6 ipin_x8y9_0
port 31 nsew signal input
rlabel metal2 s 177578 679200 177634 680000 6 ipin_x8y9_1
port 32 nsew signal input
rlabel metal3 s 549200 7080 550000 7200 6 ipin_x9y1_0
port 33 nsew signal input
rlabel metal3 s 549200 21224 550000 21344 6 ipin_x9y1_1
port 34 nsew signal input
rlabel metal3 s 549200 35368 550000 35488 6 ipin_x9y2_0
port 35 nsew signal input
rlabel metal3 s 549200 49512 550000 49632 6 ipin_x9y2_1
port 36 nsew signal input
rlabel metal3 s 549200 63656 550000 63776 6 ipin_x9y3_0
port 37 nsew signal input
rlabel metal3 s 549200 77800 550000 77920 6 ipin_x9y3_1
port 38 nsew signal input
rlabel metal3 s 549200 92080 550000 92200 6 ipin_x9y4_0
port 39 nsew signal input
rlabel metal3 s 549200 106224 550000 106344 6 ipin_x9y4_1
port 40 nsew signal input
rlabel metal3 s 549200 120368 550000 120488 6 ipin_x9y5_0
port 41 nsew signal input
rlabel metal3 s 549200 134512 550000 134632 6 ipin_x9y5_1
port 42 nsew signal input
rlabel metal3 s 549200 148656 550000 148776 6 ipin_x9y6_0
port 43 nsew signal input
rlabel metal3 s 549200 162800 550000 162920 6 ipin_x9y6_1
port 44 nsew signal input
rlabel metal3 s 549200 177080 550000 177200 6 ipin_x9y7_0
port 45 nsew signal input
rlabel metal3 s 549200 191224 550000 191344 6 ipin_x9y7_1
port 46 nsew signal input
rlabel metal3 s 549200 205368 550000 205488 6 ipin_x9y8_0
port 47 nsew signal input
rlabel metal3 s 549200 219512 550000 219632 6 ipin_x9y8_1
port 48 nsew signal input
rlabel metal3 s 0 460368 800 460488 6 oe_x0y1_0
port 49 nsew signal output
rlabel metal3 s 0 474512 800 474632 6 oe_x0y1_1
port 50 nsew signal output
rlabel metal3 s 0 488656 800 488776 6 oe_x0y2_0
port 51 nsew signal output
rlabel metal3 s 0 502800 800 502920 6 oe_x0y2_1
port 52 nsew signal output
rlabel metal3 s 0 517080 800 517200 6 oe_x0y3_0
port 53 nsew signal output
rlabel metal3 s 0 531224 800 531344 6 oe_x0y3_1
port 54 nsew signal output
rlabel metal3 s 0 545368 800 545488 6 oe_x0y4_0
port 55 nsew signal output
rlabel metal3 s 0 559512 800 559632 6 oe_x0y4_1
port 56 nsew signal output
rlabel metal3 s 0 573656 800 573776 6 oe_x0y5_0
port 57 nsew signal output
rlabel metal3 s 0 587800 800 587920 6 oe_x0y5_1
port 58 nsew signal output
rlabel metal3 s 0 602080 800 602200 6 oe_x0y6_0
port 59 nsew signal output
rlabel metal3 s 0 616224 800 616344 6 oe_x0y6_1
port 60 nsew signal output
rlabel metal3 s 0 630368 800 630488 6 oe_x0y7_0
port 61 nsew signal output
rlabel metal3 s 0 644512 800 644632 6 oe_x0y7_1
port 62 nsew signal output
rlabel metal3 s 0 658656 800 658776 6 oe_x0y8_0
port 63 nsew signal output
rlabel metal3 s 0 672800 800 672920 6 oe_x0y8_1
port 64 nsew signal output
rlabel metal2 s 372342 679200 372398 680000 6 oe_x1y9_0
port 65 nsew signal output
rlabel metal2 s 383750 679200 383806 680000 6 oe_x1y9_1
port 66 nsew signal output
rlabel metal2 s 395250 679200 395306 680000 6 oe_x2y9_0
port 67 nsew signal output
rlabel metal2 s 406658 679200 406714 680000 6 oe_x2y9_1
port 68 nsew signal output
rlabel metal2 s 418158 679200 418214 680000 6 oe_x3y9_0
port 69 nsew signal output
rlabel metal2 s 429658 679200 429714 680000 6 oe_x3y9_1
port 70 nsew signal output
rlabel metal2 s 441066 679200 441122 680000 6 oe_x4y9_0
port 71 nsew signal output
rlabel metal2 s 452566 679200 452622 680000 6 oe_x4y9_1
port 72 nsew signal output
rlabel metal2 s 463974 679200 464030 680000 6 oe_x5y9_0
port 73 nsew signal output
rlabel metal2 s 475474 679200 475530 680000 6 oe_x5y9_1
port 74 nsew signal output
rlabel metal2 s 486882 679200 486938 680000 6 oe_x6y9_0
port 75 nsew signal output
rlabel metal2 s 498382 679200 498438 680000 6 oe_x6y9_1
port 76 nsew signal output
rlabel metal2 s 509790 679200 509846 680000 6 oe_x7y9_0
port 77 nsew signal output
rlabel metal2 s 521290 679200 521346 680000 6 oe_x7y9_1
port 78 nsew signal output
rlabel metal2 s 532698 679200 532754 680000 6 oe_x8y9_0
port 79 nsew signal output
rlabel metal2 s 544198 679200 544254 680000 6 oe_x8y9_1
port 80 nsew signal output
rlabel metal3 s 549200 460368 550000 460488 6 oe_x9y1_0
port 81 nsew signal output
rlabel metal3 s 549200 474512 550000 474632 6 oe_x9y1_1
port 82 nsew signal output
rlabel metal3 s 549200 488656 550000 488776 6 oe_x9y2_0
port 83 nsew signal output
rlabel metal3 s 549200 502800 550000 502920 6 oe_x9y2_1
port 84 nsew signal output
rlabel metal3 s 549200 517080 550000 517200 6 oe_x9y3_0
port 85 nsew signal output
rlabel metal3 s 549200 531224 550000 531344 6 oe_x9y3_1
port 86 nsew signal output
rlabel metal3 s 549200 545368 550000 545488 6 oe_x9y4_0
port 87 nsew signal output
rlabel metal3 s 549200 559512 550000 559632 6 oe_x9y4_1
port 88 nsew signal output
rlabel metal3 s 549200 573656 550000 573776 6 oe_x9y5_0
port 89 nsew signal output
rlabel metal3 s 549200 587800 550000 587920 6 oe_x9y5_1
port 90 nsew signal output
rlabel metal3 s 549200 602080 550000 602200 6 oe_x9y6_0
port 91 nsew signal output
rlabel metal3 s 549200 616224 550000 616344 6 oe_x9y6_1
port 92 nsew signal output
rlabel metal3 s 549200 630368 550000 630488 6 oe_x9y7_0
port 93 nsew signal output
rlabel metal3 s 549200 644512 550000 644632 6 oe_x9y7_1
port 94 nsew signal output
rlabel metal3 s 549200 658656 550000 658776 6 oe_x9y8_0
port 95 nsew signal output
rlabel metal3 s 549200 672800 550000 672920 6 oe_x9y8_1
port 96 nsew signal output
rlabel metal3 s 0 233656 800 233776 6 opin_x0y1_0
port 97 nsew signal output
rlabel metal3 s 0 247800 800 247920 6 opin_x0y1_1
port 98 nsew signal output
rlabel metal3 s 0 262080 800 262200 6 opin_x0y2_0
port 99 nsew signal output
rlabel metal3 s 0 276224 800 276344 6 opin_x0y2_1
port 100 nsew signal output
rlabel metal3 s 0 290368 800 290488 6 opin_x0y3_0
port 101 nsew signal output
rlabel metal3 s 0 304512 800 304632 6 opin_x0y3_1
port 102 nsew signal output
rlabel metal3 s 0 318656 800 318776 6 opin_x0y4_0
port 103 nsew signal output
rlabel metal3 s 0 332800 800 332920 6 opin_x0y4_1
port 104 nsew signal output
rlabel metal3 s 0 347080 800 347200 6 opin_x0y5_0
port 105 nsew signal output
rlabel metal3 s 0 361224 800 361344 6 opin_x0y5_1
port 106 nsew signal output
rlabel metal3 s 0 375368 800 375488 6 opin_x0y6_0
port 107 nsew signal output
rlabel metal3 s 0 389512 800 389632 6 opin_x0y6_1
port 108 nsew signal output
rlabel metal3 s 0 403656 800 403776 6 opin_x0y7_0
port 109 nsew signal output
rlabel metal3 s 0 417800 800 417920 6 opin_x0y7_1
port 110 nsew signal output
rlabel metal3 s 0 432080 800 432200 6 opin_x0y8_0
port 111 nsew signal output
rlabel metal3 s 0 446224 800 446344 6 opin_x0y8_1
port 112 nsew signal output
rlabel metal2 s 188986 679200 189042 680000 6 opin_x1y9_0
port 113 nsew signal output
rlabel metal2 s 200486 679200 200542 680000 6 opin_x1y9_1
port 114 nsew signal output
rlabel metal2 s 211894 679200 211950 680000 6 opin_x2y9_0
port 115 nsew signal output
rlabel metal2 s 223394 679200 223450 680000 6 opin_x2y9_1
port 116 nsew signal output
rlabel metal2 s 234802 679200 234858 680000 6 opin_x3y9_0
port 117 nsew signal output
rlabel metal2 s 246302 679200 246358 680000 6 opin_x3y9_1
port 118 nsew signal output
rlabel metal2 s 257710 679200 257766 680000 6 opin_x4y9_0
port 119 nsew signal output
rlabel metal2 s 269210 679200 269266 680000 6 opin_x4y9_1
port 120 nsew signal output
rlabel metal2 s 280710 679200 280766 680000 6 opin_x5y9_0
port 121 nsew signal output
rlabel metal2 s 292118 679200 292174 680000 6 opin_x5y9_1
port 122 nsew signal output
rlabel metal2 s 303618 679200 303674 680000 6 opin_x6y9_0
port 123 nsew signal output
rlabel metal2 s 315026 679200 315082 680000 6 opin_x6y9_1
port 124 nsew signal output
rlabel metal2 s 326526 679200 326582 680000 6 opin_x7y9_0
port 125 nsew signal output
rlabel metal2 s 337934 679200 337990 680000 6 opin_x7y9_1
port 126 nsew signal output
rlabel metal2 s 349434 679200 349490 680000 6 opin_x8y9_0
port 127 nsew signal output
rlabel metal2 s 360842 679200 360898 680000 6 opin_x8y9_1
port 128 nsew signal output
rlabel metal3 s 549200 233656 550000 233776 6 opin_x9y1_0
port 129 nsew signal output
rlabel metal3 s 549200 247800 550000 247920 6 opin_x9y1_1
port 130 nsew signal output
rlabel metal3 s 549200 262080 550000 262200 6 opin_x9y2_0
port 131 nsew signal output
rlabel metal3 s 549200 276224 550000 276344 6 opin_x9y2_1
port 132 nsew signal output
rlabel metal3 s 549200 290368 550000 290488 6 opin_x9y3_0
port 133 nsew signal output
rlabel metal3 s 549200 304512 550000 304632 6 opin_x9y3_1
port 134 nsew signal output
rlabel metal3 s 549200 318656 550000 318776 6 opin_x9y4_0
port 135 nsew signal output
rlabel metal3 s 549200 332800 550000 332920 6 opin_x9y4_1
port 136 nsew signal output
rlabel metal3 s 549200 347080 550000 347200 6 opin_x9y5_0
port 137 nsew signal output
rlabel metal3 s 549200 361224 550000 361344 6 opin_x9y5_1
port 138 nsew signal output
rlabel metal3 s 549200 375368 550000 375488 6 opin_x9y6_0
port 139 nsew signal output
rlabel metal3 s 549200 389512 550000 389632 6 opin_x9y6_1
port 140 nsew signal output
rlabel metal3 s 549200 403656 550000 403776 6 opin_x9y7_0
port 141 nsew signal output
rlabel metal3 s 549200 417800 550000 417920 6 opin_x9y7_1
port 142 nsew signal output
rlabel metal3 s 549200 432080 550000 432200 6 opin_x9y8_0
port 143 nsew signal output
rlabel metal3 s 549200 446224 550000 446344 6 opin_x9y8_1
port 144 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 prog_clk
port 145 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 prog_din
port 146 nsew signal input
rlabel metal2 s 196438 0 196494 800 6 prog_done
port 147 nsew signal input
rlabel metal2 s 275006 0 275062 800 6 prog_dout
port 148 nsew signal output
rlabel metal2 s 353574 0 353630 800 6 prog_rst
port 149 nsew signal input
rlabel metal2 s 432142 0 432198 800 6 prog_we
port 150 nsew signal input
rlabel metal2 s 510710 0 510766 800 6 prog_we_o
port 151 nsew signal output
rlabel metal4 s 4208 2128 4528 677872 6 vccd1
port 152 nsew power input
rlabel metal4 s 34928 2128 35248 677872 6 vccd1
port 152 nsew power input
rlabel metal4 s 65648 2128 65968 677872 6 vccd1
port 152 nsew power input
rlabel metal4 s 96368 2128 96688 677872 6 vccd1
port 152 nsew power input
rlabel metal4 s 127088 2128 127408 677872 6 vccd1
port 152 nsew power input
rlabel metal4 s 157808 2128 158128 677872 6 vccd1
port 152 nsew power input
rlabel metal4 s 188528 2128 188848 677872 6 vccd1
port 152 nsew power input
rlabel metal4 s 219248 2128 219568 677872 6 vccd1
port 152 nsew power input
rlabel metal4 s 249968 2128 250288 677872 6 vccd1
port 152 nsew power input
rlabel metal4 s 280688 2128 281008 677872 6 vccd1
port 152 nsew power input
rlabel metal4 s 311408 2128 311728 677872 6 vccd1
port 152 nsew power input
rlabel metal4 s 342128 2128 342448 677872 6 vccd1
port 152 nsew power input
rlabel metal4 s 372848 2128 373168 677872 6 vccd1
port 152 nsew power input
rlabel metal4 s 403568 2128 403888 677872 6 vccd1
port 152 nsew power input
rlabel metal4 s 434288 2128 434608 677872 6 vccd1
port 152 nsew power input
rlabel metal4 s 465008 2128 465328 677872 6 vccd1
port 152 nsew power input
rlabel metal4 s 495728 2128 496048 677872 6 vccd1
port 152 nsew power input
rlabel metal4 s 526448 2128 526768 677872 6 vccd1
port 152 nsew power input
rlabel metal4 s 19568 2128 19888 677872 6 vssd1
port 153 nsew ground input
rlabel metal4 s 50288 2128 50608 677872 6 vssd1
port 153 nsew ground input
rlabel metal4 s 81008 2128 81328 677872 6 vssd1
port 153 nsew ground input
rlabel metal4 s 111728 2128 112048 677872 6 vssd1
port 153 nsew ground input
rlabel metal4 s 142448 2128 142768 677872 6 vssd1
port 153 nsew ground input
rlabel metal4 s 173168 2128 173488 677872 6 vssd1
port 153 nsew ground input
rlabel metal4 s 203888 2128 204208 677872 6 vssd1
port 153 nsew ground input
rlabel metal4 s 234608 2128 234928 677872 6 vssd1
port 153 nsew ground input
rlabel metal4 s 265328 2128 265648 677872 6 vssd1
port 153 nsew ground input
rlabel metal4 s 296048 2128 296368 677872 6 vssd1
port 153 nsew ground input
rlabel metal4 s 326768 2128 327088 677872 6 vssd1
port 153 nsew ground input
rlabel metal4 s 357488 2128 357808 677872 6 vssd1
port 153 nsew ground input
rlabel metal4 s 388208 2128 388528 677872 6 vssd1
port 153 nsew ground input
rlabel metal4 s 418928 2128 419248 677872 6 vssd1
port 153 nsew ground input
rlabel metal4 s 449648 2128 449968 677872 6 vssd1
port 153 nsew ground input
rlabel metal4 s 480368 2128 480688 677872 6 vssd1
port 153 nsew ground input
rlabel metal4 s 511088 2128 511408 677872 6 vssd1
port 153 nsew ground input
rlabel metal4 s 541808 2128 542128 677872 6 vssd1
port 153 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 550000 680000
string LEFview TRUE
string GDS_FILE /files/research/projects/tapeout/caravel_mpw5_prga/openlane/prga/runs/prga/results/magic/top.gds
string GDS_END 261387618
string GDS_START 6170262
<< end >>

